magic
tech sky130A
magscale 1 2
timestamp 1671820617
<< viali >>
rect 7849 13481 7883 13515
rect 8401 13481 8435 13515
rect 10241 13481 10275 13515
rect 13553 13481 13587 13515
rect 17233 13481 17267 13515
rect 17969 13481 18003 13515
rect 18705 13481 18739 13515
rect 20637 13481 20671 13515
rect 22385 13481 22419 13515
rect 27629 13481 27663 13515
rect 28365 13481 28399 13515
rect 29101 13481 29135 13515
rect 32781 13481 32815 13515
rect 33425 13481 33459 13515
rect 37841 13481 37875 13515
rect 44649 13481 44683 13515
rect 55689 13481 55723 13515
rect 60105 13481 60139 13515
rect 65993 13481 66027 13515
rect 66637 13481 66671 13515
rect 67649 13481 67683 13515
rect 68845 13481 68879 13515
rect 69489 13481 69523 13515
rect 70225 13481 70259 13515
rect 71329 13481 71363 13515
rect 72065 13481 72099 13515
rect 72801 13481 72835 13515
rect 73905 13481 73939 13515
rect 74641 13481 74675 13515
rect 75469 13481 75503 13515
rect 76205 13481 76239 13515
rect 78045 13481 78079 13515
rect 78965 13481 78999 13515
rect 79793 13481 79827 13515
rect 80437 13481 80471 13515
rect 81449 13481 81483 13515
rect 82829 13481 82863 13515
rect 83933 13481 83967 13515
rect 85405 13481 85439 13515
rect 90649 13481 90683 13515
rect 94237 13481 94271 13515
rect 97549 13481 97583 13515
rect 99389 13481 99423 13515
rect 104541 13481 104575 13515
rect 106105 13481 106139 13515
rect 107025 13481 107059 13515
rect 110429 13481 110463 13515
rect 112269 13481 112303 13515
rect 113741 13481 113775 13515
rect 114937 13481 114971 13515
rect 118157 13481 118191 13515
rect 119997 13481 120031 13515
rect 121469 13481 121503 13515
rect 125149 13481 125183 13515
rect 126621 13481 126655 13515
rect 129197 13481 129231 13515
rect 131037 13481 131071 13515
rect 131773 13481 131807 13515
rect 132969 13481 133003 13515
rect 135453 13481 135487 13515
rect 136281 13481 136315 13515
rect 137017 13481 137051 13515
rect 138029 13481 138063 13515
rect 138765 13481 138799 13515
rect 139593 13481 139627 13515
rect 140605 13481 140639 13515
rect 141433 13481 141467 13515
rect 147321 13481 147355 13515
rect 153577 13481 153611 13515
rect 154313 13481 154347 13515
rect 156153 13481 156187 13515
rect 9597 13413 9631 13447
rect 12173 13413 12207 13447
rect 19901 13413 19935 13447
rect 21281 13413 21315 13447
rect 23121 13413 23155 13447
rect 34161 13413 34195 13447
rect 34897 13413 34931 13447
rect 48421 13413 48455 13447
rect 54953 13413 54987 13447
rect 62221 13413 62255 13447
rect 82093 13413 82127 13447
rect 87061 13413 87095 13447
rect 91753 13413 91787 13447
rect 95709 13413 95743 13447
rect 96813 13413 96847 13447
rect 98377 13413 98411 13447
rect 100217 13413 100251 13447
rect 103161 13413 103195 13447
rect 105277 13413 105311 13447
rect 109693 13413 109727 13447
rect 111165 13413 111199 13447
rect 113097 13413 113131 13447
rect 116409 13413 116443 13447
rect 117513 13413 117547 13447
rect 118893 13413 118927 13447
rect 120733 13413 120767 13447
rect 123861 13413 123895 13447
rect 125885 13413 125919 13447
rect 127725 13413 127759 13447
rect 128461 13413 128495 13447
rect 130301 13413 130335 13447
rect 133705 13413 133739 13447
rect 134441 13413 134475 13447
rect 142169 13413 142203 13447
rect 149621 13413 149655 13447
rect 150081 13413 150115 13447
rect 150817 13413 150851 13447
rect 156889 13413 156923 13447
rect 122481 13345 122515 13379
rect 143089 13345 143123 13379
rect 8585 13277 8619 13311
rect 9413 13277 9447 13311
rect 10425 13277 10459 13311
rect 11161 13277 11195 13311
rect 11989 13277 12023 13311
rect 12725 13277 12759 13311
rect 13737 13277 13771 13311
rect 15669 13277 15703 13311
rect 17417 13277 17451 13311
rect 18153 13277 18187 13311
rect 18889 13277 18923 13311
rect 19717 13277 19751 13311
rect 20453 13277 20487 13311
rect 21465 13277 21499 13311
rect 22569 13277 22603 13311
rect 23305 13277 23339 13311
rect 23765 13277 23799 13311
rect 25237 13277 25271 13311
rect 27445 13277 27479 13311
rect 28181 13277 28215 13311
rect 28917 13277 28951 13311
rect 30205 13277 30239 13311
rect 32597 13277 32631 13311
rect 33609 13277 33643 13311
rect 34345 13277 34379 13311
rect 36021 13277 36055 13311
rect 36277 13277 36311 13311
rect 38025 13277 38059 13311
rect 38761 13277 38795 13311
rect 39497 13277 39531 13311
rect 40233 13277 40267 13311
rect 40417 13277 40451 13311
rect 41245 13277 41279 13311
rect 41705 13277 41739 13311
rect 41889 13277 41923 13311
rect 42073 13277 42107 13311
rect 42625 13277 42659 13311
rect 43269 13277 43303 13311
rect 46581 13277 46615 13311
rect 47961 13277 47995 13311
rect 49801 13277 49835 13311
rect 52377 13277 52411 13311
rect 53573 13277 53607 13311
rect 55505 13277 55539 13311
rect 56149 13277 56183 13311
rect 56405 13277 56439 13311
rect 58725 13277 58759 13311
rect 60841 13277 60875 13311
rect 63417 13277 63451 13311
rect 63509 13277 63543 13311
rect 65809 13277 65843 13311
rect 67833 13277 67867 13311
rect 68661 13277 68695 13311
rect 69673 13277 69707 13311
rect 70409 13277 70443 13311
rect 71513 13277 71547 13311
rect 72249 13277 72283 13311
rect 72985 13277 73019 13311
rect 74089 13277 74123 13311
rect 74825 13277 74859 13311
rect 75285 13277 75319 13311
rect 76389 13277 76423 13311
rect 77235 13277 77269 13311
rect 77861 13277 77895 13311
rect 79149 13277 79183 13311
rect 79609 13277 79643 13311
rect 80621 13277 80655 13311
rect 81265 13277 81299 13311
rect 82277 13277 82311 13311
rect 83013 13277 83047 13311
rect 84117 13277 84151 13311
rect 84853 13277 84887 13311
rect 85589 13277 85623 13311
rect 88441 13277 88475 13311
rect 89637 13277 89671 13311
rect 90833 13277 90867 13311
rect 93133 13277 93167 13311
rect 94421 13277 94455 13311
rect 95157 13277 95191 13311
rect 95893 13277 95927 13311
rect 96997 13277 97031 13311
rect 97733 13277 97767 13311
rect 98193 13277 98227 13311
rect 99573 13277 99607 13311
rect 100033 13277 100067 13311
rect 101045 13277 101079 13311
rect 102333 13277 102367 13311
rect 102425 13277 102459 13311
rect 103345 13277 103379 13311
rect 104725 13277 104759 13311
rect 105461 13277 105495 13311
rect 105921 13277 105955 13311
rect 107669 13277 107703 13311
rect 109877 13277 109911 13311
rect 110613 13277 110647 13311
rect 111349 13277 111383 13311
rect 112453 13277 112487 13311
rect 112919 13277 112953 13311
rect 113925 13277 113959 13311
rect 114753 13277 114787 13311
rect 115765 13277 115799 13311
rect 116225 13277 116259 13311
rect 117329 13277 117363 13311
rect 118341 13277 118375 13311
rect 119077 13277 119111 13311
rect 120181 13277 120215 13311
rect 120917 13277 120951 13311
rect 121653 13277 121687 13311
rect 125333 13277 125367 13311
rect 126069 13277 126103 13311
rect 126805 13277 126839 13311
rect 127909 13277 127943 13311
rect 128645 13277 128679 13311
rect 129381 13277 129415 13311
rect 130485 13277 130519 13311
rect 131221 13277 131255 13311
rect 131957 13277 131991 13311
rect 132785 13277 132819 13311
rect 133521 13277 133555 13311
rect 134257 13277 134291 13311
rect 135637 13277 135671 13311
rect 136097 13277 136131 13311
rect 136833 13277 136867 13311
rect 138213 13277 138247 13311
rect 138949 13277 138983 13311
rect 139409 13277 139443 13311
rect 140789 13277 140823 13311
rect 141249 13277 141283 13311
rect 141985 13277 142019 13311
rect 143733 13277 143767 13311
rect 145941 13277 145975 13311
rect 148241 13277 148275 13311
rect 150265 13277 150299 13311
rect 152197 13277 152231 13311
rect 152841 13277 152875 13311
rect 153393 13277 153427 13311
rect 154129 13277 154163 13311
rect 154865 13277 154899 13311
rect 155969 13277 156003 13311
rect 156705 13277 156739 13311
rect 157441 13277 157475 13311
rect 15402 13209 15436 13243
rect 16313 13209 16347 13243
rect 25504 13209 25538 13243
rect 30472 13209 30506 13243
rect 43536 13209 43570 13243
rect 46314 13209 46348 13243
rect 49534 13209 49568 13243
rect 52132 13209 52166 13243
rect 53840 13209 53874 13243
rect 58970 13209 59004 13243
rect 61108 13209 61142 13243
rect 64337 13209 64371 13243
rect 65165 13209 65199 13243
rect 66913 13209 66947 13243
rect 88196 13209 88230 13243
rect 90005 13209 90039 13243
rect 92888 13209 92922 13243
rect 107936 13209 107970 13243
rect 122748 13209 122782 13243
rect 144000 13209 144034 13243
rect 146208 13209 146242 13243
rect 148508 13209 148542 13243
rect 151930 13209 151964 13243
rect 7297 13141 7331 13175
rect 10977 13141 11011 13175
rect 12909 13141 12943 13175
rect 14289 13141 14323 13175
rect 23949 13141 23983 13175
rect 24777 13141 24811 13175
rect 26617 13141 26651 13175
rect 31585 13141 31619 13175
rect 36829 13141 36863 13175
rect 38577 13141 38611 13175
rect 39313 13141 39347 13175
rect 40049 13141 40083 13175
rect 41061 13141 41095 13175
rect 42809 13141 42843 13175
rect 45201 13141 45235 13175
rect 47225 13141 47259 13175
rect 50537 13141 50571 13175
rect 50997 13141 51031 13175
rect 53113 13141 53147 13175
rect 57529 13141 57563 13175
rect 58265 13141 58299 13175
rect 63693 13141 63727 13175
rect 65073 13141 65107 13175
rect 76941 13141 76975 13175
rect 84669 13141 84703 13175
rect 86417 13141 86451 13175
rect 88993 13141 89027 13175
rect 94973 13141 95007 13175
rect 100861 13141 100895 13175
rect 102609 13141 102643 13175
rect 103805 13141 103839 13175
rect 109049 13141 109083 13175
rect 115581 13141 115615 13175
rect 124321 13141 124355 13175
rect 145113 13141 145147 13175
rect 152657 13141 152691 13175
rect 155049 13141 155083 13175
rect 157625 13141 157659 13175
rect 7297 12937 7331 12971
rect 9505 12937 9539 12971
rect 10241 12937 10275 12971
rect 15577 12937 15611 12971
rect 16129 12937 16163 12971
rect 17509 12937 17543 12971
rect 18705 12937 18739 12971
rect 19441 12937 19475 12971
rect 22661 12937 22695 12971
rect 23489 12937 23523 12971
rect 26433 12937 26467 12971
rect 32505 12937 32539 12971
rect 33517 12937 33551 12971
rect 36829 12937 36863 12971
rect 37933 12937 37967 12971
rect 38577 12937 38611 12971
rect 39405 12937 39439 12971
rect 44005 12937 44039 12971
rect 50353 12937 50387 12971
rect 57529 12937 57563 12971
rect 58909 12937 58943 12971
rect 63877 12937 63911 12971
rect 64613 12937 64647 12971
rect 65441 12937 65475 12971
rect 66085 12937 66119 12971
rect 67005 12937 67039 12971
rect 67649 12937 67683 12971
rect 68385 12937 68419 12971
rect 72249 12937 72283 12971
rect 72801 12937 72835 12971
rect 74641 12937 74675 12971
rect 75561 12937 75595 12971
rect 76573 12937 76607 12971
rect 77677 12937 77711 12971
rect 78781 12937 78815 12971
rect 79517 12937 79551 12971
rect 83013 12937 83047 12971
rect 83933 12937 83967 12971
rect 84577 12937 84611 12971
rect 88073 12937 88107 12971
rect 89085 12937 89119 12971
rect 94237 12937 94271 12971
rect 97365 12937 97399 12971
rect 98193 12937 98227 12971
rect 100953 12937 100987 12971
rect 102425 12937 102459 12971
rect 103161 12937 103195 12971
rect 104541 12937 104575 12971
rect 108313 12937 108347 12971
rect 109693 12937 109727 12971
rect 112913 12937 112947 12971
rect 113649 12937 113683 12971
rect 118525 12937 118559 12971
rect 119997 12937 120031 12971
rect 120733 12937 120767 12971
rect 121469 12937 121503 12971
rect 125149 12937 125183 12971
rect 128829 12937 128863 12971
rect 129565 12937 129599 12971
rect 130301 12937 130335 12971
rect 131037 12937 131071 12971
rect 131865 12937 131899 12971
rect 134165 12937 134199 12971
rect 135545 12937 135579 12971
rect 136833 12937 136867 12971
rect 137937 12937 137971 12971
rect 139593 12937 139627 12971
rect 140881 12937 140915 12971
rect 142905 12937 142939 12971
rect 149437 12937 149471 12971
rect 156153 12937 156187 12971
rect 156889 12937 156923 12971
rect 158085 12937 158119 12971
rect 14758 12869 14792 12903
rect 31524 12869 31558 12903
rect 34406 12869 34440 12903
rect 41806 12869 41840 12903
rect 42870 12869 42904 12903
rect 106780 12869 106814 12903
rect 112116 12869 112150 12903
rect 115020 12869 115054 12903
rect 127164 12869 127198 12903
rect 146800 12869 146834 12903
rect 9689 12801 9723 12835
rect 10425 12801 10459 12835
rect 10885 12801 10919 12835
rect 11897 12801 11931 12835
rect 13001 12801 13035 12835
rect 16313 12801 16347 12835
rect 17693 12801 17727 12835
rect 18889 12801 18923 12835
rect 19625 12801 19659 12835
rect 21209 12801 21243 12835
rect 22845 12801 22879 12835
rect 23305 12801 23339 12835
rect 25165 12801 25199 12835
rect 26617 12801 26651 12835
rect 28650 12801 28684 12835
rect 28917 12801 28951 12835
rect 29653 12801 29687 12835
rect 32321 12801 32355 12835
rect 33701 12801 33735 12835
rect 36645 12801 36679 12835
rect 37749 12801 37783 12835
rect 38761 12801 38795 12835
rect 39221 12801 39255 12835
rect 40233 12801 40267 12835
rect 42625 12801 42659 12835
rect 45109 12801 45143 12835
rect 45836 12801 45870 12835
rect 48044 12801 48078 12835
rect 50537 12801 50571 12835
rect 52110 12801 52144 12835
rect 53573 12801 53607 12835
rect 54033 12801 54067 12835
rect 54300 12801 54334 12835
rect 56405 12801 56439 12835
rect 58265 12801 58299 12835
rect 58725 12801 58759 12835
rect 60574 12801 60608 12835
rect 60841 12801 60875 12835
rect 61568 12801 61602 12835
rect 63325 12801 63359 12835
rect 64061 12801 64095 12835
rect 64797 12801 64831 12835
rect 65257 12801 65291 12835
rect 66269 12801 66303 12835
rect 66821 12801 66855 12835
rect 67833 12801 67867 12835
rect 69498 12801 69532 12835
rect 71136 12801 71170 12835
rect 72985 12801 73019 12835
rect 74089 12801 74123 12835
rect 74825 12801 74859 12835
rect 75377 12801 75411 12835
rect 76757 12801 76791 12835
rect 77861 12801 77895 12835
rect 78965 12801 78999 12835
rect 81348 12801 81382 12835
rect 83197 12801 83231 12835
rect 84117 12801 84151 12835
rect 85313 12801 85347 12835
rect 87162 12801 87196 12835
rect 87889 12801 87923 12835
rect 89269 12801 89303 12835
rect 89729 12801 89763 12835
rect 90649 12801 90683 12835
rect 91293 12801 91327 12835
rect 91560 12801 91594 12835
rect 93409 12801 93443 12835
rect 94421 12801 94455 12835
rect 95433 12801 95467 12835
rect 95700 12801 95734 12835
rect 97549 12801 97583 12835
rect 98009 12801 98043 12835
rect 99481 12801 99515 12835
rect 100125 12801 100159 12835
rect 101137 12801 101171 12835
rect 101873 12801 101907 12835
rect 102609 12801 102643 12835
rect 103345 12801 103379 12835
rect 104725 12801 104759 12835
rect 107761 12801 107795 12835
rect 108497 12801 108531 12835
rect 109049 12801 109083 12835
rect 109877 12801 109911 12835
rect 113097 12801 113131 12835
rect 113833 12801 113867 12835
rect 116593 12801 116627 12835
rect 116860 12801 116894 12835
rect 118709 12801 118743 12835
rect 120181 12801 120215 12835
rect 120917 12801 120951 12835
rect 121653 12801 121687 12835
rect 122472 12801 122506 12835
rect 124321 12801 124355 12835
rect 125333 12801 125367 12835
rect 126069 12801 126103 12835
rect 129013 12801 129047 12835
rect 130485 12801 130519 12835
rect 131221 12801 131255 12835
rect 131681 12801 131715 12835
rect 134349 12801 134383 12835
rect 135386 12801 135420 12835
rect 136649 12801 136683 12835
rect 137753 12801 137787 12835
rect 138949 12801 138983 12835
rect 139409 12801 139443 12835
rect 142005 12801 142039 12835
rect 142721 12801 142755 12835
rect 144857 12801 144891 12835
rect 145113 12801 145147 12835
rect 147045 12801 147079 12835
rect 147505 12801 147539 12835
rect 147772 12801 147806 12835
rect 149621 12801 149655 12835
rect 150265 12801 150299 12835
rect 151930 12801 151964 12835
rect 152197 12801 152231 12835
rect 153770 12801 153804 12835
rect 154037 12801 154071 12835
rect 154589 12801 154623 12835
rect 154681 12801 154715 12835
rect 155969 12801 156003 12835
rect 156705 12801 156739 12835
rect 157625 12801 157659 12835
rect 158269 12801 158303 12835
rect 8953 12733 8987 12767
rect 11713 12733 11747 12767
rect 12817 12733 12851 12767
rect 15025 12733 15059 12767
rect 16865 12733 16899 12767
rect 21465 12733 21499 12767
rect 25421 12733 25455 12767
rect 31769 12733 31803 12767
rect 34161 12733 34195 12767
rect 42073 12733 42107 12767
rect 45569 12733 45603 12767
rect 47777 12733 47811 12767
rect 52377 12733 52411 12767
rect 56149 12733 56183 12767
rect 61301 12733 61335 12767
rect 69765 12733 69799 12767
rect 70317 12733 70351 12767
rect 70869 12733 70903 12767
rect 81081 12733 81115 12767
rect 85497 12733 85531 12767
rect 87429 12733 87463 12767
rect 90465 12733 90499 12767
rect 99665 12733 99699 12767
rect 103897 12733 103931 12767
rect 107025 12733 107059 12767
rect 112361 12733 112395 12767
rect 114753 12733 114787 12767
rect 122205 12733 122239 12767
rect 126897 12733 126931 12767
rect 132785 12733 132819 12767
rect 133061 12733 133095 12767
rect 136097 12733 136131 12767
rect 142261 12733 142295 12767
rect 154865 12733 154899 12767
rect 8401 12665 8435 12699
rect 11069 12665 11103 12699
rect 24041 12665 24075 12699
rect 30389 12665 30423 12699
rect 35541 12665 35575 12699
rect 40049 12665 40083 12699
rect 46949 12665 46983 12699
rect 80529 12665 80563 12699
rect 86049 12665 86083 12699
rect 89913 12665 89947 12699
rect 92673 12665 92707 12699
rect 96813 12665 96847 12699
rect 100309 12665 100343 12699
rect 101689 12665 101723 12699
rect 105645 12665 105679 12699
rect 117973 12665 118007 12699
rect 123585 12665 123619 12699
rect 143733 12665 143767 12699
rect 148885 12665 148919 12699
rect 150081 12665 150115 12699
rect 150817 12665 150851 12699
rect 152657 12665 152691 12699
rect 155325 12665 155359 12699
rect 157441 12665 157475 12699
rect 7849 12597 7883 12631
rect 12081 12597 12115 12631
rect 13185 12597 13219 12631
rect 13645 12597 13679 12631
rect 20085 12597 20119 12631
rect 22109 12597 22143 12631
rect 27537 12597 27571 12631
rect 29837 12597 29871 12631
rect 36185 12597 36219 12631
rect 40693 12597 40727 12631
rect 44925 12597 44959 12631
rect 49157 12597 49191 12631
rect 49801 12597 49835 12631
rect 50997 12597 51031 12631
rect 53389 12597 53423 12631
rect 55413 12597 55447 12631
rect 58081 12597 58115 12631
rect 59461 12597 59495 12631
rect 62681 12597 62715 12631
rect 73905 12597 73939 12631
rect 80069 12597 80103 12631
rect 82461 12597 82495 12631
rect 85129 12597 85163 12631
rect 90833 12597 90867 12631
rect 93225 12597 93259 12631
rect 94881 12597 94915 12631
rect 99297 12597 99331 12631
rect 107577 12597 107611 12631
rect 110429 12597 110463 12631
rect 110981 12597 111015 12631
rect 116133 12597 116167 12631
rect 119169 12597 119203 12631
rect 124137 12597 124171 12631
rect 125885 12597 125919 12631
rect 128277 12597 128311 12631
rect 138765 12597 138799 12631
rect 145665 12597 145699 12631
rect 10517 12393 10551 12427
rect 13645 12393 13679 12427
rect 22109 12393 22143 12427
rect 23029 12393 23063 12427
rect 23857 12393 23891 12427
rect 27261 12393 27295 12427
rect 27997 12393 28031 12427
rect 29929 12393 29963 12427
rect 30665 12393 30699 12427
rect 32689 12393 32723 12427
rect 34069 12393 34103 12427
rect 35173 12393 35207 12427
rect 36369 12393 36403 12427
rect 37381 12393 37415 12427
rect 38577 12393 38611 12427
rect 39405 12393 39439 12427
rect 44557 12393 44591 12427
rect 49801 12393 49835 12427
rect 56425 12393 56459 12427
rect 59277 12393 59311 12427
rect 63233 12393 63267 12427
rect 63969 12393 64003 12427
rect 64981 12393 65015 12427
rect 68845 12393 68879 12427
rect 70041 12393 70075 12427
rect 72433 12393 72467 12427
rect 75377 12393 75411 12427
rect 77769 12393 77803 12427
rect 85405 12393 85439 12427
rect 86601 12393 86635 12427
rect 87797 12393 87831 12427
rect 96813 12393 96847 12427
rect 98745 12393 98779 12427
rect 99389 12393 99423 12427
rect 105369 12393 105403 12427
rect 106013 12393 106047 12427
rect 107117 12393 107151 12427
rect 110245 12393 110279 12427
rect 112269 12393 112303 12427
rect 121745 12393 121779 12427
rect 127817 12393 127851 12427
rect 128461 12393 128495 12427
rect 129013 12393 129047 12427
rect 132877 12393 132911 12427
rect 135545 12393 135579 12427
rect 141341 12393 141375 12427
rect 146953 12393 146987 12427
rect 149989 12393 150023 12427
rect 7757 12325 7791 12359
rect 26433 12325 26467 12359
rect 42257 12325 42291 12359
rect 43821 12325 43855 12359
rect 50813 12325 50847 12359
rect 54033 12325 54067 12359
rect 62405 12325 62439 12359
rect 66637 12325 66671 12359
rect 89821 12325 89855 12359
rect 90557 12325 90591 12359
rect 122481 12325 122515 12359
rect 141893 12325 141927 12359
rect 153393 12325 153427 12359
rect 156245 12325 156279 12359
rect 32045 12257 32079 12291
rect 42717 12257 42751 12291
rect 56793 12257 56827 12291
rect 76665 12257 76699 12291
rect 81265 12257 81299 12291
rect 83749 12257 83783 12291
rect 87153 12257 87187 12291
rect 94145 12257 94179 12291
rect 117881 12257 117915 12291
rect 120273 12257 120307 12291
rect 137017 12257 137051 12291
rect 155601 12257 155635 12291
rect 4629 12189 4663 12223
rect 6377 12189 6411 12223
rect 9873 12189 9907 12223
rect 10333 12189 10367 12223
rect 11069 12189 11103 12223
rect 13461 12189 13495 12223
rect 14841 12189 14875 12223
rect 15577 12189 15611 12223
rect 17417 12189 17451 12223
rect 20729 12189 20763 12223
rect 23213 12189 23247 12223
rect 24041 12189 24075 12223
rect 24593 12189 24627 12223
rect 27445 12189 27479 12223
rect 28181 12189 28215 12223
rect 29745 12189 29779 12223
rect 32505 12189 32539 12223
rect 34253 12189 34287 12223
rect 35357 12189 35391 12223
rect 36185 12189 36219 12223
rect 37565 12189 37599 12223
rect 38393 12189 38427 12223
rect 39221 12189 39255 12223
rect 40233 12189 40267 12223
rect 42073 12189 42107 12223
rect 42901 12189 42935 12223
rect 43637 12189 43671 12223
rect 44373 12189 44407 12223
rect 45477 12189 45511 12223
rect 45937 12189 45971 12223
rect 49157 12189 49191 12223
rect 50629 12189 50663 12223
rect 51641 12189 51675 12223
rect 52101 12189 52135 12223
rect 54217 12189 54251 12223
rect 55689 12189 55723 12223
rect 55873 12189 55907 12223
rect 56609 12189 56643 12223
rect 57253 12189 57287 12223
rect 59461 12189 59495 12223
rect 59553 12189 59587 12223
rect 61025 12189 61059 12223
rect 63049 12189 63083 12223
rect 63785 12189 63819 12223
rect 65165 12189 65199 12223
rect 67741 12189 67775 12223
rect 69029 12189 69063 12223
rect 69857 12189 69891 12223
rect 72893 12189 72927 12223
rect 73997 12189 74031 12223
rect 74264 12189 74298 12223
rect 79149 12189 79183 12223
rect 81449 12189 81483 12223
rect 82093 12189 82127 12223
rect 85589 12189 85623 12223
rect 86417 12189 86451 12223
rect 89177 12189 89211 12223
rect 89637 12189 89671 12223
rect 90373 12189 90407 12223
rect 92949 12189 92983 12223
rect 93685 12189 93719 12223
rect 96169 12189 96203 12223
rect 96997 12189 97031 12223
rect 97733 12189 97767 12223
rect 99941 12189 99975 12223
rect 102977 12189 103011 12223
rect 104357 12189 104391 12223
rect 104541 12189 104575 12223
rect 105185 12189 105219 12223
rect 106197 12189 106231 12223
rect 107301 12189 107335 12223
rect 109693 12189 109727 12223
rect 110429 12189 110463 12223
rect 110889 12189 110923 12223
rect 111073 12189 111107 12223
rect 112453 12189 112487 12223
rect 115397 12189 115431 12223
rect 116501 12189 116535 12223
rect 121929 12189 121963 12223
rect 123861 12189 123895 12223
rect 124597 12189 124631 12223
rect 125701 12189 125735 12223
rect 127633 12189 127667 12223
rect 130025 12189 130059 12223
rect 134165 12189 134199 12223
rect 134432 12189 134466 12223
rect 136557 12189 136591 12223
rect 138029 12189 138063 12223
rect 140513 12189 140547 12223
rect 141157 12189 141191 12223
rect 144561 12189 144595 12223
rect 146401 12189 146435 12223
rect 147137 12189 147171 12223
rect 148517 12189 148551 12223
rect 148977 12189 149011 12223
rect 151369 12189 151403 12223
rect 152013 12189 152047 12223
rect 152657 12189 152691 12223
rect 152841 12189 152875 12223
rect 154773 12189 154807 12223
rect 155417 12189 155451 12223
rect 156061 12189 156095 12223
rect 156797 12189 156831 12223
rect 157717 12189 157751 12223
rect 6644 12121 6678 12155
rect 9321 12121 9355 12155
rect 11336 12121 11370 12155
rect 13001 12121 13035 12155
rect 14381 12121 14415 12155
rect 15822 12121 15856 12155
rect 17662 12121 17696 12155
rect 20177 12121 20211 12155
rect 20974 12121 21008 12155
rect 24860 12121 24894 12155
rect 26617 12121 26651 12155
rect 31778 12121 31812 12155
rect 40478 12121 40512 12155
rect 46204 12121 46238 12155
rect 48912 12121 48946 12155
rect 52368 12121 52402 12155
rect 54769 12121 54803 12155
rect 57520 12121 57554 12155
rect 61292 12121 61326 12155
rect 67189 12121 67223 12155
rect 73537 12121 73571 12155
rect 77309 12121 77343 12155
rect 78882 12121 78916 12155
rect 88910 12121 88944 12155
rect 92704 12121 92738 12155
rect 95924 12121 95958 12155
rect 98193 12121 98227 12155
rect 109426 12121 109460 12155
rect 113005 12121 113039 12155
rect 120017 12121 120051 12155
rect 123616 12121 123650 12155
rect 140268 12121 140302 12155
rect 142077 12121 142111 12155
rect 144294 12121 144328 12155
rect 146134 12121 146168 12155
rect 151102 12121 151136 12155
rect 154506 12121 154540 12155
rect 4445 12053 4479 12087
rect 8585 12053 8619 12087
rect 12449 12053 12483 12087
rect 15025 12053 15059 12087
rect 16957 12053 16991 12087
rect 18797 12053 18831 12087
rect 19625 12053 19659 12087
rect 25973 12053 26007 12087
rect 29193 12053 29227 12087
rect 33517 12053 33551 12087
rect 41613 12053 41647 12087
rect 43085 12053 43119 12087
rect 45293 12053 45327 12087
rect 47317 12053 47351 12087
rect 47777 12053 47811 12087
rect 51457 12053 51491 12087
rect 53481 12053 53515 12087
rect 54861 12053 54895 12087
rect 55505 12053 55539 12087
rect 58633 12053 58667 12087
rect 66085 12053 66119 12087
rect 68293 12053 68327 12087
rect 71053 12053 71087 12087
rect 71697 12053 71731 12087
rect 81633 12053 81667 12087
rect 82645 12053 82679 12087
rect 83289 12053 83323 12087
rect 84393 12053 84427 12087
rect 91569 12053 91603 12087
rect 93501 12053 93535 12087
rect 94789 12053 94823 12087
rect 97549 12053 97583 12087
rect 100401 12053 100435 12087
rect 101321 12053 101355 12087
rect 101965 12053 101999 12087
rect 102793 12053 102827 12087
rect 103529 12053 103563 12087
rect 104725 12053 104759 12087
rect 107853 12053 107887 12087
rect 108313 12053 108347 12087
rect 111257 12053 111291 12087
rect 113557 12053 113591 12087
rect 114109 12053 114143 12087
rect 114569 12053 114603 12087
rect 115213 12053 115247 12087
rect 116317 12053 116351 12087
rect 117329 12053 117363 12087
rect 118893 12053 118927 12087
rect 120825 12053 120859 12087
rect 124413 12053 124447 12087
rect 125057 12053 125091 12087
rect 126253 12053 126287 12087
rect 126805 12053 126839 12087
rect 129473 12053 129507 12087
rect 130669 12053 130703 12087
rect 131221 12053 131255 12087
rect 131773 12053 131807 12087
rect 133337 12053 133371 12087
rect 136373 12053 136407 12087
rect 138489 12053 138523 12087
rect 139133 12053 139167 12087
rect 143181 12053 143215 12087
rect 145021 12053 145055 12087
rect 147597 12053 147631 12087
rect 148333 12053 148367 12087
rect 149161 12053 149195 12087
rect 151829 12053 151863 12087
rect 152473 12053 152507 12087
rect 155233 12053 155267 12087
rect 156981 12053 157015 12087
rect 157533 12053 157567 12087
rect 10517 11849 10551 11883
rect 18521 11849 18555 11883
rect 20821 11849 20855 11883
rect 23949 11849 23983 11883
rect 26249 11849 26283 11883
rect 31033 11849 31067 11883
rect 31677 11849 31711 11883
rect 32873 11849 32907 11883
rect 36369 11849 36403 11883
rect 39681 11849 39715 11883
rect 41889 11849 41923 11883
rect 44373 11849 44407 11883
rect 45109 11849 45143 11883
rect 47041 11849 47075 11883
rect 48421 11849 48455 11883
rect 52101 11849 52135 11883
rect 52929 11849 52963 11883
rect 53757 11849 53791 11883
rect 54309 11849 54343 11883
rect 59461 11849 59495 11883
rect 63417 11849 63451 11883
rect 71145 11849 71179 11883
rect 79149 11849 79183 11883
rect 85405 11849 85439 11883
rect 87429 11849 87463 11883
rect 88993 11849 89027 11883
rect 94973 11849 95007 11883
rect 97825 11849 97859 11883
rect 98469 11849 98503 11883
rect 99941 11849 99975 11883
rect 103529 11849 103563 11883
rect 104541 11849 104575 11883
rect 108589 11849 108623 11883
rect 109693 11849 109727 11883
rect 113281 11849 113315 11883
rect 114845 11849 114879 11883
rect 119077 11849 119111 11883
rect 125609 11849 125643 11883
rect 129289 11849 129323 11883
rect 130209 11849 130243 11883
rect 135361 11849 135395 11883
rect 152657 11849 152691 11883
rect 156797 11849 156831 11883
rect 157625 11849 157659 11883
rect 13277 11781 13311 11815
rect 17386 11781 17420 11815
rect 19165 11781 19199 11815
rect 25114 11781 25148 11815
rect 28080 11781 28114 11815
rect 45928 11781 45962 11815
rect 56405 11781 56439 11815
rect 69480 11781 69514 11815
rect 72341 11781 72375 11815
rect 74365 11781 74399 11815
rect 90106 11781 90140 11815
rect 126529 11781 126563 11815
rect 138848 11781 138882 11815
rect 142660 11781 142694 11815
rect 151062 11781 151096 11815
rect 4068 11713 4102 11747
rect 8401 11713 8435 11747
rect 10977 11713 11011 11747
rect 11897 11713 11931 11747
rect 12817 11713 12851 11747
rect 13461 11713 13495 11747
rect 14473 11713 14507 11747
rect 14729 11713 14763 11747
rect 21005 11713 21039 11747
rect 22937 11713 22971 11747
rect 24133 11713 24167 11747
rect 24869 11713 24903 11747
rect 27353 11713 27387 11747
rect 29909 11713 29943 11747
rect 31493 11713 31527 11747
rect 38557 11713 38591 11747
rect 40509 11713 40543 11747
rect 40693 11713 40727 11747
rect 42073 11713 42107 11747
rect 42717 11713 42751 11747
rect 43453 11713 43487 11747
rect 44189 11713 44223 11747
rect 44925 11713 44959 11747
rect 45661 11713 45695 11747
rect 48605 11713 48639 11747
rect 49341 11713 49375 11747
rect 50068 11713 50102 11747
rect 51917 11713 51951 11747
rect 53113 11713 53147 11747
rect 53573 11713 53607 11747
rect 55422 11713 55456 11747
rect 58081 11713 58115 11747
rect 58348 11713 58382 11747
rect 60657 11713 60691 11747
rect 61568 11713 61602 11747
rect 63233 11713 63267 11747
rect 63969 11713 64003 11747
rect 65625 11713 65659 11747
rect 65881 11713 65915 11747
rect 67833 11713 67867 11747
rect 68569 11713 68603 11747
rect 74917 11713 74951 11747
rect 76380 11713 76414 11747
rect 80273 11713 80307 11747
rect 80529 11713 80563 11747
rect 83013 11713 83047 11747
rect 84025 11713 84059 11747
rect 86529 11713 86563 11747
rect 86785 11713 86819 11747
rect 87245 11713 87279 11747
rect 91468 11713 91502 11747
rect 93133 11713 93167 11747
rect 94421 11713 94455 11747
rect 95157 11713 95191 11747
rect 96169 11713 96203 11747
rect 97273 11713 97307 11747
rect 101790 11713 101824 11747
rect 105665 11713 105699 11747
rect 108129 11713 108163 11747
rect 112545 11713 112579 11747
rect 113465 11713 113499 11747
rect 115673 11713 115707 11747
rect 117441 11713 117475 11747
rect 118341 11713 118375 11747
rect 120457 11713 120491 11747
rect 121193 11713 121227 11747
rect 122113 11713 122147 11747
rect 125057 11713 125091 11747
rect 126345 11713 126379 11747
rect 126989 11713 127023 11747
rect 127173 11713 127207 11747
rect 127357 11713 127391 11747
rect 128001 11713 128035 11747
rect 128645 11713 128679 11747
rect 130761 11713 130795 11747
rect 134185 11713 134219 11747
rect 136474 11713 136508 11747
rect 140697 11713 140731 11747
rect 144478 11713 144512 11747
rect 144745 11713 144779 11747
rect 146789 11713 146823 11747
rect 147045 11713 147079 11747
rect 148629 11713 148663 11747
rect 148885 11713 148919 11747
rect 149437 11713 149471 11747
rect 150265 11713 150299 11747
rect 153781 11713 153815 11747
rect 154681 11713 154715 11747
rect 156153 11711 156187 11745
rect 156981 11713 157015 11747
rect 157809 11713 157843 11747
rect 3801 11645 3835 11679
rect 8585 11645 8619 11679
rect 13645 11645 13679 11679
rect 17141 11645 17175 11679
rect 19625 11645 19659 11679
rect 23121 11645 23155 11679
rect 24317 11645 24351 11679
rect 27813 11645 27847 11679
rect 29653 11645 29687 11679
rect 38301 11645 38335 11679
rect 40877 11645 40911 11679
rect 49801 11645 49835 11679
rect 51733 11645 51767 11679
rect 55689 11645 55723 11679
rect 56149 11645 56183 11679
rect 60013 11645 60047 11679
rect 60841 11645 60875 11679
rect 61301 11645 61335 11679
rect 68753 11645 68787 11679
rect 69213 11645 69247 11679
rect 73905 11645 73939 11679
rect 76113 11645 76147 11679
rect 84209 11645 84243 11679
rect 87981 11645 88015 11679
rect 90373 11645 90407 11679
rect 91201 11645 91235 11679
rect 96813 11645 96847 11679
rect 99389 11645 99423 11679
rect 102057 11645 102091 11679
rect 105921 11645 105955 11679
rect 115489 11645 115523 11679
rect 117697 11645 117731 11679
rect 118525 11645 118559 11679
rect 119997 11645 120031 11679
rect 121377 11645 121411 11679
rect 126161 11645 126195 11679
rect 128829 11645 128863 11679
rect 132509 11645 132543 11679
rect 134441 11645 134475 11679
rect 136741 11645 136775 11679
rect 137201 11645 137235 11679
rect 138581 11645 138615 11679
rect 140513 11645 140547 11679
rect 142905 11645 142939 11679
rect 150817 11645 150851 11679
rect 154037 11645 154071 11679
rect 154497 11645 154531 11679
rect 154865 11645 154899 11679
rect 155969 11645 156003 11679
rect 157165 11645 157199 11679
rect 8217 11577 8251 11611
rect 9413 11577 9447 11611
rect 11161 11577 11195 11611
rect 22753 11577 22787 11611
rect 34805 11577 34839 11611
rect 36921 11577 36955 11611
rect 43637 11577 43671 11611
rect 57529 11577 57563 11611
rect 64153 11577 64187 11611
rect 67005 11577 67039 11611
rect 75101 11577 75135 11611
rect 77493 11577 77527 11611
rect 81081 11577 81115 11611
rect 92581 11577 92615 11611
rect 94237 11577 94271 11611
rect 106381 11577 106415 11611
rect 111257 11577 111291 11611
rect 116317 11577 116351 11611
rect 139961 11577 139995 11611
rect 150081 11577 150115 11611
rect 5181 11509 5215 11543
rect 5733 11509 5767 11543
rect 7757 11509 7791 11543
rect 9965 11509 9999 11543
rect 12081 11509 12115 11543
rect 12633 11509 12667 11543
rect 15853 11509 15887 11543
rect 20177 11509 20211 11543
rect 22293 11509 22327 11543
rect 29193 11509 29227 11543
rect 32321 11509 32355 11543
rect 33609 11509 33643 11543
rect 34253 11509 34287 11543
rect 37841 11509 37875 11543
rect 42901 11509 42935 11543
rect 47777 11509 47811 11543
rect 49157 11509 49191 11543
rect 51181 11509 51215 11543
rect 60473 11509 60507 11543
rect 62681 11509 62715 11543
rect 65073 11509 65107 11543
rect 67649 11509 67683 11543
rect 68385 11509 68419 11543
rect 70593 11509 70627 11543
rect 72985 11509 73019 11543
rect 78045 11509 78079 11543
rect 82829 11509 82863 11543
rect 83841 11509 83875 11543
rect 84853 11509 84887 11543
rect 95617 11509 95651 11543
rect 100677 11509 100711 11543
rect 102609 11509 102643 11543
rect 107025 11509 107059 11543
rect 107945 11509 107979 11543
rect 110245 11509 110279 11543
rect 113925 11509 113959 11543
rect 115857 11509 115891 11543
rect 118157 11509 118191 11543
rect 121009 11509 121043 11543
rect 121929 11509 121963 11543
rect 122665 11509 122699 11543
rect 123217 11509 123251 11543
rect 123677 11509 123711 11543
rect 124229 11509 124263 11543
rect 127817 11509 127851 11543
rect 128461 11509 128495 11543
rect 131405 11509 131439 11543
rect 131957 11509 131991 11543
rect 133061 11509 133095 11543
rect 138121 11509 138155 11543
rect 140881 11509 140915 11543
rect 141525 11509 141559 11543
rect 143365 11509 143399 11543
rect 145665 11509 145699 11543
rect 147505 11509 147539 11543
rect 149529 11509 149563 11543
rect 152197 11509 152231 11543
rect 155325 11509 155359 11543
rect 156337 11509 156371 11543
rect 158269 11509 158303 11543
rect 4445 11305 4479 11339
rect 10149 11305 10183 11339
rect 13737 11305 13771 11339
rect 26157 11305 26191 11339
rect 31125 11305 31159 11339
rect 33057 11305 33091 11339
rect 36277 11305 36311 11339
rect 38761 11305 38795 11339
rect 40693 11305 40727 11339
rect 41981 11305 42015 11339
rect 42625 11305 42659 11339
rect 44649 11305 44683 11339
rect 53573 11305 53607 11339
rect 57897 11305 57931 11339
rect 60013 11305 60047 11339
rect 62589 11305 62623 11339
rect 65901 11305 65935 11339
rect 68017 11305 68051 11339
rect 82461 11305 82495 11339
rect 88533 11305 88567 11339
rect 107117 11305 107151 11339
rect 107669 11305 107703 11339
rect 108773 11305 108807 11339
rect 109601 11305 109635 11339
rect 113833 11305 113867 11339
rect 119629 11305 119663 11339
rect 123033 11305 123067 11339
rect 129105 11305 129139 11339
rect 132233 11305 132267 11339
rect 134533 11305 134567 11339
rect 138489 11305 138523 11339
rect 147321 11305 147355 11339
rect 149253 11305 149287 11339
rect 151093 11305 151127 11339
rect 153393 11305 153427 11339
rect 156889 11305 156923 11339
rect 9229 11237 9263 11271
rect 11897 11237 11931 11271
rect 17601 11237 17635 11271
rect 23029 11237 23063 11271
rect 38301 11237 38335 11271
rect 39497 11237 39531 11271
rect 45385 11237 45419 11271
rect 47593 11237 47627 11271
rect 53113 11237 53147 11271
rect 56885 11237 56919 11271
rect 66637 11237 66671 11271
rect 73261 11237 73295 11271
rect 76573 11237 76607 11271
rect 80713 11237 80747 11271
rect 82001 11237 82035 11271
rect 88993 11237 89027 11271
rect 90833 11237 90867 11271
rect 92489 11237 92523 11271
rect 95433 11237 95467 11271
rect 96077 11237 96111 11271
rect 96813 11237 96847 11271
rect 101965 11237 101999 11271
rect 111441 11237 111475 11271
rect 117329 11237 117363 11271
rect 124045 11237 124079 11271
rect 126805 11237 126839 11271
rect 139501 11237 139535 11271
rect 157533 11237 157567 11271
rect 5365 11169 5399 11203
rect 10701 11169 10735 11203
rect 16221 11169 16255 11203
rect 19441 11169 19475 11203
rect 28549 11169 28583 11203
rect 34253 11169 34287 11203
rect 51733 11169 51767 11203
rect 65257 11169 65291 11203
rect 69765 11169 69799 11203
rect 71421 11169 71455 11203
rect 71881 11169 71915 11203
rect 77953 11169 77987 11203
rect 79333 11169 79367 11203
rect 87153 11169 87187 11203
rect 98193 11169 98227 11203
rect 99297 11169 99331 11203
rect 103805 11169 103839 11203
rect 106289 11169 106323 11203
rect 113373 11169 113407 11203
rect 115213 11169 115247 11203
rect 115765 11169 115799 11203
rect 118341 11169 118375 11203
rect 122481 11169 122515 11203
rect 131865 11169 131899 11203
rect 133153 11169 133187 11203
rect 137385 11169 137419 11203
rect 144837 11169 144871 11203
rect 148609 11169 148643 11203
rect 150633 11169 150667 11203
rect 152473 11169 152507 11203
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 5917 11101 5951 11135
rect 11713 11101 11747 11135
rect 12357 11101 12391 11135
rect 14381 11101 14415 11135
rect 16488 11101 16522 11135
rect 18613 11101 18647 11135
rect 21649 11101 21683 11135
rect 23949 11101 23983 11135
rect 26617 11101 26651 11135
rect 26801 11101 26835 11135
rect 29745 11101 29779 11135
rect 30012 11101 30046 11135
rect 31677 11101 31711 11135
rect 33701 11101 33735 11135
rect 34897 11101 34931 11135
rect 35164 11101 35198 11135
rect 36921 11101 36955 11135
rect 37105 11101 37139 11135
rect 39313 11101 39347 11135
rect 40877 11101 40911 11135
rect 41797 11101 41831 11135
rect 42809 11101 42843 11135
rect 43269 11101 43303 11135
rect 45569 11101 45603 11135
rect 45753 11101 45787 11135
rect 46213 11101 46247 11135
rect 48697 11101 48731 11135
rect 49433 11101 49467 11135
rect 49617 11111 49651 11145
rect 50813 11101 50847 11135
rect 50997 11101 51031 11135
rect 54953 11101 54987 11135
rect 55505 11101 55539 11135
rect 55772 11101 55806 11135
rect 57713 11101 57747 11135
rect 58449 11101 58483 11135
rect 58633 11101 58667 11135
rect 58817 11101 58851 11135
rect 59829 11101 59863 11135
rect 60657 11101 60691 11135
rect 62773 11101 62807 11135
rect 66821 11101 66855 11135
rect 69949 11101 69983 11135
rect 70041 11101 70075 11135
rect 72148 11101 72182 11135
rect 75285 11101 75319 11135
rect 78873 11101 78907 11135
rect 81265 11101 81299 11135
rect 83841 11101 83875 11135
rect 84761 11101 84795 11135
rect 85865 11101 85899 11135
rect 86509 11101 86543 11135
rect 90373 11101 90407 11135
rect 93869 11101 93903 11135
rect 94881 11101 94915 11135
rect 98837 11101 98871 11135
rect 103345 11101 103379 11135
rect 108313 11101 108347 11135
rect 108957 11101 108991 11135
rect 109141 11101 109175 11135
rect 110981 11101 111015 11135
rect 111625 11101 111659 11135
rect 117513 11101 117547 11135
rect 118617 11101 118651 11135
rect 120181 11101 120215 11135
rect 120917 11101 120951 11135
rect 121009 11101 121043 11135
rect 121561 11101 121595 11135
rect 125158 11101 125192 11135
rect 125418 11101 125452 11135
rect 126161 11101 126195 11135
rect 126253 11101 126287 11135
rect 127817 11101 127851 11135
rect 128093 11101 128127 11135
rect 130218 11101 130252 11135
rect 130485 11101 130519 11135
rect 132049 11101 132083 11135
rect 141249 11101 141283 11135
rect 141433 11101 141467 11135
rect 142169 11101 142203 11135
rect 142353 11101 142387 11135
rect 146677 11101 146711 11135
rect 147137 11101 147171 11135
rect 148425 11101 148459 11135
rect 154506 11101 154540 11135
rect 154773 11101 154807 11135
rect 155417 11101 155451 11135
rect 155601 11101 155635 11135
rect 156061 11101 156095 11135
rect 156245 11101 156279 11135
rect 157073 11101 157107 11135
rect 157717 11101 157751 11135
rect 7941 11033 7975 11067
rect 11253 11033 11287 11067
rect 12602 11033 12636 11067
rect 14626 11033 14660 11067
rect 21189 11033 21223 11067
rect 21916 11033 21950 11067
rect 25145 11033 25179 11067
rect 25329 11033 25363 11067
rect 26985 11033 27019 11067
rect 31944 11033 31978 11067
rect 36737 11033 36771 11067
rect 37657 11033 37691 11067
rect 40141 11033 40175 11067
rect 43514 11033 43548 11067
rect 46480 11033 46514 11067
rect 51181 11033 51215 11067
rect 52000 11033 52034 11067
rect 54686 11033 54720 11067
rect 60924 11033 60958 11067
rect 64990 11033 65024 11067
rect 69305 11033 69339 11067
rect 74641 11033 74675 11067
rect 77686 11033 77720 11067
rect 79600 11033 79634 11067
rect 83596 11033 83630 11067
rect 85497 11033 85531 11067
rect 87420 11033 87454 11067
rect 90128 11033 90162 11067
rect 91569 11033 91603 11067
rect 93624 11033 93658 11067
rect 94421 11033 94455 11067
rect 97948 11033 97982 11067
rect 99849 11033 99883 11067
rect 103100 11033 103134 11067
rect 104072 11033 104106 11067
rect 105737 11033 105771 11067
rect 110736 11033 110770 11067
rect 112177 11033 112211 11067
rect 112821 11033 112855 11067
rect 114968 11033 115002 11067
rect 120733 11033 120767 11067
rect 125977 11033 126011 11067
rect 131313 11033 131347 11067
rect 133420 11033 133454 11067
rect 135545 11033 135579 11067
rect 136097 11033 136131 11067
rect 136833 11033 136867 11067
rect 139777 11033 139811 11067
rect 140421 11033 140455 11067
rect 141065 11033 141099 11067
rect 141985 11033 142019 11067
rect 144570 11033 144604 11067
rect 146432 11033 146466 11067
rect 148241 11033 148275 11067
rect 150366 11033 150400 11067
rect 152206 11033 152240 11067
rect 155233 11033 155267 11067
rect 156429 11033 156463 11067
rect 15761 10965 15795 10999
rect 18429 10965 18463 10999
rect 27629 10965 27663 10999
rect 29101 10965 29135 10999
rect 33517 10965 33551 10999
rect 48513 10965 48547 10999
rect 49801 10965 49835 10999
rect 59277 10965 59311 10999
rect 62037 10965 62071 10999
rect 63417 10965 63451 10999
rect 63877 10965 63911 10999
rect 74089 10965 74123 10999
rect 75469 10965 75503 10999
rect 84853 10965 84887 10999
rect 98653 10965 98687 10999
rect 105185 10965 105219 10999
rect 116225 10965 116259 10999
rect 121745 10965 121779 10999
rect 134993 10965 135027 10999
rect 143457 10965 143491 10999
rect 145297 10965 145331 10999
rect 5733 10761 5767 10795
rect 11069 10761 11103 10795
rect 13829 10761 13863 10795
rect 15301 10761 15335 10795
rect 18797 10761 18831 10795
rect 19349 10761 19383 10795
rect 19809 10761 19843 10795
rect 22109 10761 22143 10795
rect 24869 10761 24903 10795
rect 26617 10761 26651 10795
rect 27813 10761 27847 10795
rect 36921 10761 36955 10795
rect 37565 10761 37599 10795
rect 40049 10761 40083 10795
rect 45109 10761 45143 10795
rect 45845 10761 45879 10795
rect 49801 10761 49835 10795
rect 51089 10761 51123 10795
rect 55689 10761 55723 10795
rect 57529 10761 57563 10795
rect 60657 10761 60691 10795
rect 81081 10761 81115 10795
rect 87705 10761 87739 10795
rect 89729 10761 89763 10795
rect 93225 10761 93259 10795
rect 100861 10761 100895 10795
rect 103529 10761 103563 10795
rect 106473 10761 106507 10795
rect 108681 10761 108715 10795
rect 112637 10761 112671 10795
rect 113649 10761 113683 10795
rect 114845 10761 114879 10795
rect 115949 10761 115983 10795
rect 117789 10761 117823 10795
rect 125333 10761 125367 10795
rect 126713 10761 126747 10795
rect 130209 10761 130243 10795
rect 136741 10761 136775 10795
rect 139133 10761 139167 10795
rect 140973 10761 141007 10795
rect 148885 10761 148919 10795
rect 150817 10761 150851 10795
rect 155325 10761 155359 10795
rect 157625 10761 157659 10795
rect 158269 10761 158303 10795
rect 4068 10693 4102 10727
rect 12072 10693 12106 10727
rect 17662 10693 17696 10727
rect 25513 10693 25547 10727
rect 38853 10693 38887 10727
rect 61362 10693 61396 10727
rect 68569 10693 68603 10727
rect 72709 10693 72743 10727
rect 79149 10693 79183 10727
rect 79946 10693 79980 10727
rect 86448 10693 86482 10727
rect 101996 10693 102030 10727
rect 102793 10693 102827 10727
rect 104541 10693 104575 10727
rect 117084 10693 117118 10727
rect 131580 10693 131614 10727
rect 141801 10693 141835 10727
rect 144837 10693 144871 10727
rect 145910 10693 145944 10727
rect 8309 10625 8343 10659
rect 9321 10625 9355 10659
rect 11805 10625 11839 10659
rect 13645 10625 13679 10659
rect 14657 10625 14691 10659
rect 15485 10625 15519 10659
rect 16865 10625 16899 10659
rect 17417 10625 17451 10659
rect 28937 10625 28971 10659
rect 29193 10625 29227 10659
rect 30277 10625 30311 10659
rect 32965 10625 32999 10659
rect 33885 10625 33919 10659
rect 35797 10625 35831 10659
rect 40509 10625 40543 10659
rect 41337 10625 41371 10659
rect 41889 10625 41923 10659
rect 43749 10625 43783 10659
rect 44005 10625 44039 10659
rect 44465 10625 44499 10659
rect 45293 10625 45327 10659
rect 46958 10625 46992 10659
rect 47225 10625 47259 10659
rect 47777 10625 47811 10659
rect 48421 10625 48455 10659
rect 48688 10625 48722 10659
rect 50445 10625 50479 10659
rect 50905 10625 50939 10659
rect 51825 10625 51859 10659
rect 51917 10625 51951 10659
rect 54309 10625 54343 10659
rect 54576 10625 54610 10659
rect 56405 10625 56439 10659
rect 58633 10615 58667 10649
rect 58817 10625 58851 10659
rect 59277 10625 59311 10659
rect 59544 10625 59578 10659
rect 61117 10625 61151 10659
rect 63877 10625 63911 10659
rect 64521 10625 64555 10659
rect 66933 10625 66967 10659
rect 69940 10625 69974 10659
rect 72525 10625 72559 10659
rect 73721 10625 73755 10659
rect 73905 10625 73939 10659
rect 75938 10625 75972 10659
rect 76205 10625 76239 10659
rect 76757 10625 76791 10659
rect 77024 10625 77058 10659
rect 82093 10625 82127 10659
rect 82737 10625 82771 10659
rect 86693 10625 86727 10659
rect 89085 10625 89119 10659
rect 89269 10625 89303 10659
rect 91773 10625 91807 10659
rect 102241 10625 102275 10659
rect 103345 10625 103379 10659
rect 105093 10625 105127 10659
rect 105360 10625 105394 10659
rect 107025 10625 107059 10659
rect 107761 10625 107795 10659
rect 107945 10625 107979 10659
rect 110613 10625 110647 10659
rect 111441 10625 111475 10659
rect 111533 10625 111567 10659
rect 113833 10625 113867 10659
rect 118913 10625 118947 10659
rect 120549 10625 120583 10659
rect 122122 10625 122156 10659
rect 123033 10625 123067 10659
rect 124229 10625 124263 10659
rect 125885 10625 125919 10659
rect 126069 10625 126103 10659
rect 126897 10625 126931 10659
rect 128001 10625 128035 10659
rect 128553 10625 128587 10659
rect 128829 10625 128863 10659
rect 130853 10625 130887 10659
rect 138417 10625 138451 10659
rect 138673 10625 138707 10659
rect 141157 10625 141191 10659
rect 144009 10625 144043 10659
rect 144193 10625 144227 10659
rect 145665 10625 145699 10659
rect 147772 10625 147806 10659
rect 149437 10625 149471 10659
rect 149621 10625 149655 10659
rect 150265 10625 150299 10659
rect 151930 10625 151964 10659
rect 152197 10625 152231 10659
rect 153770 10625 153804 10659
rect 154681 10625 154715 10659
rect 155969 10625 156003 10659
rect 156153 10625 156187 10659
rect 156981 10625 157015 10659
rect 157809 10625 157843 10659
rect 3801 10557 3835 10591
rect 9137 10557 9171 10591
rect 23029 10557 23063 10591
rect 30021 10557 30055 10591
rect 33701 10557 33735 10591
rect 34989 10557 35023 10591
rect 35541 10557 35575 10591
rect 52929 10557 52963 10591
rect 53205 10557 53239 10591
rect 56149 10557 56183 10591
rect 63693 10557 63727 10591
rect 67189 10557 67223 10591
rect 69673 10557 69707 10591
rect 72341 10557 72375 10591
rect 73537 10557 73571 10591
rect 79701 10557 79735 10591
rect 82553 10557 82587 10591
rect 92029 10557 92063 10591
rect 109693 10557 109727 10591
rect 110429 10557 110463 10591
rect 117329 10557 117363 10591
rect 119169 10557 119203 10591
rect 122389 10557 122423 10591
rect 131313 10557 131347 10591
rect 139685 10557 139719 10591
rect 144377 10557 144411 10591
rect 147505 10557 147539 10591
rect 154037 10557 154071 10591
rect 154865 10557 154899 10591
rect 156797 10557 156831 10591
rect 13185 10489 13219 10523
rect 14841 10489 14875 10523
rect 31401 10489 31435 10523
rect 32413 10489 32447 10523
rect 41153 10489 41187 10523
rect 50261 10489 50295 10523
rect 51641 10489 51675 10523
rect 62497 10489 62531 10523
rect 65809 10489 65843 10523
rect 71053 10489 71087 10523
rect 78137 10489 78171 10523
rect 87245 10489 87279 10523
rect 90649 10489 90683 10523
rect 127817 10489 127851 10523
rect 133245 10489 133279 10523
rect 135637 10489 135671 10523
rect 152657 10489 152691 10523
rect 156337 10489 156371 10523
rect 5181 10421 5215 10455
rect 8125 10421 8159 10455
rect 9505 10421 9539 10455
rect 10057 10421 10091 10455
rect 16129 10421 16163 10455
rect 21373 10421 21407 10455
rect 23765 10421 23799 10455
rect 25973 10421 26007 10455
rect 27261 10421 27295 10455
rect 33149 10421 33183 10455
rect 34069 10421 34103 10455
rect 39405 10421 39439 10455
rect 40693 10421 40727 10455
rect 41981 10421 42015 10455
rect 42625 10421 42659 10455
rect 47961 10421 47995 10455
rect 58449 10421 58483 10455
rect 64061 10421 64095 10455
rect 64705 10421 64739 10455
rect 65257 10421 65291 10455
rect 67833 10421 67867 10455
rect 69121 10421 69155 10455
rect 71789 10421 71823 10455
rect 74825 10421 74859 10455
rect 81909 10421 81943 10455
rect 82921 10421 82955 10455
rect 85313 10421 85347 10455
rect 88441 10421 88475 10455
rect 92765 10421 92799 10455
rect 94329 10421 94363 10455
rect 94881 10421 94915 10455
rect 95433 10421 95467 10455
rect 95985 10421 96019 10455
rect 96721 10421 96755 10455
rect 98285 10421 98319 10455
rect 108129 10421 108163 10455
rect 110797 10421 110831 10455
rect 111257 10421 111291 10455
rect 112177 10421 112211 10455
rect 115305 10421 115339 10455
rect 120365 10421 120399 10455
rect 121009 10421 121043 10455
rect 122941 10421 122975 10455
rect 123677 10421 123711 10455
rect 126253 10421 126287 10455
rect 132693 10421 132727 10455
rect 133705 10421 133739 10455
rect 134809 10421 134843 10455
rect 136189 10421 136223 10455
rect 137293 10421 137327 10455
rect 143089 10421 143123 10455
rect 147045 10421 147079 10455
rect 150081 10421 150115 10455
rect 154497 10421 154531 10455
rect 157165 10421 157199 10455
rect 1961 10217 1995 10251
rect 5825 10217 5859 10251
rect 25421 10217 25455 10251
rect 29193 10217 29227 10251
rect 40325 10217 40359 10251
rect 41429 10217 41463 10251
rect 44649 10217 44683 10251
rect 46121 10217 46155 10251
rect 47869 10217 47903 10251
rect 50445 10217 50479 10251
rect 51273 10217 51307 10251
rect 52193 10217 52227 10251
rect 82645 10217 82679 10251
rect 96813 10217 96847 10251
rect 100769 10217 100803 10251
rect 101321 10217 101355 10251
rect 104357 10217 104391 10251
rect 107117 10217 107151 10251
rect 107669 10217 107703 10251
rect 112545 10217 112579 10251
rect 137385 10217 137419 10251
rect 147045 10217 147079 10251
rect 157349 10217 157383 10251
rect 12633 10149 12667 10183
rect 15669 10149 15703 10183
rect 37657 10149 37691 10183
rect 54033 10149 54067 10183
rect 55597 10149 55631 10183
rect 56241 10149 56275 10183
rect 57897 10149 57931 10183
rect 59001 10149 59035 10183
rect 60013 10149 60047 10183
rect 62037 10149 62071 10183
rect 75101 10149 75135 10183
rect 77309 10149 77343 10183
rect 84853 10149 84887 10183
rect 85589 10149 85623 10183
rect 89729 10149 89763 10183
rect 90833 10149 90867 10183
rect 92857 10149 92891 10183
rect 98837 10149 98871 10183
rect 101873 10149 101907 10183
rect 109785 10149 109819 10183
rect 118709 10149 118743 10183
rect 120549 10149 120583 10183
rect 121469 10149 121503 10183
rect 123217 10149 123251 10183
rect 128369 10149 128403 10183
rect 148241 10149 148275 10183
rect 153853 10149 153887 10183
rect 25973 10081 26007 10115
rect 27813 10081 27847 10115
rect 38853 10081 38887 10115
rect 45569 10081 45603 10115
rect 52653 10081 52687 10115
rect 54493 10081 54527 10115
rect 60657 10081 60691 10115
rect 65257 10081 65291 10115
rect 67189 10081 67223 10115
rect 100217 10081 100251 10115
rect 103253 10081 103287 10115
rect 127725 10081 127759 10115
rect 132785 10081 132819 10115
rect 145205 10081 145239 10115
rect 149621 10081 149655 10115
rect 151921 10081 151955 10115
rect 155693 10081 155727 10115
rect 156061 10081 156095 10115
rect 3985 10013 4019 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 13093 10013 13127 10047
rect 14289 10013 14323 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 17325 10013 17359 10047
rect 19441 10013 19475 10047
rect 31217 10013 31251 10047
rect 31861 10013 31895 10047
rect 32781 10013 32815 10047
rect 33425 10013 33459 10047
rect 33517 10013 33551 10047
rect 33701 10013 33735 10047
rect 36277 10013 36311 10047
rect 38117 10013 38151 10047
rect 40785 10013 40819 10047
rect 42542 10013 42576 10047
rect 42809 10013 42843 10047
rect 43269 10013 43303 10047
rect 43536 10013 43570 10047
rect 46305 10013 46339 10047
rect 46949 10013 46983 10047
rect 47133 10013 47167 10047
rect 47685 10013 47719 10047
rect 49801 10013 49835 10047
rect 50629 10013 50663 10047
rect 51089 10013 51123 10047
rect 51825 10013 51859 10047
rect 52009 10013 52043 10047
rect 54677 10013 54711 10047
rect 56057 10013 56091 10047
rect 56793 10013 56827 10047
rect 56977 10013 57011 10047
rect 58817 10013 58851 10047
rect 59829 10013 59863 10047
rect 63049 10013 63083 10047
rect 63233 10013 63267 10047
rect 71237 10013 71271 10047
rect 73721 10013 73755 10047
rect 76297 10013 76331 10047
rect 76389 10013 76423 10047
rect 78321 10013 78355 10047
rect 80713 10013 80747 10047
rect 81265 10013 81299 10047
rect 84217 10013 84251 10047
rect 85405 10013 85439 10047
rect 89269 10013 89303 10047
rect 91661 10013 91695 10047
rect 94237 10013 94271 10047
rect 94789 10013 94823 10047
rect 95056 10013 95090 10047
rect 96997 10013 97031 10047
rect 97089 10013 97123 10047
rect 97825 10013 97859 10047
rect 108405 10013 108439 10047
rect 110245 10013 110279 10047
rect 111349 10013 111383 10047
rect 114385 10013 114419 10047
rect 114569 10013 114603 10047
rect 115673 10013 115707 10047
rect 116133 10013 116167 10047
rect 116317 10013 116351 10047
rect 117329 10013 117363 10047
rect 119169 10013 119203 10047
rect 119905 10013 119939 10047
rect 121101 10013 121135 10047
rect 121271 10013 121305 10047
rect 122665 10013 122699 10047
rect 125149 10013 125183 10047
rect 129749 10013 129783 10047
rect 130025 10013 130059 10047
rect 130485 10013 130519 10047
rect 130761 10013 130795 10047
rect 132969 10013 133003 10047
rect 135545 10013 135579 10047
rect 136005 10013 136039 10047
rect 138857 10013 138891 10047
rect 140605 10013 140639 10047
rect 142537 10013 142571 10047
rect 143365 10013 143399 10047
rect 145472 10013 145506 10047
rect 147597 10013 147631 10047
rect 149354 10013 149388 10047
rect 151461 10013 151495 10047
rect 152105 10013 152139 10047
rect 152289 10013 152323 10047
rect 154977 10013 155011 10047
rect 155233 10013 155267 10047
rect 155877 10013 155911 10047
rect 156613 10013 156647 10047
rect 156705 10013 156739 10047
rect 157533 10013 157567 10047
rect 1685 9945 1719 9979
rect 4252 9945 4286 9979
rect 10333 9945 10367 9979
rect 10977 9945 11011 9979
rect 14534 9945 14568 9979
rect 16221 9945 16255 9979
rect 26218 9945 26252 9979
rect 28080 9945 28114 9979
rect 30972 9945 31006 9979
rect 36544 9945 36578 9979
rect 49534 9945 49568 9979
rect 52920 9945 52954 9979
rect 57713 9945 57747 9979
rect 60924 9945 60958 9979
rect 64990 9945 65024 9979
rect 66922 9945 66956 9979
rect 73988 9945 74022 9979
rect 78588 9945 78622 9979
rect 81532 9945 81566 9979
rect 87337 9945 87371 9979
rect 89002 9945 89036 9979
rect 92213 9945 92247 9979
rect 93970 9945 94004 9979
rect 99972 9945 100006 9979
rect 103008 9945 103042 9979
rect 108672 9945 108706 9979
rect 117596 9945 117630 9979
rect 123861 9945 123895 9979
rect 125416 9945 125450 9979
rect 126989 9945 127023 9979
rect 132141 9945 132175 9979
rect 135300 9945 135334 9979
rect 136272 9945 136306 9979
rect 138121 9945 138155 9979
rect 139317 9945 139351 9979
rect 142292 9945 142326 9979
rect 143632 9945 143666 9979
rect 151194 9945 151228 9979
rect 5365 9877 5399 9911
rect 8401 9877 8435 9911
rect 11805 9877 11839 9911
rect 13277 9877 13311 9911
rect 17141 9877 17175 9911
rect 17877 9877 17911 9911
rect 18429 9877 18463 9911
rect 19625 9877 19659 9911
rect 20085 9877 20119 9911
rect 27353 9877 27387 9911
rect 29837 9877 29871 9911
rect 32045 9877 32079 9911
rect 32597 9877 32631 9911
rect 34161 9877 34195 9911
rect 34989 9877 35023 9911
rect 35817 9877 35851 9911
rect 39405 9877 39439 9911
rect 40969 9877 41003 9911
rect 46765 9877 46799 9911
rect 48421 9877 48455 9911
rect 54861 9877 54895 9911
rect 57161 9877 57195 9911
rect 62497 9877 62531 9911
rect 63417 9877 63451 9911
rect 63877 9877 63911 9911
rect 65809 9877 65843 9911
rect 69581 9877 69615 9911
rect 72617 9877 72651 9911
rect 73169 9877 73203 9911
rect 76113 9877 76147 9911
rect 77861 9877 77895 9911
rect 79701 9877 79735 9911
rect 83105 9877 83139 9911
rect 84025 9877 84059 9911
rect 87889 9877 87923 9911
rect 90373 9877 90407 9911
rect 96169 9877 96203 9911
rect 98009 9877 98043 9911
rect 103805 9877 103839 9911
rect 104817 9877 104851 9911
rect 110889 9877 110923 9911
rect 113097 9877 113131 9911
rect 113649 9877 113683 9911
rect 114201 9877 114235 9911
rect 115489 9877 115523 9911
rect 116501 9877 116535 9911
rect 119353 9877 119387 9911
rect 122481 9877 122515 9911
rect 124413 9877 124447 9911
rect 126529 9877 126563 9911
rect 133521 9877 133555 9911
rect 134165 9877 134199 9911
rect 138213 9877 138247 9911
rect 139961 9877 139995 9911
rect 140421 9877 140455 9911
rect 141157 9877 141191 9911
rect 144745 9877 144779 9911
rect 146585 9877 146619 9911
rect 150081 9877 150115 9911
rect 152749 9877 152783 9911
rect 156889 9877 156923 9911
rect 1593 9673 1627 9707
rect 5733 9673 5767 9707
rect 31677 9673 31711 9707
rect 35817 9673 35851 9707
rect 36829 9673 36863 9707
rect 47225 9673 47259 9707
rect 55965 9673 55999 9707
rect 56793 9673 56827 9707
rect 65533 9673 65567 9707
rect 88349 9673 88383 9707
rect 96353 9673 96387 9707
rect 117421 9673 117455 9707
rect 132601 9673 132635 9707
rect 149805 9673 149839 9707
rect 151277 9673 151311 9707
rect 158269 9673 158303 9707
rect 11989 9605 12023 9639
rect 15393 9605 15427 9639
rect 21097 9605 21131 9639
rect 28374 9605 28408 9639
rect 30941 9605 30975 9639
rect 39589 9605 39623 9639
rect 40233 9605 40267 9639
rect 40960 9605 40994 9639
rect 43422 9605 43456 9639
rect 49341 9605 49375 9639
rect 62221 9605 62255 9639
rect 66729 9605 66763 9639
rect 72893 9605 72927 9639
rect 74733 9605 74767 9639
rect 77677 9605 77711 9639
rect 84954 9605 84988 9639
rect 85773 9605 85807 9639
rect 92038 9605 92072 9639
rect 93593 9605 93627 9639
rect 95534 9605 95568 9639
rect 98745 9605 98779 9639
rect 116602 9605 116636 9639
rect 130301 9605 130335 9639
rect 136833 9605 136867 9639
rect 153945 9605 153979 9639
rect 3801 9537 3835 9571
rect 4068 9537 4102 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 13820 9537 13854 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 17233 9537 17267 9571
rect 19001 9537 19035 9571
rect 19257 9537 19291 9571
rect 19717 9537 19751 9571
rect 19901 9537 19935 9571
rect 26085 9537 26119 9571
rect 29368 9537 29402 9571
rect 31493 9537 31527 9571
rect 32689 9537 32723 9571
rect 32956 9537 32990 9571
rect 34529 9537 34563 9571
rect 38689 9537 38723 9571
rect 38945 9537 38979 9571
rect 40693 9537 40727 9571
rect 45017 9537 45051 9571
rect 46857 9537 46891 9571
rect 47041 9537 47075 9571
rect 48237 9537 48271 9571
rect 48421 9537 48455 9571
rect 49157 9537 49191 9571
rect 50261 9537 50295 9571
rect 50528 9537 50562 9571
rect 52929 9537 52963 9571
rect 53196 9537 53230 9571
rect 55137 9537 55171 9571
rect 56149 9537 56183 9571
rect 56609 9537 56643 9571
rect 57529 9537 57563 9571
rect 58265 9537 58299 9571
rect 60482 9537 60516 9571
rect 60749 9537 60783 9571
rect 63601 9537 63635 9571
rect 64705 9537 64739 9571
rect 64889 9537 64923 9571
rect 64981 9537 65015 9571
rect 67649 9537 67683 9571
rect 73721 9537 73755 9571
rect 76306 9537 76340 9571
rect 77033 9537 77067 9571
rect 83197 9537 83231 9571
rect 85221 9537 85255 9571
rect 89085 9537 89119 9571
rect 89341 9537 89375 9571
rect 95801 9537 95835 9571
rect 98561 9537 98595 9571
rect 99564 9537 99598 9571
rect 104449 9537 104483 9571
rect 104633 9537 104667 9571
rect 105645 9537 105679 9571
rect 108405 9537 108439 9571
rect 111533 9537 111567 9571
rect 113465 9537 113499 9571
rect 121009 9537 121043 9571
rect 121837 9537 121871 9571
rect 122104 9537 122138 9571
rect 123677 9537 123711 9571
rect 124413 9537 124447 9571
rect 125517 9537 125551 9571
rect 129401 9537 129435 9571
rect 129657 9537 129691 9571
rect 131221 9537 131255 9571
rect 131477 9537 131511 9571
rect 133685 9537 133719 9571
rect 138193 9537 138227 9571
rect 140973 9537 141007 9571
rect 141157 9537 141191 9571
rect 143017 9537 143051 9571
rect 143273 9537 143307 9571
rect 144857 9537 144891 9571
rect 146881 9537 146915 9571
rect 147853 9537 147887 9571
rect 149437 9537 149471 9571
rect 149621 9537 149655 9571
rect 152401 9537 152435 9571
rect 153301 9537 153335 9571
rect 154143 9535 154177 9569
rect 154957 9537 154991 9571
rect 155049 9537 155083 9571
rect 156153 9537 156187 9571
rect 156981 9537 157015 9571
rect 157809 9537 157843 9571
rect 16221 9469 16255 9503
rect 17049 9469 17083 9503
rect 20085 9469 20119 9503
rect 26341 9469 26375 9503
rect 28641 9469 28675 9503
rect 29101 9469 29135 9503
rect 43177 9469 43211 9503
rect 73905 9469 73939 9503
rect 76573 9469 76607 9503
rect 92305 9469 92339 9503
rect 98377 9469 98411 9503
rect 99297 9469 99331 9503
rect 112729 9469 112763 9503
rect 113281 9469 113315 9503
rect 114753 9469 114787 9503
rect 116869 9469 116903 9503
rect 118341 9469 118375 9503
rect 125701 9469 125735 9503
rect 133429 9469 133463 9503
rect 137937 9469 137971 9503
rect 145113 9469 145147 9503
rect 147137 9469 147171 9503
rect 147597 9469 147631 9503
rect 152657 9469 152691 9503
rect 153485 9469 153519 9503
rect 154313 9469 154347 9503
rect 155969 9469 156003 9503
rect 156797 9469 156831 9503
rect 14933 9401 14967 9435
rect 27261 9401 27295 9435
rect 30481 9401 30515 9435
rect 37565 9401 37599 9435
rect 42073 9401 42107 9435
rect 51641 9401 51675 9435
rect 55321 9401 55355 9435
rect 58449 9401 58483 9435
rect 75193 9401 75227 9435
rect 77217 9401 77251 9435
rect 83841 9401 83875 9435
rect 90925 9401 90959 9435
rect 101229 9401 101263 9435
rect 108589 9401 108623 9435
rect 113649 9401 113683 9435
rect 123217 9401 123251 9435
rect 125333 9401 125367 9435
rect 127725 9401 127759 9435
rect 135729 9401 135763 9435
rect 136373 9401 136407 9435
rect 139317 9401 139351 9435
rect 5181 9333 5215 9367
rect 12725 9333 12759 9367
rect 17417 9333 17451 9367
rect 17877 9333 17911 9367
rect 20637 9333 20671 9367
rect 24961 9333 24995 9367
rect 34069 9333 34103 9367
rect 42717 9333 42751 9367
rect 44557 9333 44591 9367
rect 45201 9333 45235 9367
rect 45753 9333 45787 9367
rect 46305 9333 46339 9367
rect 48605 9333 48639 9367
rect 52285 9333 52319 9367
rect 54309 9333 54343 9367
rect 57345 9333 57379 9367
rect 59369 9333 59403 9367
rect 61669 9333 61703 9367
rect 63785 9333 63819 9367
rect 66085 9333 66119 9367
rect 67465 9333 67499 9367
rect 73537 9333 73571 9367
rect 79885 9333 79919 9367
rect 90465 9333 90499 9367
rect 94421 9333 94455 9367
rect 97825 9333 97859 9367
rect 100677 9333 100711 9367
rect 103437 9333 103471 9367
rect 104817 9333 104851 9367
rect 105461 9333 105495 9367
rect 107209 9333 107243 9367
rect 110061 9333 110095 9367
rect 111349 9333 111383 9367
rect 114109 9333 114143 9367
rect 115489 9333 115523 9367
rect 118801 9333 118835 9367
rect 119905 9333 119939 9367
rect 126161 9333 126195 9367
rect 126713 9333 126747 9367
rect 128277 9333 128311 9367
rect 134809 9333 134843 9367
rect 137385 9333 137419 9367
rect 139869 9333 139903 9367
rect 140789 9333 140823 9367
rect 141893 9333 141927 9367
rect 143733 9333 143767 9367
rect 145757 9333 145791 9367
rect 148977 9333 149011 9367
rect 153117 9333 153151 9367
rect 154773 9333 154807 9367
rect 156337 9333 156371 9367
rect 157165 9333 157199 9367
rect 157625 9333 157659 9367
rect 3985 9129 4019 9163
rect 13737 9129 13771 9163
rect 21373 9129 21407 9163
rect 26433 9129 26467 9163
rect 39405 9129 39439 9163
rect 43913 9129 43947 9163
rect 48697 9129 48731 9163
rect 53389 9129 53423 9163
rect 55689 9129 55723 9163
rect 57069 9129 57103 9163
rect 64521 9129 64555 9163
rect 65165 9129 65199 9163
rect 67189 9129 67223 9163
rect 74457 9129 74491 9163
rect 87797 9129 87831 9163
rect 88809 9129 88843 9163
rect 101229 9129 101263 9163
rect 114937 9129 114971 9163
rect 115489 9129 115523 9163
rect 117973 9129 118007 9163
rect 131681 9129 131715 9163
rect 148793 9129 148827 9163
rect 155417 9129 155451 9163
rect 10701 9061 10735 9095
rect 18613 9061 18647 9095
rect 29193 9061 29227 9095
rect 33149 9061 33183 9095
rect 47225 9061 47259 9095
rect 49801 9061 49835 9095
rect 59093 9061 59127 9095
rect 94789 9061 94823 9095
rect 96721 9061 96755 9095
rect 98561 9061 98595 9095
rect 104909 9061 104943 9095
rect 126989 9061 127023 9095
rect 130577 9061 130611 9095
rect 131129 9061 131163 9095
rect 138121 9061 138155 9095
rect 138673 9061 138707 9095
rect 139317 9061 139351 9095
rect 139869 9061 139903 9095
rect 144929 9061 144963 9095
rect 145665 9061 145699 9095
rect 153761 9061 153795 9095
rect 157533 9061 157567 9095
rect 11253 8993 11287 9027
rect 14289 8993 14323 9027
rect 15117 8993 15151 9027
rect 16957 8993 16991 9027
rect 19441 8993 19475 9027
rect 27813 8993 27847 9027
rect 31769 8993 31803 9027
rect 33977 8993 34011 9027
rect 36737 8993 36771 9027
rect 37197 8993 37231 9027
rect 41797 8993 41831 9027
rect 50721 8993 50755 9027
rect 62129 8993 62163 9027
rect 90833 8993 90867 9027
rect 92949 8993 92983 9027
rect 93409 8993 93443 9027
rect 96077 8993 96111 9027
rect 100769 8993 100803 9027
rect 124781 8993 124815 9027
rect 126621 8993 126655 9027
rect 129197 8993 129231 9027
rect 147045 8993 147079 9027
rect 150633 8993 150667 9027
rect 5365 8925 5399 8959
rect 5825 8925 5859 8959
rect 11437 8925 11471 8959
rect 12357 8925 12391 8959
rect 14473 8925 14507 8959
rect 17141 8925 17175 8959
rect 17785 8925 17819 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 27169 8925 27203 8959
rect 29745 8925 29779 8959
rect 33793 8925 33827 8959
rect 42533 8925 42567 8959
rect 45201 8925 45235 8959
rect 45845 8925 45879 8959
rect 53573 8925 53607 8959
rect 54309 8925 54343 8959
rect 54493 8925 54527 8959
rect 56241 8925 56275 8959
rect 57253 8925 57287 8959
rect 57713 8925 57747 8959
rect 57980 8925 58014 8959
rect 65809 8925 65843 8959
rect 66065 8925 66099 8959
rect 68109 8925 68143 8959
rect 68845 8925 68879 8959
rect 75101 8925 75135 8959
rect 76297 8925 76331 8959
rect 76481 8925 76515 8959
rect 76941 8925 76975 8959
rect 86417 8925 86451 8959
rect 90566 8925 90600 8959
rect 98101 8925 98135 8959
rect 100502 8925 100536 8959
rect 107393 8925 107427 8959
rect 107577 8925 107611 8959
rect 107761 8925 107795 8959
rect 108405 8925 108439 8959
rect 111073 8925 111107 8959
rect 112361 8925 112395 8959
rect 118157 8925 118191 8959
rect 119629 8925 119663 8959
rect 121837 8925 121871 8959
rect 122665 8925 122699 8959
rect 122849 8925 122883 8959
rect 126805 8925 126839 8959
rect 127633 8925 127667 8959
rect 132969 8925 133003 8959
rect 133153 8925 133187 8959
rect 135637 8925 135671 8959
rect 137937 8925 137971 8959
rect 140329 8925 140363 8959
rect 140973 8925 141007 8959
rect 141709 8925 141743 8959
rect 141985 8925 142019 8959
rect 144213 8925 144247 8959
rect 144469 8925 144503 8959
rect 150173 8925 150207 8959
rect 150817 8925 150851 8959
rect 151553 8925 151587 8959
rect 151645 8925 151679 8959
rect 151829 8925 151863 8959
rect 152473 8925 152507 8959
rect 152565 8925 152599 8959
rect 153485 8925 153519 8959
rect 153577 8925 153611 8959
rect 154221 8925 154255 8959
rect 154405 8925 154439 8959
rect 155141 8925 155175 8959
rect 155233 8925 155267 8959
rect 156061 8925 156095 8959
rect 156153 8925 156187 8959
rect 156705 8925 156739 8959
rect 156889 8925 156923 8959
rect 157717 8925 157751 8959
rect 5120 8857 5154 8891
rect 12602 8857 12636 8891
rect 15384 8857 15418 8891
rect 19686 8857 19720 8891
rect 28058 8857 28092 8891
rect 29990 8857 30024 8891
rect 32036 8857 32070 8891
rect 36492 8857 36526 8891
rect 37464 8857 37498 8891
rect 41530 8857 41564 8891
rect 42778 8857 42812 8891
rect 46090 8857 46124 8891
rect 50966 8857 51000 8891
rect 60841 8857 60875 8891
rect 62396 8857 62430 8891
rect 86684 8857 86718 8891
rect 92682 8857 92716 8891
rect 93676 8857 93710 8891
rect 97834 8857 97868 8891
rect 104265 8857 104299 8891
rect 116777 8857 116811 8891
rect 119445 8857 119479 8891
rect 128737 8857 128771 8891
rect 129442 8857 129476 8891
rect 132141 8857 132175 8891
rect 146800 8857 146834 8891
rect 149928 8857 149962 8891
rect 152289 8857 152323 8891
rect 154589 8857 154623 8891
rect 11621 8789 11655 8823
rect 14657 8789 14691 8823
rect 16497 8789 16531 8823
rect 17325 8789 17359 8823
rect 20821 8789 20855 8823
rect 27353 8789 27387 8823
rect 31125 8789 31159 8823
rect 33609 8789 33643 8823
rect 35357 8789 35391 8823
rect 38577 8789 38611 8823
rect 40417 8789 40451 8823
rect 44649 8789 44683 8823
rect 45385 8789 45419 8823
rect 48053 8789 48087 8823
rect 49249 8789 49283 8823
rect 52101 8789 52135 8823
rect 52837 8789 52871 8823
rect 54677 8789 54711 8823
rect 56425 8789 56459 8823
rect 59553 8789 59587 8823
rect 61669 8789 61703 8823
rect 63509 8789 63543 8823
rect 68293 8789 68327 8823
rect 74917 8789 74951 8823
rect 76113 8789 76147 8823
rect 88349 8789 88383 8823
rect 89453 8789 89487 8823
rect 91569 8789 91603 8823
rect 99389 8789 99423 8823
rect 108221 8789 108255 8823
rect 110889 8789 110923 8823
rect 112545 8789 112579 8823
rect 113097 8789 113131 8823
rect 115949 8789 115983 8823
rect 117329 8789 117363 8823
rect 118709 8789 118743 8823
rect 120181 8789 120215 8823
rect 120733 8789 120767 8823
rect 121377 8789 121411 8823
rect 122481 8789 122515 8823
rect 123401 8789 123435 8823
rect 124229 8789 124263 8823
rect 125241 8789 125275 8823
rect 125885 8789 125919 8823
rect 132785 8789 132819 8823
rect 133613 8789 133647 8823
rect 134165 8789 134199 8823
rect 135177 8789 135211 8823
rect 135821 8789 135855 8823
rect 136465 8789 136499 8823
rect 137293 8789 137327 8823
rect 140513 8789 140547 8823
rect 141157 8789 141191 8823
rect 143089 8789 143123 8823
rect 147505 8789 147539 8823
rect 148333 8789 148367 8823
rect 151001 8789 151035 8823
rect 155877 8789 155911 8823
rect 157073 8789 157107 8823
rect 5181 8585 5215 8619
rect 11805 8585 11839 8619
rect 18429 8585 18463 8619
rect 19441 8585 19475 8619
rect 28549 8585 28583 8619
rect 29561 8585 29595 8619
rect 33333 8585 33367 8619
rect 35909 8585 35943 8619
rect 45293 8585 45327 8619
rect 48789 8585 48823 8619
rect 49433 8585 49467 8619
rect 51457 8585 51491 8619
rect 53481 8585 53515 8619
rect 56057 8585 56091 8619
rect 60013 8585 60047 8619
rect 61393 8585 61427 8619
rect 62681 8585 62715 8619
rect 63785 8585 63819 8619
rect 67465 8585 67499 8619
rect 69765 8585 69799 8619
rect 88993 8585 89027 8619
rect 117421 8585 117455 8619
rect 122389 8585 122423 8619
rect 130577 8585 130611 8619
rect 131589 8585 131623 8619
rect 135729 8585 135763 8619
rect 145021 8585 145055 8619
rect 149713 8585 149747 8619
rect 150817 8585 150851 8619
rect 155325 8585 155359 8619
rect 13470 8517 13504 8551
rect 29009 8517 29043 8551
rect 30113 8517 30147 8551
rect 38936 8517 38970 8551
rect 40693 8517 40727 8551
rect 46406 8517 46440 8551
rect 55054 8517 55088 8551
rect 58348 8517 58382 8551
rect 64245 8517 64279 8551
rect 87898 8517 87932 8551
rect 112177 8517 112211 8551
rect 115305 8517 115339 8551
rect 120724 8517 120758 8551
rect 133674 8517 133708 8551
rect 4537 8449 4571 8483
rect 6009 8449 6043 8483
rect 6745 8449 6779 8483
rect 13737 8449 13771 8483
rect 14657 8449 14691 8483
rect 14924 8449 14958 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 27169 8449 27203 8483
rect 27425 8449 27459 8483
rect 30852 8439 30886 8473
rect 33517 8449 33551 8483
rect 35090 8449 35124 8483
rect 35357 8449 35391 8483
rect 36553 8449 36587 8483
rect 36737 8449 36771 8483
rect 37841 8449 37875 8483
rect 38025 8449 38059 8483
rect 38669 8449 38703 8483
rect 41245 8449 41279 8483
rect 41429 8449 41463 8483
rect 41521 8449 41555 8483
rect 43749 8449 43783 8483
rect 44649 8449 44683 8483
rect 48329 8449 48363 8483
rect 48973 8449 49007 8483
rect 50546 8449 50580 8483
rect 52193 8449 52227 8483
rect 52285 8449 52319 8483
rect 55321 8449 55355 8483
rect 56701 8449 56735 8483
rect 57161 8449 57195 8483
rect 57345 8449 57379 8483
rect 60657 8449 60691 8483
rect 60749 8449 60783 8483
rect 67649 8449 67683 8483
rect 68652 8449 68686 8483
rect 70225 8449 70259 8483
rect 76030 8449 76064 8483
rect 76297 8449 76331 8483
rect 76757 8449 76791 8483
rect 77024 8449 77058 8483
rect 83841 8449 83875 8483
rect 88165 8449 88199 8483
rect 90106 8449 90140 8483
rect 91946 8449 91980 8483
rect 92206 8449 92240 8483
rect 94329 8449 94363 8483
rect 98193 8449 98227 8483
rect 107025 8449 107059 8483
rect 108313 8449 108347 8483
rect 108957 8449 108991 8483
rect 109601 8449 109635 8483
rect 109868 8449 109902 8483
rect 112821 8449 112855 8483
rect 118157 8449 118191 8483
rect 118985 8449 119019 8483
rect 122573 8449 122607 8483
rect 123300 8449 123334 8483
rect 126529 8449 126563 8483
rect 127265 8449 127299 8483
rect 128553 8449 128587 8483
rect 130393 8449 130427 8483
rect 132713 8449 132747 8483
rect 137477 8449 137511 8483
rect 140513 8449 140547 8483
rect 141341 8449 141375 8483
rect 142914 8449 142948 8483
rect 143181 8449 143215 8483
rect 143641 8449 143675 8483
rect 143908 8449 143942 8483
rect 145665 8449 145699 8483
rect 145932 8449 145966 8483
rect 147505 8449 147539 8483
rect 147772 8449 147806 8483
rect 149529 8449 149563 8483
rect 151001 8449 151035 8483
rect 152841 8449 152875 8483
rect 153853 8449 153887 8483
rect 154681 8449 154715 8483
rect 156153 8449 156187 8483
rect 156337 8449 156371 8483
rect 156797 8449 156831 8483
rect 156981 8449 157015 8483
rect 158085 8449 158119 8483
rect 3893 8381 3927 8415
rect 4353 8381 4387 8415
rect 6929 8381 6963 8415
rect 16865 8381 16899 8415
rect 17233 8381 17267 8415
rect 30665 8381 30699 8415
rect 31033 8381 31067 8415
rect 31769 8381 31803 8415
rect 44005 8381 44039 8415
rect 46673 8381 46707 8415
rect 50813 8381 50847 8415
rect 57529 8381 57563 8415
rect 58081 8381 58115 8415
rect 67833 8381 67867 8415
rect 68385 8381 68419 8415
rect 90373 8381 90407 8415
rect 94145 8381 94179 8415
rect 111533 8381 111567 8415
rect 116409 8381 116443 8415
rect 117973 8381 118007 8415
rect 118341 8381 118375 8415
rect 118801 8381 118835 8415
rect 119169 8381 119203 8415
rect 119905 8381 119939 8415
rect 120457 8381 120491 8415
rect 123033 8381 123067 8415
rect 125149 8381 125183 8415
rect 126805 8381 126839 8415
rect 128829 8381 128863 8415
rect 132969 8381 133003 8415
rect 133429 8381 133463 8415
rect 136925 8381 136959 8415
rect 139409 8381 139443 8415
rect 139961 8381 139995 8415
rect 149345 8381 149379 8415
rect 152013 8381 152047 8415
rect 152289 8381 152323 8415
rect 154037 8381 154071 8415
rect 154865 8381 154899 8415
rect 6561 8313 6595 8347
rect 7481 8313 7515 8347
rect 12357 8313 12391 8347
rect 16037 8313 16071 8347
rect 17693 8313 17727 8347
rect 33977 8313 34011 8347
rect 36369 8313 36403 8347
rect 38209 8313 38243 8347
rect 40049 8313 40083 8347
rect 44465 8313 44499 8347
rect 52009 8313 52043 8347
rect 53941 8313 53975 8347
rect 56517 8313 56551 8347
rect 59461 8313 59495 8347
rect 66913 8313 66947 8347
rect 73537 8313 73571 8347
rect 74917 8313 74951 8347
rect 78137 8313 78171 8347
rect 84025 8313 84059 8347
rect 86785 8313 86819 8347
rect 93317 8313 93351 8347
rect 94513 8313 94547 8347
rect 108129 8313 108163 8347
rect 110981 8313 111015 8347
rect 115857 8313 115891 8347
rect 121837 8313 121871 8347
rect 124413 8313 124447 8347
rect 128093 8313 128127 8347
rect 134809 8313 134843 8347
rect 138029 8313 138063 8347
rect 138581 8313 138615 8347
rect 140697 8313 140731 8347
rect 141157 8313 141191 8347
rect 141801 8313 141835 8347
rect 147045 8313 147079 8347
rect 148885 8313 148919 8347
rect 154497 8313 154531 8347
rect 155969 8313 156003 8347
rect 157165 8313 157199 8347
rect 158269 8313 158303 8347
rect 4721 8245 4755 8279
rect 18889 8245 18923 8279
rect 32873 8245 32907 8279
rect 42625 8245 42659 8279
rect 47133 8245 47167 8279
rect 60473 8245 60507 8279
rect 65533 8245 65567 8279
rect 74365 8245 74399 8279
rect 90833 8245 90867 8279
rect 92765 8245 92799 8279
rect 108773 8245 108807 8279
rect 116869 8245 116903 8279
rect 131037 8245 131071 8279
rect 136373 8245 136407 8279
rect 150173 8245 150207 8279
rect 152933 8245 152967 8279
rect 153669 8245 153703 8279
rect 6377 8041 6411 8075
rect 12909 8041 12943 8075
rect 14381 8041 14415 8075
rect 15301 8041 15335 8075
rect 18613 8041 18647 8075
rect 21557 8041 21591 8075
rect 26065 8041 26099 8075
rect 31033 8041 31067 8075
rect 31585 8041 31619 8075
rect 36185 8041 36219 8075
rect 36737 8041 36771 8075
rect 38393 8041 38427 8075
rect 42809 8041 42843 8075
rect 43269 8041 43303 8075
rect 45385 8041 45419 8075
rect 46673 8041 46707 8075
rect 48605 8041 48639 8075
rect 49249 8041 49283 8075
rect 55873 8041 55907 8075
rect 56885 8041 56919 8075
rect 59553 8041 59587 8075
rect 63325 8041 63359 8075
rect 68937 8041 68971 8075
rect 74825 8041 74859 8075
rect 76757 8041 76791 8075
rect 80621 8041 80655 8075
rect 84485 8041 84519 8075
rect 125333 8041 125367 8075
rect 127633 8041 127667 8075
rect 137385 8041 137419 8075
rect 152105 8041 152139 8075
rect 157257 8041 157291 8075
rect 5733 7973 5767 8007
rect 32505 7973 32539 8007
rect 35541 7973 35575 8007
rect 39129 7973 39163 8007
rect 50997 7973 51031 8007
rect 53021 7973 53055 8007
rect 57437 7973 57471 8007
rect 61209 7973 61243 8007
rect 65901 7973 65935 8007
rect 86969 7973 87003 8007
rect 90465 7973 90499 8007
rect 91569 7973 91603 8007
rect 93501 7973 93535 8007
rect 99757 7973 99791 8007
rect 110521 7973 110555 8007
rect 112637 7973 112671 8007
rect 122481 7973 122515 8007
rect 132141 7973 132175 8007
rect 141433 7973 141467 8007
rect 144469 7973 144503 8007
rect 144929 7973 144963 8007
rect 150357 7973 150391 8007
rect 12357 7905 12391 7939
rect 37749 7905 37783 7939
rect 40049 7905 40083 7939
rect 41429 7905 41463 7939
rect 47225 7905 47259 7939
rect 48053 7905 48087 7939
rect 50445 7905 50479 7939
rect 52377 7905 52411 7939
rect 67005 7905 67039 7939
rect 67557 7905 67591 7939
rect 85865 7905 85899 7939
rect 118617 7905 118651 7939
rect 121653 7905 121687 7939
rect 129013 7905 129047 7939
rect 132785 7905 132819 7939
rect 133061 7905 133095 7939
rect 140145 7905 140179 7939
rect 147137 7905 147171 7939
rect 147505 7905 147539 7939
rect 156797 7905 156831 7939
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 6193 7837 6227 7871
rect 13553 7837 13587 7871
rect 14933 7837 14967 7871
rect 15117 7837 15151 7871
rect 16129 7837 16163 7871
rect 18153 7837 18187 7871
rect 20177 7837 20211 7871
rect 22109 7837 22143 7871
rect 25881 7837 25915 7871
rect 31769 7837 31803 7871
rect 34345 7837 34379 7871
rect 35357 7837 35391 7871
rect 36921 7837 36955 7871
rect 38577 7837 38611 7871
rect 39313 7837 39347 7871
rect 40233 7837 40267 7871
rect 40417 7837 40451 7871
rect 40877 7837 40911 7871
rect 41696 7837 41730 7871
rect 44649 7837 44683 7871
rect 45845 7837 45879 7871
rect 46029 7839 46063 7873
rect 47409 7837 47443 7871
rect 52837 7837 52871 7871
rect 54125 7837 54159 7871
rect 54217 7837 54251 7871
rect 54953 7837 54987 7871
rect 58817 7837 58851 7871
rect 62333 7837 62367 7871
rect 62589 7837 62623 7871
rect 64705 7837 64739 7871
rect 66085 7837 66119 7871
rect 72065 7837 72099 7871
rect 72617 7837 72651 7871
rect 72884 7837 72918 7871
rect 74457 7837 74491 7871
rect 74641 7837 74675 7871
rect 76297 7837 76331 7871
rect 81265 7837 81299 7871
rect 86785 7837 86819 7871
rect 87429 7837 87463 7871
rect 87613 7837 87647 7871
rect 87705 7837 87739 7871
rect 91017 7837 91051 7871
rect 92949 7837 92983 7871
rect 95341 7837 95375 7871
rect 98377 7837 98411 7871
rect 105737 7837 105771 7871
rect 109141 7837 109175 7871
rect 111165 7837 111199 7871
rect 112821 7837 112855 7871
rect 112913 7837 112947 7871
rect 113741 7837 113775 7871
rect 115581 7837 115615 7871
rect 117881 7837 117915 7871
rect 118801 7837 118835 7871
rect 119445 7837 119479 7871
rect 123953 7837 123987 7871
rect 124229 7837 124263 7871
rect 129749 7837 129783 7871
rect 129933 7837 129967 7871
rect 130117 7837 130151 7871
rect 130669 7837 130703 7871
rect 130761 7837 130795 7871
rect 131497 7837 131531 7871
rect 135821 7837 135855 7871
rect 138121 7837 138155 7871
rect 140789 7837 140823 7871
rect 140973 7837 141007 7871
rect 141617 7837 141651 7871
rect 143089 7837 143123 7871
rect 146309 7837 146343 7871
rect 147321 7837 147355 7871
rect 148241 7837 148275 7871
rect 150817 7837 150851 7871
rect 151093 7837 151127 7871
rect 152289 7837 152323 7871
rect 152381 7837 152415 7871
rect 153577 7837 153611 7871
rect 153761 7837 153795 7871
rect 154497 7837 154531 7871
rect 154753 7837 154787 7871
rect 156613 7837 156647 7871
rect 157441 7837 157475 7871
rect 7021 7769 7055 7803
rect 17886 7769 17920 7803
rect 20444 7769 20478 7803
rect 34078 7769 34112 7803
rect 44382 7769 44416 7803
rect 52110 7769 52144 7803
rect 56333 7769 56367 7803
rect 58550 7769 58584 7803
rect 64438 7769 64472 7803
rect 67802 7769 67836 7803
rect 85598 7769 85632 7803
rect 92682 7769 92716 7803
rect 98644 7769 98678 7803
rect 109408 7769 109442 7803
rect 114008 7769 114042 7803
rect 116225 7769 116259 7803
rect 121193 7769 121227 7803
rect 122665 7769 122699 7803
rect 128746 7769 128780 7803
rect 135576 7769 135610 7803
rect 136373 7769 136407 7803
rect 139878 7769 139912 7803
rect 142169 7769 142203 7803
rect 143356 7769 143390 7803
rect 146042 7769 146076 7803
rect 148508 7769 148542 7803
rect 150173 7769 150207 7803
rect 4813 7701 4847 7735
rect 13369 7701 13403 7735
rect 16313 7701 16347 7735
rect 16773 7701 16807 7735
rect 19441 7701 19475 7735
rect 22293 7701 22327 7735
rect 32965 7701 32999 7735
rect 46213 7701 46247 7735
rect 47593 7701 47627 7735
rect 49801 7701 49835 7735
rect 53941 7701 53975 7735
rect 54769 7701 54803 7735
rect 60749 7701 60783 7735
rect 65257 7701 65291 7735
rect 73997 7701 74031 7735
rect 76113 7701 76147 7735
rect 82553 7701 82587 7735
rect 94053 7701 94087 7735
rect 95157 7701 95191 7735
rect 97825 7701 97859 7735
rect 100309 7701 100343 7735
rect 105921 7701 105955 7735
rect 110981 7701 111015 7735
rect 115121 7701 115155 7735
rect 116777 7701 116811 7735
rect 117697 7701 117731 7735
rect 118985 7701 119019 7735
rect 123217 7701 123251 7735
rect 125885 7701 125919 7735
rect 126437 7701 126471 7735
rect 127081 7701 127115 7735
rect 130945 7701 130979 7735
rect 134441 7701 134475 7735
rect 137937 7701 137971 7735
rect 138765 7701 138799 7735
rect 140605 7701 140639 7735
rect 142445 7701 142479 7735
rect 149621 7701 149655 7735
rect 153393 7701 153427 7735
rect 155877 7701 155911 7735
rect 156429 7701 156463 7735
rect 157993 7701 158027 7735
rect 5273 7497 5307 7531
rect 6009 7497 6043 7531
rect 14105 7497 14139 7531
rect 15117 7497 15151 7531
rect 16865 7497 16899 7531
rect 21097 7497 21131 7531
rect 32873 7497 32907 7531
rect 34713 7497 34747 7531
rect 36737 7497 36771 7531
rect 38577 7497 38611 7531
rect 40509 7497 40543 7531
rect 41429 7497 41463 7531
rect 41981 7497 42015 7531
rect 43085 7497 43119 7531
rect 45201 7497 45235 7531
rect 49341 7497 49375 7531
rect 50445 7497 50479 7531
rect 57437 7497 57471 7531
rect 58081 7497 58115 7531
rect 58725 7497 58759 7531
rect 59737 7497 59771 7531
rect 63233 7497 63267 7531
rect 64797 7497 64831 7531
rect 65257 7497 65291 7531
rect 67097 7497 67131 7531
rect 71605 7497 71639 7531
rect 74089 7497 74123 7531
rect 76573 7497 76607 7531
rect 97365 7497 97399 7531
rect 127173 7497 127207 7531
rect 127725 7497 127759 7531
rect 128737 7497 128771 7531
rect 129381 7497 129415 7531
rect 130209 7497 130243 7531
rect 130853 7497 130887 7531
rect 131773 7497 131807 7531
rect 133429 7497 133463 7531
rect 136097 7497 136131 7531
rect 141893 7497 141927 7531
rect 150817 7497 150851 7531
rect 155325 7497 155359 7531
rect 157625 7497 157659 7531
rect 15761 7429 15795 7463
rect 30113 7429 30147 7463
rect 31125 7429 31159 7463
rect 32413 7429 32447 7463
rect 39374 7429 39408 7463
rect 46489 7429 46523 7463
rect 52132 7429 52166 7463
rect 66085 7429 66119 7463
rect 79324 7429 79358 7463
rect 111616 7429 111650 7463
rect 122950 7429 122984 7463
rect 132877 7429 132911 7463
rect 134542 7429 134576 7463
rect 144000 7429 144034 7463
rect 147352 7429 147386 7463
rect 148508 7429 148542 7463
rect 151930 7429 151964 7463
rect 158269 7429 158303 7463
rect 4813 7361 4847 7395
rect 5457 7361 5491 7395
rect 13461 7361 13495 7395
rect 13645 7361 13679 7395
rect 14289 7361 14323 7395
rect 16313 7361 16347 7395
rect 17417 7361 17451 7395
rect 18245 7361 18279 7395
rect 21281 7361 21315 7395
rect 26074 7361 26108 7395
rect 29285 7361 29319 7395
rect 29469 7361 29503 7395
rect 33986 7361 34020 7395
rect 34253 7361 34287 7395
rect 35826 7361 35860 7395
rect 36553 7361 36587 7395
rect 41245 7361 41279 7395
rect 53205 7361 53239 7395
rect 53849 7361 53883 7395
rect 54861 7361 54895 7395
rect 58265 7361 58299 7395
rect 60565 7361 60599 7395
rect 63417 7361 63451 7395
rect 64613 7361 64647 7395
rect 66913 7361 66947 7395
rect 72729 7361 72763 7395
rect 75213 7361 75247 7395
rect 81440 7361 81474 7395
rect 84669 7361 84703 7395
rect 91569 7361 91603 7395
rect 91836 7361 91870 7395
rect 96546 7361 96580 7395
rect 96813 7361 96847 7395
rect 110521 7361 110555 7395
rect 110705 7361 110739 7395
rect 114109 7361 114143 7395
rect 116777 7361 116811 7395
rect 117237 7361 117271 7395
rect 119097 7361 119131 7395
rect 121121 7361 121155 7395
rect 127909 7361 127943 7395
rect 128553 7361 128587 7395
rect 130393 7361 130427 7395
rect 134809 7361 134843 7395
rect 135361 7361 135395 7395
rect 138397 7361 138431 7395
rect 139225 7361 139259 7395
rect 140881 7361 140915 7395
rect 141065 7361 141099 7395
rect 143017 7361 143051 7395
rect 147597 7361 147631 7395
rect 148241 7361 148275 7395
rect 150081 7361 150115 7395
rect 153485 7361 153519 7395
rect 154313 7361 154347 7395
rect 155141 7361 155175 7395
rect 156153 7361 156187 7395
rect 156981 7361 157015 7395
rect 157809 7361 157843 7395
rect 12817 7293 12851 7327
rect 13277 7293 13311 7327
rect 18061 7293 18095 7327
rect 18429 7293 18463 7327
rect 26341 7293 26375 7327
rect 29653 7293 29687 7327
rect 36093 7293 36127 7327
rect 38025 7293 38059 7327
rect 39129 7293 39163 7327
rect 52377 7293 52411 7327
rect 62589 7293 62623 7327
rect 72985 7293 73019 7327
rect 75469 7293 75503 7327
rect 75929 7293 75963 7327
rect 79057 7293 79091 7327
rect 81173 7293 81207 7327
rect 110889 7293 110923 7327
rect 111349 7293 111383 7327
rect 113189 7293 113223 7327
rect 119353 7293 119387 7327
rect 121377 7293 121411 7327
rect 123217 7293 123251 7327
rect 125609 7293 125643 7327
rect 126621 7293 126655 7327
rect 128093 7293 128127 7327
rect 137753 7293 137787 7327
rect 138581 7293 138615 7327
rect 139041 7293 139075 7327
rect 143273 7293 143307 7327
rect 143733 7293 143767 7327
rect 152197 7293 152231 7327
rect 153209 7293 153243 7327
rect 154129 7293 154163 7327
rect 154957 7293 154991 7327
rect 155969 7293 156003 7327
rect 156797 7293 156831 7327
rect 24961 7225 24995 7259
rect 50997 7225 51031 7259
rect 82553 7225 82587 7259
rect 117973 7225 118007 7259
rect 121837 7225 121871 7259
rect 123769 7225 123803 7259
rect 138213 7225 138247 7259
rect 139409 7225 139443 7259
rect 145113 7225 145147 7259
rect 157165 7225 157199 7259
rect 4629 7157 4663 7191
rect 17601 7157 17635 7191
rect 18981 7157 19015 7191
rect 22109 7157 22143 7191
rect 45845 7157 45879 7191
rect 60749 7157 60783 7191
rect 68385 7157 68419 7191
rect 80437 7157 80471 7191
rect 83105 7157 83139 7191
rect 84485 7157 84519 7191
rect 86049 7157 86083 7191
rect 87245 7157 87279 7191
rect 92949 7157 92983 7191
rect 93501 7157 93535 7191
rect 95433 7157 95467 7191
rect 110061 7157 110095 7191
rect 112729 7157 112763 7191
rect 113925 7157 113959 7191
rect 117421 7157 117455 7191
rect 119997 7157 120031 7191
rect 124413 7157 124447 7191
rect 126161 7157 126195 7191
rect 132325 7157 132359 7191
rect 135545 7157 135579 7191
rect 136649 7157 136683 7191
rect 137109 7157 137143 7191
rect 139961 7157 139995 7191
rect 140697 7157 140731 7191
rect 146217 7157 146251 7191
rect 149621 7157 149655 7191
rect 154497 7157 154531 7191
rect 156337 7157 156371 7191
rect 13001 6953 13035 6987
rect 34897 6953 34931 6987
rect 37657 6953 37691 6987
rect 51641 6953 51675 6987
rect 54493 6953 54527 6987
rect 63693 6953 63727 6987
rect 130209 6953 130243 6987
rect 130853 6953 130887 6987
rect 134257 6953 134291 6987
rect 138213 6953 138247 6987
rect 138765 6953 138799 6987
rect 146769 6953 146803 6987
rect 148241 6953 148275 6987
rect 156981 6953 157015 6987
rect 18337 6885 18371 6919
rect 24869 6885 24903 6919
rect 50721 6885 50755 6919
rect 110613 6885 110647 6919
rect 111073 6885 111107 6919
rect 115397 6885 115431 6919
rect 127081 6885 127115 6919
rect 140329 6885 140363 6919
rect 143089 6885 143123 6919
rect 150265 6885 150299 6919
rect 151461 6885 151495 6919
rect 16221 6817 16255 6851
rect 18705 6817 18739 6851
rect 19441 6817 19475 6851
rect 20085 6817 20119 6851
rect 26249 6817 26283 6851
rect 32781 6817 32815 6851
rect 33517 6817 33551 6851
rect 33885 6817 33919 6851
rect 38117 6817 38151 6851
rect 52101 6817 52135 6851
rect 68477 6817 68511 6851
rect 88257 6817 88291 6851
rect 93317 6817 93351 6851
rect 93869 6817 93903 6851
rect 108405 6817 108439 6851
rect 108865 6817 108899 6851
rect 112821 6817 112855 6851
rect 114569 6817 114603 6851
rect 114937 6817 114971 6851
rect 116777 6817 116811 6851
rect 118801 6817 118835 6851
rect 121653 6817 121687 6851
rect 122481 6817 122515 6851
rect 129749 6817 129783 6851
rect 133705 6817 133739 6851
rect 142169 6817 142203 6851
rect 155325 6817 155359 6851
rect 156521 6817 156555 6851
rect 4721 6749 4755 6783
rect 11897 6749 11931 6783
rect 14381 6749 14415 6783
rect 15025 6749 15059 6783
rect 15209 6749 15243 6783
rect 16488 6749 16522 6783
rect 18521 6749 18555 6783
rect 22109 6749 22143 6783
rect 27077 6749 27111 6783
rect 33701 6749 33735 6783
rect 36553 6749 36587 6783
rect 37013 6749 37047 6783
rect 43545 6749 43579 6783
rect 43729 6749 43763 6783
rect 53849 6749 53883 6783
rect 54033 6749 54067 6783
rect 55505 6749 55539 6783
rect 57621 6749 57655 6783
rect 59461 6749 59495 6783
rect 59645 6749 59679 6783
rect 64806 6749 64840 6783
rect 65073 6749 65107 6783
rect 66545 6749 66579 6783
rect 73721 6749 73755 6783
rect 75561 6749 75595 6783
rect 76113 6749 76147 6783
rect 78873 6749 78907 6783
rect 82645 6749 82679 6783
rect 87797 6749 87831 6783
rect 108149 6749 108183 6783
rect 111237 6751 111271 6785
rect 111441 6749 111475 6783
rect 114753 6749 114787 6783
rect 118249 6749 118283 6783
rect 119537 6749 119571 6783
rect 122665 6749 122699 6783
rect 122849 6749 122883 6783
rect 124873 6749 124907 6783
rect 129482 6749 129516 6783
rect 132233 6749 132267 6783
rect 136557 6749 136591 6783
rect 139501 6749 139535 6783
rect 140145 6749 140179 6783
rect 144469 6749 144503 6783
rect 145389 6749 145423 6783
rect 147229 6749 147263 6783
rect 147413 6743 147447 6777
rect 147505 6749 147539 6783
rect 149354 6749 149388 6783
rect 149621 6749 149655 6783
rect 150081 6749 150115 6783
rect 151001 6749 151035 6783
rect 151645 6749 151679 6783
rect 152289 6749 152323 6783
rect 154865 6749 154899 6783
rect 155509 6749 155543 6783
rect 156337 6749 156371 6783
rect 157165 6749 157199 6783
rect 157809 6749 157843 6783
rect 13737 6681 13771 6715
rect 20330 6681 20364 6715
rect 25982 6681 26016 6715
rect 38384 6681 38418 6715
rect 43913 6681 43947 6715
rect 52745 6681 52779 6715
rect 65901 6681 65935 6715
rect 66812 6681 66846 6715
rect 73454 6681 73488 6715
rect 75316 6681 75350 6715
rect 82389 6681 82423 6715
rect 85773 6681 85807 6715
rect 87552 6681 87586 6715
rect 93050 6681 93084 6715
rect 121386 6681 121420 6715
rect 124628 6681 124662 6715
rect 131681 6681 131715 6715
rect 136312 6681 136346 6715
rect 137109 6681 137143 6715
rect 141902 6681 141936 6715
rect 144224 6681 144258 6715
rect 145656 6681 145690 6715
rect 154620 6681 154654 6715
rect 155693 6681 155727 6715
rect 4537 6613 4571 6647
rect 11713 6613 11747 6647
rect 14565 6613 14599 6647
rect 15393 6613 15427 6647
rect 17601 6613 17635 6647
rect 21465 6613 21499 6647
rect 22293 6613 22327 6647
rect 22753 6613 22787 6647
rect 23949 6613 23983 6647
rect 26893 6613 26927 6647
rect 36369 6613 36403 6647
rect 39497 6613 39531 6647
rect 44373 6613 44407 6647
rect 53665 6613 53699 6647
rect 59277 6613 59311 6647
rect 67925 6613 67959 6647
rect 72341 6613 72375 6647
rect 74181 6613 74215 6647
rect 81265 6613 81299 6647
rect 83197 6613 83231 6647
rect 86417 6613 86451 6647
rect 91937 6613 91971 6647
rect 107025 6613 107059 6647
rect 117789 6613 117823 6647
rect 119721 6613 119755 6647
rect 120273 6613 120307 6647
rect 123493 6613 123527 6647
rect 125425 6613 125459 6647
rect 125977 6613 126011 6647
rect 126529 6613 126563 6647
rect 127725 6613 127759 6647
rect 128369 6613 128403 6647
rect 133153 6613 133187 6647
rect 135177 6613 135211 6647
rect 139685 6613 139719 6647
rect 140789 6613 140823 6647
rect 150817 6613 150851 6647
rect 152105 6613 152139 6647
rect 152841 6613 152875 6647
rect 153485 6613 153519 6647
rect 156153 6613 156187 6647
rect 157625 6613 157659 6647
rect 8033 6409 8067 6443
rect 15025 6409 15059 6443
rect 15669 6409 15703 6443
rect 19349 6409 19383 6443
rect 20361 6409 20395 6443
rect 21281 6409 21315 6443
rect 23857 6409 23891 6443
rect 37841 6409 37875 6443
rect 40601 6409 40635 6443
rect 44649 6409 44683 6443
rect 46489 6409 46523 6443
rect 53205 6409 53239 6443
rect 54125 6409 54159 6443
rect 59737 6409 59771 6443
rect 63601 6409 63635 6443
rect 64153 6409 64187 6443
rect 66085 6409 66119 6443
rect 66637 6409 66671 6443
rect 69305 6409 69339 6443
rect 72893 6409 72927 6443
rect 73813 6409 73847 6443
rect 75009 6409 75043 6443
rect 78873 6409 78907 6443
rect 85681 6409 85715 6443
rect 106473 6409 106507 6443
rect 108773 6409 108807 6443
rect 109601 6409 109635 6443
rect 117145 6409 117179 6443
rect 119905 6409 119939 6443
rect 121745 6409 121779 6443
rect 126897 6409 126931 6443
rect 129565 6409 129599 6443
rect 130209 6409 130243 6443
rect 137661 6409 137695 6443
rect 145665 6409 145699 6443
rect 148885 6409 148919 6443
rect 150081 6409 150115 6443
rect 152657 6409 152691 6443
rect 157441 6409 157475 6443
rect 18153 6341 18187 6375
rect 28825 6341 28859 6375
rect 30490 6341 30524 6375
rect 33548 6341 33582 6375
rect 70124 6341 70158 6375
rect 71789 6341 71823 6375
rect 87368 6341 87402 6375
rect 88165 6341 88199 6375
rect 105360 6341 105394 6375
rect 107638 6341 107672 6375
rect 110705 6341 110739 6375
rect 111257 6341 111291 6375
rect 119261 6341 119295 6375
rect 129013 6341 129047 6375
rect 134257 6341 134291 6375
rect 134809 6341 134843 6375
rect 138857 6341 138891 6375
rect 141249 6341 141283 6375
rect 147750 6341 147784 6375
rect 155141 6341 155175 6375
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 9321 6273 9355 6307
rect 14013 6273 14047 6307
rect 15209 6273 15243 6307
rect 15853 6273 15887 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 17785 6273 17819 6307
rect 17969 6273 18003 6307
rect 18613 6273 18647 6307
rect 21097 6273 21131 6307
rect 22201 6273 22235 6307
rect 24970 6273 25004 6307
rect 25697 6273 25731 6307
rect 25973 6273 26007 6307
rect 30757 6273 30791 6307
rect 38393 6273 38427 6307
rect 38660 6273 38694 6307
rect 40233 6273 40267 6307
rect 40417 6273 40451 6307
rect 41061 6273 41095 6307
rect 45762 6273 45796 6307
rect 46673 6273 46707 6307
rect 51641 6273 51675 6307
rect 53389 6273 53423 6307
rect 55238 6273 55272 6307
rect 55505 6273 55539 6307
rect 56517 6273 56551 6307
rect 65277 6273 65311 6307
rect 66821 6273 66855 6307
rect 67281 6273 67315 6307
rect 69857 6273 69891 6307
rect 76133 6273 76167 6307
rect 76941 6273 76975 6307
rect 89812 6273 89846 6307
rect 91477 6273 91511 6307
rect 92121 6273 92155 6307
rect 97356 6273 97390 6307
rect 101597 6273 101631 6307
rect 101873 6273 101907 6307
rect 105093 6273 105127 6307
rect 107393 6273 107427 6307
rect 114017 6273 114051 6307
rect 114201 6273 114235 6307
rect 115866 6273 115900 6307
rect 121029 6273 121063 6307
rect 122869 6273 122903 6307
rect 123125 6273 123159 6307
rect 125517 6273 125551 6307
rect 125784 6273 125818 6307
rect 127357 6273 127391 6307
rect 142813 6273 142847 6307
rect 144581 6273 144615 6307
rect 144837 6273 144871 6307
rect 146789 6273 146823 6307
rect 149345 6273 149379 6307
rect 150265 6273 150299 6307
rect 151001 6273 151035 6307
rect 151829 6273 151863 6307
rect 152841 6273 152875 6307
rect 153669 6273 153703 6307
rect 154865 6273 154899 6307
rect 154957 6273 154991 6307
rect 156153 6273 156187 6307
rect 156981 6273 157015 6307
rect 157625 6273 157659 6307
rect 158269 6273 158303 6307
rect 8677 6205 8711 6239
rect 9505 6205 9539 6239
rect 20913 6205 20947 6239
rect 22017 6205 22051 6239
rect 25237 6205 25271 6239
rect 33793 6205 33827 6239
rect 46029 6205 46063 6239
rect 51457 6205 51491 6239
rect 52285 6205 52319 6239
rect 65533 6205 65567 6239
rect 76389 6205 76423 6239
rect 87613 6205 87647 6239
rect 88993 6205 89027 6239
rect 89545 6205 89579 6239
rect 91937 6205 91971 6239
rect 97089 6205 97123 6239
rect 100953 6205 100987 6239
rect 116133 6205 116167 6239
rect 116685 6205 116719 6239
rect 121285 6205 121319 6239
rect 128001 6205 128035 6239
rect 130945 6205 130979 6239
rect 132601 6205 132635 6239
rect 133613 6205 133647 6239
rect 140513 6205 140547 6239
rect 147045 6205 147079 6239
rect 147505 6205 147539 6239
rect 155969 6205 156003 6239
rect 1777 6137 1811 6171
rect 14565 6137 14599 6171
rect 18797 6137 18831 6171
rect 29377 6137 29411 6171
rect 32413 6137 32447 6171
rect 39773 6137 39807 6171
rect 44189 6137 44223 6171
rect 51825 6137 51859 6171
rect 56701 6137 56735 6171
rect 71237 6137 71271 6171
rect 86233 6137 86267 6171
rect 90925 6137 90959 6171
rect 98469 6137 98503 6171
rect 114753 6137 114787 6171
rect 123677 6137 123711 6171
rect 124413 6137 124447 6171
rect 151645 6137 151679 6171
rect 5549 6069 5583 6103
rect 9137 6069 9171 6103
rect 17233 6069 17267 6103
rect 22385 6069 22419 6103
rect 34253 6069 34287 6103
rect 50905 6069 50939 6103
rect 92305 6069 92339 6103
rect 96629 6069 96663 6103
rect 113281 6069 113315 6103
rect 113833 6069 113867 6103
rect 118249 6069 118283 6103
rect 118801 6069 118835 6103
rect 128553 6069 128587 6103
rect 131497 6069 131531 6103
rect 132049 6069 132083 6103
rect 133061 6069 133095 6103
rect 135821 6069 135855 6103
rect 136373 6069 136407 6103
rect 136833 6069 136867 6103
rect 138213 6069 138247 6103
rect 139409 6069 139443 6103
rect 139961 6069 139995 6103
rect 143457 6069 143491 6103
rect 149529 6069 149563 6103
rect 150817 6069 150851 6103
rect 153761 6069 153795 6103
rect 156337 6069 156371 6103
rect 156797 6069 156831 6103
rect 158085 6069 158119 6103
rect 5365 5865 5399 5899
rect 5825 5865 5859 5899
rect 16129 5865 16163 5899
rect 16957 5865 16991 5899
rect 18337 5865 18371 5899
rect 19625 5865 19659 5899
rect 21833 5865 21867 5899
rect 24777 5865 24811 5899
rect 30021 5865 30055 5899
rect 32321 5865 32355 5899
rect 38025 5865 38059 5899
rect 43269 5865 43303 5899
rect 45477 5865 45511 5899
rect 52193 5865 52227 5899
rect 66637 5865 66671 5899
rect 68937 5865 68971 5899
rect 76205 5865 76239 5899
rect 91845 5865 91879 5899
rect 99389 5865 99423 5899
rect 108865 5865 108899 5899
rect 117421 5865 117455 5899
rect 120825 5865 120859 5899
rect 122481 5865 122515 5899
rect 123125 5865 123159 5899
rect 131865 5865 131899 5899
rect 132877 5865 132911 5899
rect 135729 5865 135763 5899
rect 136281 5865 136315 5899
rect 142353 5865 142387 5899
rect 146309 5865 146343 5899
rect 36001 5797 36035 5831
rect 47317 5797 47351 5831
rect 49249 5797 49283 5831
rect 65257 5797 65291 5831
rect 68477 5797 68511 5831
rect 72709 5797 72743 5831
rect 79057 5797 79091 5831
rect 108405 5797 108439 5831
rect 114385 5797 114419 5831
rect 115397 5797 115431 5831
rect 118341 5797 118375 5831
rect 120365 5797 120399 5831
rect 121745 5797 121779 5831
rect 127081 5797 127115 5831
rect 129013 5797 129047 5831
rect 129749 5797 129783 5831
rect 137293 5797 137327 5831
rect 138489 5797 138523 5831
rect 140329 5797 140363 5831
rect 144469 5797 144503 5831
rect 149621 5797 149655 5831
rect 151645 5797 151679 5831
rect 154037 5797 154071 5831
rect 155325 5797 155359 5831
rect 156981 5797 157015 5831
rect 157625 5797 157659 5831
rect 16497 5729 16531 5763
rect 35449 5729 35483 5763
rect 44649 5729 44683 5763
rect 45845 5729 45879 5763
rect 47869 5729 47903 5763
rect 53573 5729 53607 5763
rect 54677 5729 54711 5763
rect 63877 5729 63911 5763
rect 66177 5729 66211 5763
rect 75469 5729 75503 5763
rect 80437 5729 80471 5763
rect 116777 5729 116811 5763
rect 123677 5729 123711 5763
rect 124597 5729 124631 5763
rect 140973 5729 141007 5763
rect 150449 5729 150483 5763
rect 154865 5729 154899 5763
rect 3985 5661 4019 5695
rect 4252 5661 4286 5695
rect 6009 5661 6043 5695
rect 11805 5661 11839 5695
rect 13185 5661 13219 5695
rect 13737 5661 13771 5695
rect 14289 5661 14323 5695
rect 14556 5661 14590 5695
rect 16313 5661 16347 5695
rect 17141 5661 17175 5695
rect 17325 5661 17359 5695
rect 19809 5661 19843 5695
rect 24593 5661 24627 5695
rect 30205 5661 30239 5695
rect 30389 5661 30423 5695
rect 37114 5661 37148 5695
rect 37381 5661 37415 5695
rect 37841 5661 37875 5695
rect 45661 5661 45695 5695
rect 54217 5661 54251 5695
rect 58633 5661 58667 5695
rect 64133 5661 64167 5695
rect 65993 5661 66027 5695
rect 70050 5661 70084 5695
rect 70317 5661 70351 5695
rect 72893 5661 72927 5695
rect 73077 5661 73111 5695
rect 76757 5661 76791 5695
rect 80170 5661 80204 5695
rect 81265 5661 81299 5695
rect 95341 5661 95375 5695
rect 101321 5661 101355 5695
rect 107025 5661 107059 5695
rect 118525 5661 118559 5695
rect 118985 5661 119019 5695
rect 121009 5661 121043 5695
rect 121193 5661 121227 5695
rect 125793 5661 125827 5695
rect 127633 5661 127667 5695
rect 127900 5661 127934 5695
rect 130393 5661 130427 5695
rect 133981 5661 134015 5695
rect 134533 5661 134567 5695
rect 136741 5661 136775 5695
rect 138029 5661 138063 5695
rect 139869 5661 139903 5695
rect 140513 5661 140547 5695
rect 143089 5661 143123 5695
rect 144929 5661 144963 5695
rect 146769 5661 146803 5695
rect 146953 5661 146987 5695
rect 148241 5661 148275 5695
rect 150081 5661 150115 5695
rect 150265 5661 150299 5695
rect 151093 5661 151127 5695
rect 151829 5661 151863 5695
rect 152473 5661 152507 5695
rect 153669 5661 153703 5695
rect 153853 5661 153887 5695
rect 154589 5661 154623 5695
rect 154681 5661 154715 5695
rect 155509 5661 155543 5695
rect 155601 5661 155635 5695
rect 156153 5661 156187 5695
rect 156337 5661 156371 5695
rect 157165 5661 157199 5695
rect 157809 5661 157843 5695
rect 44382 5593 44416 5627
rect 48125 5593 48159 5627
rect 53328 5593 53362 5627
rect 73537 5593 73571 5627
rect 75224 5593 75258 5627
rect 83013 5593 83047 5627
rect 95074 5593 95108 5627
rect 101054 5593 101088 5627
rect 107292 5593 107326 5627
rect 116532 5593 116566 5627
rect 119252 5593 119286 5627
rect 130209 5593 130243 5627
rect 131313 5593 131347 5627
rect 131957 5593 131991 5627
rect 135085 5593 135119 5627
rect 139624 5593 139658 5627
rect 141218 5593 141252 5627
rect 143356 5593 143390 5627
rect 145196 5593 145230 5627
rect 148486 5593 148520 5627
rect 156521 5593 156555 5627
rect 11621 5525 11655 5559
rect 13001 5525 13035 5559
rect 15669 5525 15703 5559
rect 30849 5525 30883 5559
rect 38577 5525 38611 5559
rect 54033 5525 54067 5559
rect 58449 5525 58483 5559
rect 65809 5525 65843 5559
rect 74089 5525 74123 5559
rect 78045 5525 78079 5559
rect 93409 5525 93443 5559
rect 93961 5525 93995 5559
rect 99941 5525 99975 5559
rect 101965 5525 101999 5559
rect 125057 5525 125091 5559
rect 125609 5525 125643 5559
rect 126437 5525 126471 5559
rect 133429 5525 133463 5559
rect 147137 5525 147171 5559
rect 147689 5525 147723 5559
rect 150909 5525 150943 5559
rect 152289 5525 152323 5559
rect 6653 5321 6687 5355
rect 13645 5321 13679 5355
rect 16313 5321 16347 5355
rect 16865 5321 16899 5355
rect 17601 5321 17635 5355
rect 18153 5321 18187 5355
rect 19901 5321 19935 5355
rect 24133 5321 24167 5355
rect 27261 5321 27295 5355
rect 35357 5321 35391 5355
rect 48513 5321 48547 5355
rect 54309 5321 54343 5355
rect 62405 5321 62439 5355
rect 63325 5321 63359 5355
rect 65717 5321 65751 5355
rect 73537 5321 73571 5355
rect 75929 5321 75963 5355
rect 115673 5321 115707 5355
rect 116317 5321 116351 5355
rect 118525 5321 118559 5355
rect 121285 5321 121319 5355
rect 123125 5321 123159 5355
rect 124505 5321 124539 5355
rect 127725 5321 127759 5355
rect 129105 5321 129139 5355
rect 129657 5321 129691 5355
rect 137845 5321 137879 5355
rect 138397 5321 138431 5355
rect 139317 5321 139351 5355
rect 139961 5321 139995 5355
rect 144653 5321 144687 5355
rect 145665 5321 145699 5355
rect 153025 5321 153059 5355
rect 156797 5321 156831 5355
rect 158085 5321 158119 5355
rect 23020 5253 23054 5287
rect 24593 5253 24627 5287
rect 34897 5253 34931 5287
rect 45385 5253 45419 5287
rect 55658 5253 55692 5287
rect 75009 5253 75043 5287
rect 77217 5253 77251 5287
rect 104900 5253 104934 5287
rect 106565 5253 106599 5287
rect 120172 5253 120206 5287
rect 123861 5253 123895 5287
rect 132049 5253 132083 5287
rect 137569 5253 137603 5287
rect 151930 5253 151964 5287
rect 154957 5253 154991 5287
rect 3801 5185 3835 5219
rect 4068 5185 4102 5219
rect 5917 5185 5951 5219
rect 12265 5185 12299 5219
rect 12532 5185 12566 5219
rect 15025 5185 15059 5219
rect 15209 5185 15243 5219
rect 19717 5185 19751 5219
rect 26157 5185 26191 5219
rect 29662 5185 29696 5219
rect 31502 5185 31536 5219
rect 34253 5185 34287 5219
rect 36481 5185 36515 5219
rect 36737 5185 36771 5219
rect 48697 5185 48731 5219
rect 53196 5185 53230 5219
rect 61025 5185 61059 5219
rect 61281 5185 61315 5219
rect 79057 5185 79091 5219
rect 82553 5185 82587 5219
rect 90741 5185 90775 5219
rect 92417 5185 92451 5219
rect 92673 5185 92707 5219
rect 93133 5185 93167 5219
rect 112361 5185 112395 5219
rect 114937 5185 114971 5219
rect 117441 5185 117475 5219
rect 118709 5185 118743 5219
rect 119905 5185 119939 5219
rect 122001 5185 122035 5219
rect 125333 5185 125367 5219
rect 127173 5185 127207 5219
rect 127909 5185 127943 5219
rect 128093 5185 128127 5219
rect 131405 5185 131439 5219
rect 136833 5185 136867 5219
rect 138581 5185 138615 5219
rect 139777 5185 139811 5219
rect 141718 5185 141752 5219
rect 141985 5185 142019 5219
rect 143569 5185 143603 5219
rect 143825 5185 143859 5219
rect 144817 5185 144851 5219
rect 145021 5185 145055 5219
rect 146789 5185 146823 5219
rect 147045 5185 147079 5219
rect 148618 5185 148652 5219
rect 148885 5185 148919 5219
rect 149713 5185 149747 5219
rect 152841 5185 152875 5219
rect 153669 5185 153703 5219
rect 154681 5185 154715 5219
rect 154793 5185 154827 5219
rect 155969 5185 156003 5219
rect 156153 5185 156187 5219
rect 156981 5185 157015 5219
rect 157625 5185 157659 5219
rect 158269 5185 158303 5219
rect 22753 5117 22787 5151
rect 29929 5117 29963 5151
rect 31769 5117 31803 5151
rect 52929 5117 52963 5151
rect 55413 5117 55447 5151
rect 82369 5117 82403 5151
rect 104633 5117 104667 5151
rect 114109 5117 114143 5151
rect 114753 5117 114787 5151
rect 117697 5117 117731 5151
rect 121745 5117 121779 5151
rect 125057 5117 125091 5151
rect 133613 5117 133647 5151
rect 152197 5117 152231 5151
rect 152657 5117 152691 5151
rect 5733 5049 5767 5083
rect 15393 5049 15427 5083
rect 34069 5049 34103 5083
rect 78873 5049 78907 5083
rect 93317 5049 93351 5083
rect 130393 5049 130427 5083
rect 135729 5049 135763 5083
rect 140605 5049 140639 5083
rect 5181 4981 5215 5015
rect 14565 4981 14599 5015
rect 28549 4981 28583 5015
rect 30389 4981 30423 5015
rect 56793 4981 56827 5015
rect 81909 4981 81943 5015
rect 82737 4981 82771 5015
rect 91293 4981 91327 5015
rect 106013 4981 106047 5015
rect 112177 4981 112211 5015
rect 115121 4981 115155 5015
rect 119261 4981 119295 5015
rect 126621 4981 126655 5015
rect 130853 4981 130887 5015
rect 132509 4981 132543 5015
rect 133061 4981 133095 5015
rect 134165 4981 134199 5015
rect 134809 4981 134843 5015
rect 136373 4981 136407 5015
rect 137017 4981 137051 5015
rect 142445 4981 142479 5015
rect 147505 4981 147539 5015
rect 149897 4981 149931 5015
rect 150817 4981 150851 5015
rect 153485 4981 153519 5015
rect 156337 4981 156371 5015
rect 157441 4981 157475 5015
rect 4997 4777 5031 4811
rect 5733 4777 5767 4811
rect 12357 4777 12391 4811
rect 12817 4777 12851 4811
rect 13369 4777 13403 4811
rect 14841 4777 14875 4811
rect 15945 4777 15979 4811
rect 22753 4777 22787 4811
rect 24685 4777 24719 4811
rect 25237 4777 25271 4811
rect 26157 4777 26191 4811
rect 30757 4777 30791 4811
rect 46121 4777 46155 4811
rect 73353 4777 73387 4811
rect 82001 4777 82035 4811
rect 84485 4777 84519 4811
rect 88349 4777 88383 4811
rect 90189 4777 90223 4811
rect 96077 4777 96111 4811
rect 98101 4777 98135 4811
rect 104541 4777 104575 4811
rect 108313 4777 108347 4811
rect 117789 4777 117823 4811
rect 121929 4777 121963 4811
rect 133153 4777 133187 4811
rect 135085 4777 135119 4811
rect 136005 4777 136039 4811
rect 140237 4777 140271 4811
rect 146125 4777 146159 4811
rect 152841 4777 152875 4811
rect 156613 4777 156647 4811
rect 157993 4777 158027 4811
rect 44189 4709 44223 4743
rect 50445 4709 50479 4743
rect 124321 4709 124355 4743
rect 125885 4709 125919 4743
rect 127909 4709 127943 4743
rect 130577 4709 130611 4743
rect 139041 4709 139075 4743
rect 139777 4709 139811 4743
rect 150081 4709 150115 4743
rect 154405 4709 154439 4743
rect 25789 4641 25823 4675
rect 29929 4641 29963 4675
rect 81541 4641 81575 4675
rect 82369 4641 82403 4675
rect 88809 4641 88843 4675
rect 96721 4641 96755 4675
rect 114937 4641 114971 4675
rect 118801 4641 118835 4675
rect 122941 4641 122975 4675
rect 126989 4641 127023 4675
rect 131681 4641 131715 4675
rect 137937 4641 137971 4675
rect 138581 4641 138615 4675
rect 142445 4641 142479 4675
rect 147505 4641 147539 4675
rect 148241 4641 148275 4675
rect 155509 4641 155543 4675
rect 5181 4573 5215 4607
rect 12173 4573 12207 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 17058 4573 17092 4607
rect 17325 4573 17359 4607
rect 20646 4573 20680 4607
rect 20913 4573 20947 4607
rect 21373 4573 21407 4607
rect 25973 4573 26007 4607
rect 26617 4573 26651 4607
rect 30113 4573 30147 4607
rect 30297 4573 30331 4607
rect 30941 4573 30975 4607
rect 42349 4573 42383 4607
rect 42809 4573 42843 4607
rect 46305 4573 46339 4607
rect 52110 4573 52144 4607
rect 52377 4573 52411 4607
rect 73169 4573 73203 4607
rect 82185 4573 82219 4607
rect 84301 4573 84335 4607
rect 89065 4573 89099 4607
rect 92857 4573 92891 4607
rect 109437 4573 109471 4607
rect 109693 4573 109727 4607
rect 118985 4573 119019 4607
rect 119629 4573 119663 4607
rect 125333 4573 125367 4607
rect 129289 4573 129323 4607
rect 129749 4573 129783 4607
rect 133705 4573 133739 4607
rect 133961 4573 133995 4607
rect 137385 4573 137419 4607
rect 139593 4573 139627 4607
rect 140421 4573 140455 4607
rect 140605 4573 140639 4607
rect 143089 4573 143123 4607
rect 143273 4573 143307 4607
rect 143365 4573 143399 4607
rect 144285 4573 144319 4607
rect 144552 4573 144586 4607
rect 148508 4573 148542 4607
rect 151461 4573 151495 4607
rect 151921 4573 151955 4607
rect 152105 4573 152139 4607
rect 153577 4573 153611 4607
rect 153761 4573 153795 4607
rect 154589 4573 154623 4607
rect 155141 4573 155175 4607
rect 155325 4573 155359 4607
rect 156153 4573 156187 4607
rect 156797 4573 156831 4607
rect 157441 4573 157475 4607
rect 21640 4505 21674 4539
rect 43076 4505 43110 4539
rect 76389 4505 76423 4539
rect 96988 4505 97022 4539
rect 98561 4505 98595 4539
rect 114670 4505 114704 4539
rect 120825 4505 120859 4539
rect 123208 4505 123242 4539
rect 126437 4505 126471 4539
rect 129044 4505 129078 4539
rect 137140 4505 137174 4539
rect 142200 4505 142234 4539
rect 147260 4505 147294 4539
rect 151194 4505 151228 4539
rect 153945 4505 153979 4539
rect 14381 4437 14415 4471
rect 17877 4437 17911 4471
rect 18889 4437 18923 4471
rect 19533 4437 19567 4471
rect 50997 4437 51031 4471
rect 113557 4437 113591 4471
rect 115489 4437 115523 4471
rect 119169 4437 119203 4471
rect 120273 4437 120307 4471
rect 121285 4437 121319 4471
rect 124873 4437 124907 4471
rect 131129 4437 131163 4471
rect 132233 4437 132267 4471
rect 141065 4437 141099 4471
rect 145665 4437 145699 4471
rect 149621 4437 149655 4471
rect 152289 4437 152323 4471
rect 155969 4437 156003 4471
rect 157257 4437 157291 4471
rect 42625 4233 42659 4267
rect 62313 4233 62347 4267
rect 125057 4233 125091 4267
rect 141157 4233 141191 4267
rect 12633 4165 12667 4199
rect 16865 4165 16899 4199
rect 30389 4165 30423 4199
rect 119261 4165 119295 4199
rect 128829 4165 128863 4199
rect 144776 4165 144810 4199
rect 145665 4165 145699 4199
rect 149652 4165 149686 4199
rect 154436 4165 154470 4199
rect 8309 4097 8343 4131
rect 13829 4097 13863 4131
rect 14085 4097 14119 4131
rect 15669 4097 15703 4131
rect 15853 4097 15887 4131
rect 16037 4097 16071 4131
rect 17693 4097 17727 4131
rect 18521 4097 18555 4131
rect 18788 4097 18822 4131
rect 20361 4097 20395 4131
rect 43738 4097 43772 4131
rect 44005 4097 44039 4131
rect 47961 4097 47995 4131
rect 50905 4097 50939 4131
rect 55422 4097 55456 4131
rect 61505 4097 61539 4131
rect 61761 4097 61795 4131
rect 75929 4097 75963 4131
rect 79425 4097 79459 4131
rect 104633 4097 104667 4131
rect 104900 4097 104934 4131
rect 106473 4097 106507 4131
rect 108793 4097 108827 4131
rect 110725 4097 110759 4131
rect 118249 4097 118283 4131
rect 118433 4097 118467 4131
rect 118617 4097 118651 4131
rect 120917 4097 120951 4131
rect 121469 4097 121503 4131
rect 123605 4097 123639 4131
rect 123861 4097 123895 4131
rect 124321 4097 124355 4131
rect 125241 4097 125275 4131
rect 126069 4097 126103 4131
rect 126336 4097 126370 4131
rect 131333 4097 131367 4131
rect 133173 4097 133207 4131
rect 138296 4097 138330 4131
rect 142914 4097 142948 4131
rect 145021 4097 145055 4131
rect 145849 4097 145883 4131
rect 147801 4097 147835 4131
rect 149897 4097 149931 4131
rect 152022 4097 152056 4131
rect 152749 4097 152783 4131
rect 155325 4097 155359 4131
rect 155969 4097 156003 4131
rect 156153 4097 156187 4131
rect 156337 4097 156371 4131
rect 156981 4097 157015 4131
rect 157625 4097 157659 4131
rect 158269 4097 158303 4131
rect 12357 4029 12391 4063
rect 41981 4029 42015 4063
rect 55689 4029 55723 4063
rect 56149 4029 56183 4063
rect 76205 4029 76239 4063
rect 76665 4029 76699 4063
rect 109049 4029 109083 4063
rect 110981 4029 111015 4063
rect 111441 4029 111475 4063
rect 125425 4029 125459 4063
rect 127909 4029 127943 4063
rect 131589 4029 131623 4063
rect 133429 4029 133463 4063
rect 134165 4029 134199 4063
rect 134809 4029 134843 4063
rect 135913 4029 135947 4063
rect 136465 4029 136499 4063
rect 138029 4029 138063 4063
rect 143181 4029 143215 4063
rect 146033 4029 146067 4063
rect 148057 4029 148091 4063
rect 152289 4029 152323 4063
rect 154681 4029 154715 4063
rect 8125 3961 8159 3995
rect 54309 3961 54343 3995
rect 107669 3961 107703 3995
rect 109601 3961 109635 3995
rect 122481 3961 122515 3995
rect 127449 3961 127483 3995
rect 130209 3961 130243 3995
rect 137017 3961 137051 3995
rect 137569 3961 137603 3995
rect 139409 3961 139443 3995
rect 139961 3961 139995 3995
rect 141801 3961 141835 3995
rect 155141 3961 155175 3995
rect 158085 3961 158119 3995
rect 11713 3893 11747 3927
rect 13369 3893 13403 3927
rect 15209 3893 15243 3927
rect 17877 3893 17911 3927
rect 19901 3893 19935 3927
rect 21189 3893 21223 3927
rect 32873 3893 32907 3927
rect 47777 3893 47811 3927
rect 50721 3893 50755 3927
rect 60381 3893 60415 3927
rect 74825 3893 74859 3927
rect 79609 3893 79643 3927
rect 106013 3893 106047 3927
rect 119169 3893 119203 3927
rect 119905 3893 119939 3927
rect 122021 3893 122055 3927
rect 129289 3893 129323 3927
rect 132049 3893 132083 3927
rect 140513 3893 140547 3927
rect 143641 3893 143675 3927
rect 146677 3893 146711 3927
rect 148517 3893 148551 3927
rect 150909 3893 150943 3927
rect 153301 3893 153335 3927
rect 156797 3893 156831 3927
rect 157441 3893 157475 3927
rect 13277 3689 13311 3723
rect 16681 3689 16715 3723
rect 18889 3689 18923 3723
rect 20821 3689 20855 3723
rect 23305 3689 23339 3723
rect 24869 3689 24903 3723
rect 25697 3689 25731 3723
rect 30573 3689 30607 3723
rect 32965 3689 32999 3723
rect 37013 3689 37047 3723
rect 49801 3689 49835 3723
rect 63049 3689 63083 3723
rect 64889 3689 64923 3723
rect 73169 3689 73203 3723
rect 88441 3689 88475 3723
rect 94513 3689 94547 3723
rect 96813 3689 96847 3723
rect 101873 3689 101907 3723
rect 115397 3689 115431 3723
rect 119629 3689 119663 3723
rect 121929 3689 121963 3723
rect 126713 3689 126747 3723
rect 127633 3689 127667 3723
rect 140421 3689 140455 3723
rect 141985 3689 142019 3723
rect 142537 3689 142571 3723
rect 146309 3689 146343 3723
rect 149897 3689 149931 3723
rect 152841 3689 152875 3723
rect 16221 3621 16255 3655
rect 32505 3621 32539 3655
rect 36553 3621 36587 3655
rect 45201 3621 45235 3655
rect 72617 3621 72651 3655
rect 88993 3621 89027 3655
rect 98745 3621 98779 3655
rect 125517 3621 125551 3655
rect 129473 3621 129507 3655
rect 138489 3621 138523 3655
rect 156797 3621 156831 3655
rect 31125 3553 31159 3587
rect 58541 3553 58575 3587
rect 59001 3553 59035 3587
rect 77493 3553 77527 3587
rect 90373 3553 90407 3587
rect 103253 3553 103287 3587
rect 110153 3553 110187 3587
rect 110705 3553 110739 3587
rect 116777 3553 116811 3587
rect 121009 3553 121043 3587
rect 131405 3553 131439 3587
rect 144193 3553 144227 3587
rect 151829 3553 151863 3587
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 16865 3485 16899 3519
rect 16957 3485 16991 3519
rect 17509 3485 17543 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 21925 3485 21959 3519
rect 25329 3485 25363 3519
rect 25513 3485 25547 3519
rect 34345 3485 34379 3519
rect 37197 3485 37231 3519
rect 37381 3485 37415 3519
rect 46581 3485 46615 3519
rect 48421 3485 48455 3519
rect 53757 3485 53791 3519
rect 58285 3485 58319 3519
rect 61301 3485 61335 3519
rect 62405 3485 62439 3519
rect 65073 3485 65107 3519
rect 74282 3485 74316 3519
rect 74549 3485 74583 3519
rect 90117 3485 90151 3519
rect 95637 3485 95671 3519
rect 95893 3485 95927 3519
rect 100125 3485 100159 3519
rect 100677 3485 100711 3519
rect 109693 3485 109727 3519
rect 117789 3485 117823 3519
rect 123585 3485 123619 3519
rect 124137 3485 124171 3519
rect 125977 3485 126011 3519
rect 126897 3485 126931 3519
rect 127081 3485 127115 3519
rect 129013 3485 129047 3519
rect 130853 3485 130887 3519
rect 131865 3485 131899 3519
rect 132785 3485 132819 3519
rect 132969 3485 133003 3519
rect 133153 3485 133187 3519
rect 134165 3485 134199 3519
rect 135361 3485 135395 3519
rect 135913 3485 135947 3519
rect 138029 3485 138063 3519
rect 139869 3485 139903 3519
rect 143549 3485 143583 3519
rect 147689 3485 147723 3519
rect 148517 3485 148551 3519
rect 152473 3485 152507 3519
rect 152657 3485 152691 3519
rect 155141 3485 155175 3519
rect 155785 3485 155819 3519
rect 155877 3485 155911 3519
rect 156981 3485 157015 3519
rect 157625 3485 157659 3519
rect 17754 3417 17788 3451
rect 19686 3417 19720 3451
rect 22170 3417 22204 3451
rect 31381 3417 31415 3451
rect 34078 3417 34112 3451
rect 37841 3417 37875 3451
rect 46314 3417 46348 3451
rect 48688 3417 48722 3451
rect 62037 3417 62071 3451
rect 77226 3417 77260 3451
rect 77953 3417 77987 3451
rect 99880 3417 99914 3451
rect 102986 3417 103020 3451
rect 109448 3417 109482 3451
rect 116532 3417 116566 3451
rect 118056 3417 118090 3451
rect 120742 3417 120776 3451
rect 124404 3417 124438 3451
rect 128768 3417 128802 3451
rect 130608 3417 130642 3451
rect 133613 3417 133647 3451
rect 139624 3417 139658 3451
rect 144438 3417 144472 3451
rect 147444 3417 147478 3451
rect 148762 3417 148796 3451
rect 151562 3417 151596 3451
rect 154896 3417 154930 3451
rect 14289 3349 14323 3383
rect 15577 3349 15611 3383
rect 23857 3349 23891 3383
rect 44557 3349 44591 3383
rect 53573 3349 53607 3383
rect 57161 3349 57195 3383
rect 76113 3349 76147 3383
rect 108313 3349 108347 3383
rect 119169 3349 119203 3383
rect 122481 3349 122515 3383
rect 123033 3349 123067 3383
rect 134717 3349 134751 3383
rect 136465 3349 136499 3383
rect 136925 3349 136959 3383
rect 140973 3349 141007 3383
rect 143733 3349 143767 3383
rect 145573 3349 145607 3383
rect 150449 3349 150483 3383
rect 153761 3349 153795 3383
rect 155601 3349 155635 3383
rect 157441 3349 157475 3383
rect 11069 3145 11103 3179
rect 11713 3145 11747 3179
rect 13737 3145 13771 3179
rect 14197 3145 14231 3179
rect 17049 3145 17083 3179
rect 20085 3145 20119 3179
rect 23949 3145 23983 3179
rect 24501 3145 24535 3179
rect 31677 3145 31711 3179
rect 32689 3145 32723 3179
rect 44465 3145 44499 3179
rect 49157 3145 49191 3179
rect 62589 3145 62623 3179
rect 66269 3145 66303 3179
rect 68477 3145 68511 3179
rect 81265 3145 81299 3179
rect 96261 3145 96295 3179
rect 109601 3145 109635 3179
rect 110153 3145 110187 3179
rect 114845 3145 114879 3179
rect 115673 3145 115707 3179
rect 116961 3145 116995 3179
rect 126805 3145 126839 3179
rect 127909 3145 127943 3179
rect 129105 3145 129139 3179
rect 131129 3145 131163 3179
rect 132877 3145 132911 3179
rect 134165 3145 134199 3179
rect 134717 3145 134751 3179
rect 135453 3145 135487 3179
rect 138673 3145 138707 3179
rect 139869 3145 139903 3179
rect 140605 3145 140639 3179
rect 141433 3145 141467 3179
rect 142537 3145 142571 3179
rect 147045 3145 147079 3179
rect 150817 3145 150851 3179
rect 154589 3145 154623 3179
rect 155417 3145 155451 3179
rect 157257 3145 157291 3179
rect 12848 3077 12882 3111
rect 15393 3077 15427 3111
rect 18490 3077 18524 3111
rect 22814 3077 22848 3111
rect 46130 3077 46164 3111
rect 47225 3077 47259 3111
rect 55597 3077 55631 3111
rect 56416 3077 56450 3111
rect 64346 3077 64380 3111
rect 121101 3077 121135 3111
rect 131589 3077 131623 3111
rect 137560 3077 137594 3111
rect 141893 3077 141927 3111
rect 144776 3077 144810 3111
rect 152013 3077 152047 3111
rect 152197 3077 152231 3111
rect 13553 3009 13587 3043
rect 16865 3009 16899 3043
rect 18245 3009 18279 3043
rect 20729 3009 20763 3043
rect 22569 3009 22603 3043
rect 30553 3009 30587 3043
rect 32505 3009 32539 3043
rect 33701 3009 33735 3043
rect 41806 3009 41840 3043
rect 42073 3009 42107 3043
rect 46397 3009 46431 3043
rect 47777 3009 47811 3043
rect 48044 3009 48078 3043
rect 50730 3009 50764 3043
rect 50997 3009 51031 3043
rect 56149 3009 56183 3043
rect 64613 3009 64647 3043
rect 67382 3009 67416 3043
rect 114017 3009 114051 3043
rect 115489 3009 115523 3043
rect 118249 3009 118283 3043
rect 126161 3009 126195 3043
rect 127449 3009 127483 3043
rect 128645 3009 128679 3043
rect 130945 3009 130979 3043
rect 136566 3009 136600 3043
rect 137293 3009 137327 3043
rect 139409 3009 139443 3043
rect 143181 3009 143215 3043
rect 145932 3009 145966 3043
rect 147505 3009 147539 3043
rect 147772 3009 147806 3043
rect 149529 3009 149563 3043
rect 149713 3009 149747 3043
rect 151001 3009 151035 3043
rect 153669 3009 153703 3043
rect 154405 3009 154439 3043
rect 155233 3009 155267 3043
rect 156613 3009 156647 3043
rect 157073 3009 157107 3043
rect 158269 3009 158303 3043
rect 13093 2941 13127 2975
rect 14841 2941 14875 2975
rect 29745 2941 29779 2975
rect 30297 2941 30331 2975
rect 32321 2941 32355 2975
rect 33149 2941 33183 2975
rect 67649 2941 67683 2975
rect 72801 2941 72835 2975
rect 113833 2941 113867 2975
rect 114201 2941 114235 2975
rect 120089 2941 120123 2975
rect 120641 2941 120675 2975
rect 121653 2941 121687 2975
rect 122205 2941 122239 2975
rect 122849 2941 122883 2975
rect 130761 2941 130795 2975
rect 136833 2941 136867 2975
rect 145021 2941 145055 2975
rect 145665 2941 145699 2975
rect 149345 2941 149379 2975
rect 150265 2941 150299 2975
rect 151185 2941 151219 2975
rect 152749 2941 152783 2975
rect 154221 2941 154255 2975
rect 155049 2941 155083 2975
rect 19625 2873 19659 2907
rect 20913 2873 20947 2907
rect 40141 2873 40175 2907
rect 45017 2873 45051 2907
rect 63233 2873 63267 2907
rect 118065 2873 118099 2907
rect 118801 2873 118835 2907
rect 130209 2873 130243 2907
rect 143641 2873 143675 2907
rect 148885 2873 148919 2907
rect 153485 2873 153519 2907
rect 158085 2873 158119 2907
rect 1685 2805 1719 2839
rect 5825 2805 5859 2839
rect 17601 2805 17635 2839
rect 40693 2805 40727 2839
rect 49617 2805 49651 2839
rect 57529 2805 57563 2839
rect 65717 2805 65751 2839
rect 83013 2805 83047 2839
rect 117605 2805 117639 2839
rect 119353 2805 119387 2839
rect 123401 2805 123435 2839
rect 123861 2805 123895 2839
rect 124413 2805 124447 2839
rect 125149 2805 125183 2839
rect 125977 2805 126011 2839
rect 127265 2805 127299 2839
rect 142997 2805 143031 2839
rect 156429 2805 156463 2839
rect 5273 2601 5307 2635
rect 11161 2601 11195 2635
rect 11897 2601 11931 2635
rect 13277 2601 13311 2635
rect 18245 2601 18279 2635
rect 19809 2601 19843 2635
rect 26433 2601 26467 2635
rect 45385 2601 45419 2635
rect 49525 2601 49559 2635
rect 60105 2601 60139 2635
rect 60749 2601 60783 2635
rect 65809 2601 65843 2635
rect 74181 2601 74215 2635
rect 81449 2601 81483 2635
rect 107577 2601 107611 2635
rect 109601 2601 109635 2635
rect 113189 2601 113223 2635
rect 113649 2601 113683 2635
rect 114753 2601 114787 2635
rect 122849 2601 122883 2635
rect 123401 2601 123435 2635
rect 125977 2601 126011 2635
rect 127081 2601 127115 2635
rect 130209 2601 130243 2635
rect 132141 2601 132175 2635
rect 134625 2601 134659 2635
rect 137293 2601 137327 2635
rect 139501 2601 139535 2635
rect 142537 2601 142571 2635
rect 143089 2601 143123 2635
rect 147045 2601 147079 2635
rect 151645 2601 151679 2635
rect 152197 2601 152231 2635
rect 152749 2601 152783 2635
rect 154497 2601 154531 2635
rect 18889 2533 18923 2567
rect 25973 2533 26007 2567
rect 64889 2533 64923 2567
rect 126437 2533 126471 2567
rect 143733 2533 143767 2567
rect 153393 2533 153427 2567
rect 6561 2465 6595 2499
rect 12265 2465 12299 2499
rect 21189 2465 21223 2499
rect 24593 2465 24627 2499
rect 33793 2465 33827 2499
rect 46213 2465 46247 2499
rect 58725 2465 58759 2499
rect 63509 2465 63543 2499
rect 108957 2465 108991 2499
rect 114017 2465 114051 2499
rect 119353 2465 119387 2499
rect 129565 2465 129599 2499
rect 131589 2465 131623 2499
rect 133245 2465 133279 2499
rect 135361 2465 135395 2499
rect 141985 2465 142019 2499
rect 145113 2465 145147 2499
rect 145665 2465 145699 2499
rect 148241 2465 148275 2499
rect 151185 2465 151219 2499
rect 154129 2465 154163 2499
rect 155325 2465 155359 2499
rect 157257 2465 157291 2499
rect 1685 2397 1719 2431
rect 5457 2397 5491 2431
rect 5641 2397 5675 2431
rect 12081 2397 12115 2431
rect 18705 2397 18739 2431
rect 20933 2397 20967 2431
rect 24849 2397 24883 2431
rect 45569 2397 45603 2431
rect 45661 2397 45695 2431
rect 58981 2397 59015 2431
rect 63765 2397 63799 2431
rect 73721 2397 73755 2431
rect 75561 2397 75595 2431
rect 82829 2397 82863 2431
rect 108701 2397 108735 2431
rect 113833 2397 113867 2431
rect 118545 2397 118579 2431
rect 118801 2397 118835 2431
rect 121929 2397 121963 2431
rect 130393 2397 130427 2431
rect 130577 2397 130611 2431
rect 135628 2397 135662 2431
rect 138673 2397 138707 2431
rect 138765 2397 138799 2431
rect 138949 2397 138983 2431
rect 144857 2397 144891 2431
rect 147689 2397 147723 2431
rect 150081 2397 150115 2431
rect 151001 2397 151035 2431
rect 154313 2397 154347 2431
rect 155141 2397 155175 2431
rect 156153 2397 156187 2431
rect 156797 2397 156831 2431
rect 2237 2329 2271 2363
rect 33526 2329 33560 2363
rect 44649 2329 44683 2363
rect 75316 2329 75350 2363
rect 82584 2329 82618 2363
rect 119997 2329 120031 2363
rect 128001 2329 128035 2363
rect 129013 2329 129047 2363
rect 131129 2329 131163 2363
rect 133512 2329 133546 2363
rect 138029 2329 138063 2363
rect 141740 2329 141774 2363
rect 145932 2329 145966 2363
rect 148508 2329 148542 2363
rect 150817 2329 150851 2363
rect 154957 2329 154991 2363
rect 31769 2261 31803 2295
rect 32413 2261 32447 2295
rect 117421 2261 117455 2295
rect 120825 2261 120859 2295
rect 121377 2261 121411 2295
rect 123861 2261 123895 2295
rect 124413 2261 124447 2295
rect 125333 2261 125367 2295
rect 128553 2261 128587 2295
rect 136741 2261 136775 2295
rect 140605 2261 140639 2295
rect 147505 2261 147539 2295
rect 149621 2261 149655 2295
rect 155969 2261 156003 2295
rect 156613 2261 156647 2295
rect 157809 2261 157843 2295
<< metal1 >>
rect 146478 15036 146484 15088
rect 146536 15076 146542 15088
rect 154390 15076 154396 15088
rect 146536 15048 154396 15076
rect 146536 15036 146542 15048
rect 154390 15036 154396 15048
rect 154448 15036 154454 15088
rect 145926 14968 145932 15020
rect 145984 15008 145990 15020
rect 154298 15008 154304 15020
rect 145984 14980 154304 15008
rect 145984 14968 145990 14980
rect 154298 14968 154304 14980
rect 154356 14968 154362 15020
rect 96430 14900 96436 14952
rect 96488 14940 96494 14952
rect 149330 14940 149336 14952
rect 96488 14912 149336 14940
rect 96488 14900 96494 14912
rect 149330 14900 149336 14912
rect 149388 14900 149394 14952
rect 118050 14832 118056 14884
rect 118108 14872 118114 14884
rect 150710 14872 150716 14884
rect 118108 14844 150716 14872
rect 118108 14832 118114 14844
rect 150710 14832 150716 14844
rect 150768 14832 150774 14884
rect 109310 14764 109316 14816
rect 109368 14804 109374 14816
rect 141878 14804 141884 14816
rect 109368 14776 141884 14804
rect 109368 14764 109374 14776
rect 141878 14764 141884 14776
rect 141936 14764 141942 14816
rect 146018 14764 146024 14816
rect 146076 14804 146082 14816
rect 152458 14804 152464 14816
rect 146076 14776 152464 14804
rect 146076 14764 146082 14776
rect 152458 14764 152464 14776
rect 152516 14764 152522 14816
rect 114186 14696 114192 14748
rect 114244 14736 114250 14748
rect 157426 14736 157432 14748
rect 114244 14708 157432 14736
rect 114244 14696 114250 14708
rect 157426 14696 157432 14708
rect 157484 14696 157490 14748
rect 119062 14628 119068 14680
rect 119120 14668 119126 14680
rect 152642 14668 152648 14680
rect 119120 14640 152648 14668
rect 119120 14628 119126 14640
rect 152642 14628 152648 14640
rect 152700 14628 152706 14680
rect 130654 14560 130660 14612
rect 130712 14600 130718 14612
rect 156690 14600 156696 14612
rect 130712 14572 156696 14600
rect 130712 14560 130718 14572
rect 156690 14560 156696 14572
rect 156748 14560 156754 14612
rect 134610 14492 134616 14544
rect 134668 14532 134674 14544
rect 149514 14532 149520 14544
rect 134668 14504 149520 14532
rect 134668 14492 134674 14504
rect 149514 14492 149520 14504
rect 149572 14492 149578 14544
rect 149974 14492 149980 14544
rect 150032 14532 150038 14544
rect 154942 14532 154948 14544
rect 150032 14504 154948 14532
rect 150032 14492 150038 14504
rect 154942 14492 154948 14504
rect 155000 14492 155006 14544
rect 129090 14424 129096 14476
rect 129148 14464 129154 14476
rect 150802 14464 150808 14476
rect 129148 14436 150808 14464
rect 129148 14424 129154 14436
rect 150802 14424 150808 14436
rect 150860 14424 150866 14476
rect 107470 14356 107476 14408
rect 107528 14396 107534 14408
rect 132954 14396 132960 14408
rect 107528 14368 132960 14396
rect 107528 14356 107534 14368
rect 132954 14356 132960 14368
rect 133012 14356 133018 14408
rect 134518 14356 134524 14408
rect 134576 14396 134582 14408
rect 154850 14396 154856 14408
rect 134576 14368 154856 14396
rect 134576 14356 134582 14368
rect 154850 14356 154856 14368
rect 154908 14356 154914 14408
rect 125870 14288 125876 14340
rect 125928 14328 125934 14340
rect 153378 14328 153384 14340
rect 125928 14300 153384 14328
rect 125928 14288 125934 14300
rect 153378 14288 153384 14300
rect 153436 14288 153442 14340
rect 124306 14220 124312 14272
rect 124364 14260 124370 14272
rect 152550 14260 152556 14272
rect 124364 14232 152556 14260
rect 124364 14220 124370 14232
rect 152550 14220 152556 14232
rect 152608 14220 152614 14272
rect 129182 14152 129188 14204
rect 129240 14192 129246 14204
rect 156046 14192 156052 14204
rect 129240 14164 156052 14192
rect 129240 14152 129246 14164
rect 156046 14152 156052 14164
rect 156104 14152 156110 14204
rect 129550 14084 129556 14136
rect 129608 14124 129614 14136
rect 153194 14124 153200 14136
rect 129608 14096 153200 14124
rect 129608 14084 129614 14096
rect 153194 14084 153200 14096
rect 153252 14084 153258 14136
rect 51074 14016 51080 14068
rect 51132 14056 51138 14068
rect 53742 14056 53748 14068
rect 51132 14028 53748 14056
rect 51132 14016 51138 14028
rect 53742 14016 53748 14028
rect 53800 14016 53806 14068
rect 138474 14016 138480 14068
rect 138532 14056 138538 14068
rect 155954 14056 155960 14068
rect 138532 14028 155960 14056
rect 138532 14016 138538 14028
rect 155954 14016 155960 14028
rect 156012 14016 156018 14068
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 11238 13988 11244 14000
rect 10100 13960 11244 13988
rect 10100 13948 10106 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 41386 13960 70394 13988
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 15286 13920 15292 13932
rect 12584 13892 15292 13920
rect 12584 13880 12590 13892
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 41386 13852 41414 13960
rect 43898 13880 43904 13932
rect 43956 13920 43962 13932
rect 47118 13920 47124 13932
rect 43956 13892 47124 13920
rect 43956 13880 43962 13892
rect 47118 13880 47124 13892
rect 47176 13880 47182 13932
rect 50706 13880 50712 13932
rect 50764 13920 50770 13932
rect 50764 13892 51488 13920
rect 50764 13880 50770 13892
rect 4120 13824 41414 13852
rect 43088 13824 51396 13852
rect 4120 13812 4126 13824
rect 10410 13744 10416 13796
rect 10468 13784 10474 13796
rect 15194 13784 15200 13796
rect 10468 13756 15200 13784
rect 10468 13744 10474 13756
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 19610 13784 19616 13796
rect 15344 13756 19616 13784
rect 15344 13744 15350 13756
rect 19610 13744 19616 13756
rect 19668 13744 19674 13796
rect 24578 13784 24584 13796
rect 22066 13756 24584 13784
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 12710 13716 12716 13728
rect 7892 13688 12716 13716
rect 7892 13676 7898 13688
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 22066 13716 22094 13756
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 24762 13744 24768 13796
rect 24820 13784 24826 13796
rect 28258 13784 28264 13796
rect 24820 13756 28264 13784
rect 24820 13744 24826 13756
rect 28258 13744 28264 13756
rect 28316 13744 28322 13796
rect 36262 13744 36268 13796
rect 36320 13784 36326 13796
rect 41322 13784 41328 13796
rect 36320 13756 41328 13784
rect 36320 13744 36326 13756
rect 41322 13744 41328 13756
rect 41380 13744 41386 13796
rect 41414 13744 41420 13796
rect 41472 13784 41478 13796
rect 41472 13756 42472 13784
rect 41472 13744 41478 13756
rect 17460 13688 22094 13716
rect 17460 13676 17466 13688
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 27890 13716 27896 13728
rect 22428 13688 27896 13716
rect 22428 13676 22434 13688
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 36170 13676 36176 13728
rect 36228 13716 36234 13728
rect 42334 13716 42340 13728
rect 36228 13688 42340 13716
rect 36228 13676 36234 13688
rect 42334 13676 42340 13688
rect 42392 13676 42398 13728
rect 42444 13716 42472 13756
rect 42518 13744 42524 13796
rect 42576 13784 42582 13796
rect 43088 13784 43116 13824
rect 42576 13756 43116 13784
rect 42576 13744 42582 13756
rect 43162 13744 43168 13796
rect 43220 13784 43226 13796
rect 45094 13784 45100 13796
rect 43220 13756 45100 13784
rect 43220 13744 43226 13756
rect 45094 13744 45100 13756
rect 45152 13744 45158 13796
rect 46658 13784 46664 13796
rect 45204 13756 46664 13784
rect 45204 13716 45232 13756
rect 46658 13744 46664 13756
rect 46716 13744 46722 13796
rect 46934 13744 46940 13796
rect 46992 13784 46998 13796
rect 50614 13784 50620 13796
rect 46992 13756 50620 13784
rect 46992 13744 46998 13756
rect 50614 13744 50620 13756
rect 50672 13744 50678 13796
rect 42444 13688 45232 13716
rect 45554 13676 45560 13728
rect 45612 13716 45618 13728
rect 46106 13716 46112 13728
rect 45612 13688 46112 13716
rect 45612 13676 45618 13688
rect 46106 13676 46112 13688
rect 46164 13676 46170 13728
rect 48130 13676 48136 13728
rect 48188 13716 48194 13728
rect 50706 13716 50712 13728
rect 48188 13688 50712 13716
rect 48188 13676 48194 13688
rect 50706 13676 50712 13688
rect 50764 13676 50770 13728
rect 51368 13716 51396 13824
rect 51460 13784 51488 13892
rect 65518 13880 65524 13932
rect 65576 13920 65582 13932
rect 65576 13892 66024 13920
rect 65576 13880 65582 13892
rect 60550 13784 60556 13796
rect 51460 13756 60556 13784
rect 60550 13744 60556 13756
rect 60608 13744 60614 13796
rect 61378 13744 61384 13796
rect 61436 13784 61442 13796
rect 65886 13784 65892 13796
rect 61436 13756 65892 13784
rect 61436 13744 61442 13756
rect 65886 13744 65892 13756
rect 65944 13744 65950 13796
rect 65996 13784 66024 13892
rect 70366 13852 70394 13960
rect 100754 13948 100760 14000
rect 100812 13988 100818 14000
rect 128906 13988 128912 14000
rect 100812 13960 128912 13988
rect 100812 13948 100818 13960
rect 128906 13948 128912 13960
rect 128964 13948 128970 14000
rect 128998 13948 129004 14000
rect 129056 13988 129062 14000
rect 129056 13960 135254 13988
rect 129056 13948 129062 13960
rect 104250 13880 104256 13932
rect 104308 13920 104314 13932
rect 133046 13920 133052 13932
rect 104308 13892 133052 13920
rect 104308 13880 104314 13892
rect 133046 13880 133052 13892
rect 133104 13880 133110 13932
rect 80606 13852 80612 13864
rect 70366 13824 80612 13852
rect 80606 13812 80612 13824
rect 80664 13812 80670 13864
rect 123018 13852 123024 13864
rect 122024 13824 123024 13852
rect 65996 13756 90864 13784
rect 90836 13728 90864 13756
rect 94038 13744 94044 13796
rect 94096 13784 94102 13796
rect 95786 13784 95792 13796
rect 94096 13756 95792 13784
rect 94096 13744 94102 13756
rect 95786 13744 95792 13756
rect 95844 13744 95850 13796
rect 95878 13744 95884 13796
rect 95936 13784 95942 13796
rect 98730 13784 98736 13796
rect 95936 13756 98736 13784
rect 95936 13744 95942 13756
rect 98730 13744 98736 13756
rect 98788 13744 98794 13796
rect 102318 13744 102324 13796
rect 102376 13784 102382 13796
rect 104342 13784 104348 13796
rect 102376 13756 104348 13784
rect 102376 13744 102382 13756
rect 104342 13744 104348 13756
rect 104400 13784 104406 13796
rect 106642 13784 106648 13796
rect 104400 13756 106648 13784
rect 104400 13744 104406 13756
rect 106642 13744 106648 13756
rect 106700 13744 106706 13796
rect 106826 13744 106832 13796
rect 106884 13784 106890 13796
rect 115658 13784 115664 13796
rect 106884 13756 115664 13784
rect 106884 13744 106890 13756
rect 115658 13744 115664 13756
rect 115716 13744 115722 13796
rect 122024 13784 122052 13824
rect 123018 13812 123024 13824
rect 123076 13812 123082 13864
rect 115860 13756 122052 13784
rect 66622 13716 66628 13728
rect 51368 13688 66628 13716
rect 66622 13676 66628 13688
rect 66680 13676 66686 13728
rect 73982 13676 73988 13728
rect 74040 13716 74046 13728
rect 82078 13716 82084 13728
rect 74040 13688 82084 13716
rect 74040 13676 74046 13688
rect 82078 13676 82084 13688
rect 82136 13676 82142 13728
rect 82170 13676 82176 13728
rect 82228 13716 82234 13728
rect 87874 13716 87880 13728
rect 82228 13688 87880 13716
rect 82228 13676 82234 13688
rect 87874 13676 87880 13688
rect 87932 13676 87938 13728
rect 88058 13676 88064 13728
rect 88116 13716 88122 13728
rect 89714 13716 89720 13728
rect 88116 13688 89720 13716
rect 88116 13676 88122 13688
rect 89714 13676 89720 13688
rect 89772 13676 89778 13728
rect 90818 13676 90824 13728
rect 90876 13716 90882 13728
rect 94866 13716 94872 13728
rect 90876 13688 94872 13716
rect 90876 13676 90882 13688
rect 94866 13676 94872 13688
rect 94924 13676 94930 13728
rect 104158 13676 104164 13728
rect 104216 13716 104222 13728
rect 109586 13716 109592 13728
rect 104216 13688 109592 13716
rect 104216 13676 104222 13688
rect 109586 13676 109592 13688
rect 109644 13676 109650 13728
rect 109678 13676 109684 13728
rect 109736 13716 109742 13728
rect 115860 13716 115888 13756
rect 122098 13744 122104 13796
rect 122156 13784 122162 13796
rect 127342 13784 127348 13796
rect 122156 13756 127348 13784
rect 122156 13744 122162 13756
rect 127342 13744 127348 13756
rect 127400 13744 127406 13796
rect 135226 13784 135254 13960
rect 138750 13948 138756 14000
rect 138808 13988 138814 14000
rect 157610 13988 157616 14000
rect 138808 13960 157616 13988
rect 138808 13948 138814 13960
rect 157610 13948 157616 13960
rect 157668 13948 157674 14000
rect 138014 13880 138020 13932
rect 138072 13920 138078 13932
rect 138072 13892 147674 13920
rect 138072 13880 138078 13892
rect 146938 13852 146944 13864
rect 145300 13824 146944 13852
rect 140590 13784 140596 13796
rect 135226 13756 140596 13784
rect 140590 13744 140596 13756
rect 140648 13744 140654 13796
rect 141142 13744 141148 13796
rect 141200 13784 141206 13796
rect 145300 13784 145328 13824
rect 146938 13812 146944 13824
rect 146996 13812 147002 13864
rect 147646 13852 147674 13892
rect 148410 13880 148416 13932
rect 148468 13920 148474 13932
rect 148468 13892 152412 13920
rect 148468 13880 148474 13892
rect 149974 13852 149980 13864
rect 147646 13824 149980 13852
rect 149974 13812 149980 13824
rect 150032 13812 150038 13864
rect 150066 13812 150072 13864
rect 150124 13852 150130 13864
rect 152274 13852 152280 13864
rect 150124 13824 152280 13852
rect 150124 13812 150130 13824
rect 152274 13812 152280 13824
rect 152332 13812 152338 13864
rect 152384 13852 152412 13892
rect 152458 13880 152464 13932
rect 152516 13920 152522 13932
rect 158070 13920 158076 13932
rect 152516 13892 158076 13920
rect 152516 13880 152522 13892
rect 158070 13880 158076 13892
rect 158128 13880 158134 13932
rect 152384 13824 153700 13852
rect 141200 13756 145328 13784
rect 141200 13744 141206 13756
rect 145374 13744 145380 13796
rect 145432 13784 145438 13796
rect 153562 13784 153568 13796
rect 145432 13756 153568 13784
rect 145432 13744 145438 13756
rect 153562 13744 153568 13756
rect 153620 13744 153626 13796
rect 153672 13784 153700 13824
rect 156138 13784 156144 13796
rect 153672 13756 156144 13784
rect 156138 13744 156144 13756
rect 156196 13744 156202 13796
rect 109736 13688 115888 13716
rect 109736 13676 109742 13688
rect 120166 13676 120172 13728
rect 120224 13716 120230 13728
rect 127526 13716 127532 13728
rect 120224 13688 127532 13716
rect 120224 13676 120230 13688
rect 127526 13676 127532 13688
rect 127584 13676 127590 13728
rect 139578 13676 139584 13728
rect 139636 13716 139642 13728
rect 146202 13716 146208 13728
rect 139636 13688 146208 13716
rect 139636 13676 139642 13688
rect 146202 13676 146208 13688
rect 146260 13676 146266 13728
rect 149238 13676 149244 13728
rect 149296 13716 149302 13728
rect 153286 13716 153292 13728
rect 149296 13688 153292 13716
rect 149296 13676 149302 13688
rect 153286 13676 153292 13688
rect 153344 13676 153350 13728
rect 1104 13626 158884 13648
rect 1104 13574 20672 13626
rect 20724 13574 20736 13626
rect 20788 13574 20800 13626
rect 20852 13574 20864 13626
rect 20916 13574 20928 13626
rect 20980 13574 60117 13626
rect 60169 13574 60181 13626
rect 60233 13574 60245 13626
rect 60297 13574 60309 13626
rect 60361 13574 60373 13626
rect 60425 13574 99562 13626
rect 99614 13574 99626 13626
rect 99678 13574 99690 13626
rect 99742 13574 99754 13626
rect 99806 13574 99818 13626
rect 99870 13574 139007 13626
rect 139059 13574 139071 13626
rect 139123 13574 139135 13626
rect 139187 13574 139199 13626
rect 139251 13574 139263 13626
rect 139315 13574 158884 13626
rect 1104 13552 158884 13574
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 9214 13512 9220 13524
rect 8435 13484 9220 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10229 13515 10287 13521
rect 10229 13481 10241 13515
rect 10275 13512 10287 13515
rect 12342 13512 12348 13524
rect 10275 13484 12348 13512
rect 10275 13481 10287 13484
rect 10229 13475 10287 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 13541 13515 13599 13521
rect 12544 13484 12756 13512
rect 9585 13447 9643 13453
rect 9585 13413 9597 13447
rect 9631 13444 9643 13447
rect 10042 13444 10048 13456
rect 9631 13416 10048 13444
rect 9631 13413 9643 13416
rect 9585 13407 9643 13413
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 12161 13447 12219 13453
rect 12161 13413 12173 13447
rect 12207 13444 12219 13447
rect 12544 13444 12572 13484
rect 12207 13416 12572 13444
rect 12728 13444 12756 13484
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 15654 13512 15660 13524
rect 13587 13484 15660 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 17221 13515 17279 13521
rect 17221 13481 17233 13515
rect 17267 13512 17279 13515
rect 17862 13512 17868 13524
rect 17267 13484 17868 13512
rect 17267 13481 17279 13484
rect 17221 13475 17279 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 17957 13515 18015 13521
rect 17957 13481 17969 13515
rect 18003 13512 18015 13515
rect 18414 13512 18420 13524
rect 18003 13484 18420 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19518 13512 19524 13524
rect 18739 13484 19524 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20625 13515 20683 13521
rect 20625 13481 20637 13515
rect 20671 13512 20683 13515
rect 21726 13512 21732 13524
rect 20671 13484 21732 13512
rect 20671 13481 20683 13484
rect 20625 13475 20683 13481
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 22186 13512 22192 13524
rect 21836 13484 22192 13512
rect 14550 13444 14556 13456
rect 12728 13416 14556 13444
rect 12207 13413 12219 13416
rect 12161 13407 12219 13413
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 19889 13447 19947 13453
rect 19889 13413 19901 13447
rect 19935 13444 19947 13447
rect 21174 13444 21180 13456
rect 19935 13416 21180 13444
rect 19935 13413 19947 13416
rect 19889 13407 19947 13413
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 21269 13447 21327 13453
rect 21269 13413 21281 13447
rect 21315 13444 21327 13447
rect 21634 13444 21640 13456
rect 21315 13416 21640 13444
rect 21315 13413 21327 13416
rect 21269 13407 21327 13413
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 12526 13376 12532 13388
rect 9416 13348 12532 13376
rect 9416 13320 9444 13348
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 21836 13376 21864 13484
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22373 13515 22431 13521
rect 22373 13481 22385 13515
rect 22419 13512 22431 13515
rect 23934 13512 23940 13524
rect 22419 13484 23940 13512
rect 22419 13481 22431 13484
rect 22373 13475 22431 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 27430 13512 27436 13524
rect 24636 13484 27436 13512
rect 24636 13472 24642 13484
rect 27430 13472 27436 13484
rect 27488 13472 27494 13524
rect 27617 13515 27675 13521
rect 27617 13481 27629 13515
rect 27663 13512 27675 13515
rect 28074 13512 28080 13524
rect 27663 13484 28080 13512
rect 27663 13481 27675 13484
rect 27617 13475 27675 13481
rect 28074 13472 28080 13484
rect 28132 13472 28138 13524
rect 28353 13515 28411 13521
rect 28353 13481 28365 13515
rect 28399 13512 28411 13515
rect 28902 13512 28908 13524
rect 28399 13484 28908 13512
rect 28399 13481 28411 13484
rect 28353 13475 28411 13481
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 29089 13515 29147 13521
rect 29089 13481 29101 13515
rect 29135 13512 29147 13515
rect 30558 13512 30564 13524
rect 29135 13484 30564 13512
rect 29135 13481 29147 13484
rect 29089 13475 29147 13481
rect 30558 13472 30564 13484
rect 30616 13472 30622 13524
rect 32766 13512 32772 13524
rect 32727 13484 32772 13512
rect 32766 13472 32772 13484
rect 32824 13472 32830 13524
rect 33413 13515 33471 13521
rect 33413 13481 33425 13515
rect 33459 13512 33471 13515
rect 34422 13512 34428 13524
rect 33459 13484 34428 13512
rect 33459 13481 33471 13484
rect 33413 13475 33471 13481
rect 34422 13472 34428 13484
rect 34480 13472 34486 13524
rect 35526 13512 35532 13524
rect 34808 13484 35532 13512
rect 22002 13404 22008 13456
rect 22060 13444 22066 13456
rect 22278 13444 22284 13456
rect 22060 13416 22284 13444
rect 22060 13404 22066 13416
rect 22278 13404 22284 13416
rect 22336 13404 22342 13456
rect 23109 13447 23167 13453
rect 23109 13413 23121 13447
rect 23155 13444 23167 13447
rect 25222 13444 25228 13456
rect 23155 13416 25228 13444
rect 23155 13413 23167 13416
rect 23109 13407 23167 13413
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 29270 13444 29276 13456
rect 26528 13416 29276 13444
rect 24946 13376 24952 13388
rect 15580 13348 21864 13376
rect 22572 13348 24952 13376
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 9398 13308 9404 13320
rect 9311 13280 9404 13308
rect 8573 13271 8631 13277
rect 8588 13240 8616 13271
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 10226 13308 10232 13320
rect 9508 13280 10232 13308
rect 9508 13240 9536 13280
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10410 13308 10416 13320
rect 10371 13280 10416 13308
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 11146 13308 11152 13320
rect 10704 13280 11152 13308
rect 8588 13212 9536 13240
rect 7285 13175 7343 13181
rect 7285 13141 7297 13175
rect 7331 13172 7343 13175
rect 10704 13172 10732 13280
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13308 12035 13311
rect 12158 13308 12164 13320
rect 12023 13280 12164 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 13725 13311 13783 13317
rect 12768 13280 12813 13308
rect 12768 13268 12774 13280
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 15580 13308 15608 13348
rect 13771 13280 15608 13308
rect 15657 13311 15715 13317
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15746 13308 15752 13320
rect 15703 13280 15752 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 17402 13308 17408 13320
rect 17363 13280 17408 13308
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18598 13308 18604 13320
rect 18187 13280 18604 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 19886 13308 19892 13320
rect 19751 13280 19892 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 13906 13240 13912 13252
rect 12820 13212 13912 13240
rect 7331 13144 10732 13172
rect 7331 13141 7343 13144
rect 7285 13135 7343 13141
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 10965 13175 11023 13181
rect 10965 13172 10977 13175
rect 10836 13144 10977 13172
rect 10836 13132 10842 13144
rect 10965 13141 10977 13144
rect 11011 13172 11023 13175
rect 12820 13172 12848 13212
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 15102 13240 15108 13252
rect 14016 13212 15108 13240
rect 11011 13144 12848 13172
rect 12897 13175 12955 13181
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 12897 13141 12909 13175
rect 12943 13172 12955 13175
rect 14016 13172 14044 13212
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 15390 13243 15448 13249
rect 15390 13240 15402 13243
rect 15344 13212 15402 13240
rect 15344 13200 15350 13212
rect 15390 13209 15402 13212
rect 15436 13209 15448 13243
rect 15390 13203 15448 13209
rect 16301 13243 16359 13249
rect 16301 13209 16313 13243
rect 16347 13240 16359 13243
rect 17678 13240 17684 13252
rect 16347 13212 17684 13240
rect 16347 13209 16359 13212
rect 16301 13203 16359 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 18892 13240 18920 13271
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 20404 13280 20453 13308
rect 20404 13268 20410 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 21450 13308 21456 13320
rect 21411 13280 21456 13308
rect 20441 13271 20499 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 22572 13317 22600 13348
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 23290 13308 23296 13320
rect 23251 13280 23296 13308
rect 22557 13271 22615 13277
rect 23290 13268 23296 13280
rect 23348 13268 23354 13320
rect 23750 13308 23756 13320
rect 23711 13280 23756 13308
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 25038 13308 25044 13320
rect 23860 13280 25044 13308
rect 21358 13240 21364 13252
rect 18892 13212 21364 13240
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 22186 13200 22192 13252
rect 22244 13240 22250 13252
rect 23860 13240 23888 13280
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25188 13280 25237 13308
rect 25188 13268 25194 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25774 13308 25780 13320
rect 25225 13271 25283 13277
rect 25424 13280 25780 13308
rect 25424 13240 25452 13280
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 22244 13212 23888 13240
rect 23952 13212 25452 13240
rect 25492 13243 25550 13249
rect 22244 13200 22250 13212
rect 14274 13172 14280 13184
rect 12943 13144 14044 13172
rect 14235 13144 14280 13172
rect 12943 13141 12955 13144
rect 12897 13135 12955 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 21542 13172 21548 13184
rect 16448 13144 21548 13172
rect 16448 13132 16454 13144
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 23952 13181 23980 13212
rect 25492 13209 25504 13243
rect 25538 13240 25550 13243
rect 26528 13240 26556 13416
rect 29270 13404 29276 13416
rect 29328 13404 29334 13456
rect 34149 13447 34207 13453
rect 34149 13413 34161 13447
rect 34195 13444 34207 13447
rect 34808 13444 34836 13484
rect 35526 13472 35532 13484
rect 35584 13472 35590 13524
rect 37829 13515 37887 13521
rect 37829 13481 37841 13515
rect 37875 13512 37887 13515
rect 39390 13512 39396 13524
rect 37875 13484 39396 13512
rect 37875 13481 37887 13484
rect 37829 13475 37887 13481
rect 39390 13472 39396 13484
rect 39448 13472 39454 13524
rect 39850 13472 39856 13524
rect 39908 13512 39914 13524
rect 42978 13512 42984 13524
rect 39908 13484 42984 13512
rect 39908 13472 39914 13484
rect 42978 13472 42984 13484
rect 43036 13472 43042 13524
rect 44637 13515 44695 13521
rect 43272 13484 44220 13512
rect 34195 13416 34836 13444
rect 34885 13447 34943 13453
rect 34195 13413 34207 13416
rect 34149 13407 34207 13413
rect 34885 13413 34897 13447
rect 34931 13413 34943 13447
rect 43070 13444 43076 13456
rect 34885 13407 34943 13413
rect 38028 13416 43076 13444
rect 26786 13336 26792 13388
rect 26844 13376 26850 13388
rect 26844 13348 27660 13376
rect 26844 13336 26850 13348
rect 27433 13311 27491 13317
rect 27433 13277 27445 13311
rect 27479 13308 27491 13311
rect 27522 13308 27528 13320
rect 27479 13280 27528 13308
rect 27479 13277 27491 13280
rect 27433 13271 27491 13277
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 27632 13308 27660 13348
rect 27706 13336 27712 13388
rect 27764 13376 27770 13388
rect 30098 13376 30104 13388
rect 27764 13348 30104 13376
rect 27764 13336 27770 13348
rect 30098 13336 30104 13348
rect 30156 13336 30162 13388
rect 34900 13376 34928 13407
rect 33612 13348 34928 13376
rect 28169 13311 28227 13317
rect 28169 13308 28181 13311
rect 27632 13280 28181 13308
rect 28169 13277 28181 13280
rect 28215 13277 28227 13311
rect 28169 13271 28227 13277
rect 28258 13268 28264 13320
rect 28316 13308 28322 13320
rect 28905 13311 28963 13317
rect 28905 13308 28917 13311
rect 28316 13280 28917 13308
rect 28316 13268 28322 13280
rect 28905 13277 28917 13280
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 28994 13268 29000 13320
rect 29052 13308 29058 13320
rect 30193 13311 30251 13317
rect 30193 13308 30205 13311
rect 29052 13280 30205 13308
rect 29052 13268 29058 13280
rect 30193 13277 30205 13280
rect 30239 13277 30251 13311
rect 32582 13308 32588 13320
rect 30193 13271 30251 13277
rect 30392 13280 31754 13308
rect 32543 13280 32588 13308
rect 30392 13240 30420 13280
rect 30466 13249 30472 13252
rect 25538 13212 26556 13240
rect 26620 13212 30420 13240
rect 25538 13209 25550 13212
rect 25492 13203 25550 13209
rect 23937 13175 23995 13181
rect 23937 13141 23949 13175
rect 23983 13141 23995 13175
rect 24762 13172 24768 13184
rect 24723 13144 24768 13172
rect 23937 13135 23995 13141
rect 24762 13132 24768 13144
rect 24820 13132 24826 13184
rect 24946 13132 24952 13184
rect 25004 13172 25010 13184
rect 26510 13172 26516 13184
rect 25004 13144 26516 13172
rect 25004 13132 25010 13144
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 26620 13181 26648 13212
rect 30460 13203 30472 13249
rect 30524 13240 30530 13252
rect 30524 13212 30560 13240
rect 30466 13200 30472 13203
rect 30524 13200 30530 13212
rect 26605 13175 26663 13181
rect 26605 13141 26617 13175
rect 26651 13141 26663 13175
rect 26605 13135 26663 13141
rect 26694 13132 26700 13184
rect 26752 13172 26758 13184
rect 31573 13175 31631 13181
rect 31573 13172 31585 13175
rect 26752 13144 31585 13172
rect 26752 13132 26758 13144
rect 31573 13141 31585 13144
rect 31619 13141 31631 13175
rect 31726 13172 31754 13280
rect 32582 13268 32588 13280
rect 32640 13268 32646 13320
rect 33612 13317 33640 13348
rect 33597 13311 33655 13317
rect 33597 13277 33609 13311
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 34333 13311 34391 13317
rect 34333 13277 34345 13311
rect 34379 13308 34391 13311
rect 34790 13308 34796 13320
rect 34379 13280 34796 13308
rect 34379 13277 34391 13280
rect 34333 13271 34391 13277
rect 34790 13268 34796 13280
rect 34848 13268 34854 13320
rect 36009 13311 36067 13317
rect 36009 13277 36021 13311
rect 36055 13308 36067 13311
rect 36170 13308 36176 13320
rect 36055 13280 36176 13308
rect 36055 13277 36067 13280
rect 36009 13271 36067 13277
rect 36170 13268 36176 13280
rect 36228 13268 36234 13320
rect 38028 13317 38056 13416
rect 43070 13404 43076 13416
rect 43128 13404 43134 13456
rect 41046 13376 41052 13388
rect 38856 13348 41052 13376
rect 36265 13311 36323 13317
rect 36265 13277 36277 13311
rect 36311 13277 36323 13311
rect 36265 13271 36323 13277
rect 38013 13311 38071 13317
rect 38013 13277 38025 13311
rect 38059 13277 38071 13311
rect 38746 13308 38752 13320
rect 38707 13280 38752 13308
rect 38013 13271 38071 13277
rect 34054 13200 34060 13252
rect 34112 13240 34118 13252
rect 34422 13240 34428 13252
rect 34112 13212 34428 13240
rect 34112 13200 34118 13212
rect 34422 13200 34428 13212
rect 34480 13240 34486 13252
rect 36280 13240 36308 13271
rect 38746 13268 38752 13280
rect 38804 13268 38810 13320
rect 34480 13212 36308 13240
rect 34480 13200 34486 13212
rect 35434 13172 35440 13184
rect 31726 13144 35440 13172
rect 31573 13135 31631 13141
rect 35434 13132 35440 13144
rect 35492 13132 35498 13184
rect 36538 13132 36544 13184
rect 36596 13172 36602 13184
rect 36817 13175 36875 13181
rect 36817 13172 36829 13175
rect 36596 13144 36829 13172
rect 36596 13132 36602 13144
rect 36817 13141 36829 13144
rect 36863 13172 36875 13175
rect 37826 13172 37832 13184
rect 36863 13144 37832 13172
rect 36863 13141 36875 13144
rect 36817 13135 36875 13141
rect 37826 13132 37832 13144
rect 37884 13132 37890 13184
rect 38565 13175 38623 13181
rect 38565 13141 38577 13175
rect 38611 13172 38623 13175
rect 38856 13172 38884 13348
rect 41046 13336 41052 13348
rect 41104 13336 41110 13388
rect 43272 13376 43300 13484
rect 44192 13444 44220 13484
rect 44637 13481 44649 13515
rect 44683 13512 44695 13515
rect 50890 13512 50896 13524
rect 44683 13484 50896 13512
rect 44683 13481 44695 13484
rect 44637 13475 44695 13481
rect 50890 13472 50896 13484
rect 50948 13472 50954 13524
rect 55677 13515 55735 13521
rect 51046 13484 54616 13512
rect 45554 13444 45560 13456
rect 44192 13416 45560 13444
rect 45554 13404 45560 13416
rect 45612 13404 45618 13456
rect 46658 13404 46664 13456
rect 46716 13444 46722 13456
rect 48409 13447 48467 13453
rect 48409 13444 48421 13447
rect 46716 13416 48421 13444
rect 46716 13404 46722 13416
rect 48409 13413 48421 13416
rect 48455 13413 48467 13447
rect 48409 13407 48467 13413
rect 49786 13404 49792 13456
rect 49844 13444 49850 13456
rect 51046 13444 51074 13484
rect 49844 13416 51074 13444
rect 49844 13404 49850 13416
rect 41248 13348 43300 13376
rect 39482 13308 39488 13320
rect 39443 13280 39488 13308
rect 39482 13268 39488 13280
rect 39540 13268 39546 13320
rect 40221 13311 40279 13317
rect 40221 13277 40233 13311
rect 40267 13308 40279 13311
rect 40310 13308 40316 13320
rect 40267 13280 40316 13308
rect 40267 13277 40279 13280
rect 40221 13271 40279 13277
rect 40310 13268 40316 13280
rect 40368 13268 40374 13320
rect 40405 13311 40463 13317
rect 40405 13277 40417 13311
rect 40451 13308 40463 13311
rect 41138 13308 41144 13320
rect 40451 13280 41144 13308
rect 40451 13277 40463 13280
rect 40405 13271 40463 13277
rect 41138 13268 41144 13280
rect 41196 13268 41202 13320
rect 41248 13317 41276 13348
rect 52914 13336 52920 13388
rect 52972 13376 52978 13388
rect 54588 13376 54616 13484
rect 55677 13481 55689 13515
rect 55723 13512 55735 13515
rect 60093 13515 60151 13521
rect 55723 13484 60044 13512
rect 55723 13481 55735 13484
rect 55677 13475 55735 13481
rect 54941 13447 54999 13453
rect 54941 13413 54953 13447
rect 54987 13444 54999 13447
rect 55858 13444 55864 13456
rect 54987 13416 55864 13444
rect 54987 13413 54999 13416
rect 54941 13407 54999 13413
rect 55858 13404 55864 13416
rect 55916 13404 55922 13456
rect 60016 13444 60044 13484
rect 60093 13481 60105 13515
rect 60139 13512 60151 13515
rect 65981 13515 66039 13521
rect 60139 13484 65840 13512
rect 60139 13481 60151 13484
rect 60093 13475 60151 13481
rect 60642 13444 60648 13456
rect 60016 13416 60648 13444
rect 60642 13404 60648 13416
rect 60700 13404 60706 13456
rect 62209 13447 62267 13453
rect 62209 13413 62221 13447
rect 62255 13444 62267 13447
rect 62255 13416 65748 13444
rect 62255 13413 62267 13416
rect 62209 13407 62267 13413
rect 52972 13348 53696 13376
rect 54588 13348 56272 13376
rect 52972 13336 52978 13348
rect 41233 13311 41291 13317
rect 41233 13277 41245 13311
rect 41279 13277 41291 13311
rect 41233 13271 41291 13277
rect 41322 13268 41328 13320
rect 41380 13308 41386 13320
rect 41506 13308 41512 13320
rect 41380 13280 41512 13308
rect 41380 13268 41386 13280
rect 41506 13268 41512 13280
rect 41564 13308 41570 13320
rect 41693 13311 41751 13317
rect 41693 13308 41705 13311
rect 41564 13280 41705 13308
rect 41564 13268 41570 13280
rect 41693 13277 41705 13280
rect 41739 13277 41751 13311
rect 41874 13308 41880 13320
rect 41835 13280 41880 13308
rect 41693 13271 41751 13277
rect 41874 13268 41880 13280
rect 41932 13268 41938 13320
rect 42061 13311 42119 13317
rect 42061 13277 42073 13311
rect 42107 13308 42119 13311
rect 42613 13311 42671 13317
rect 42613 13308 42625 13311
rect 42107 13280 42625 13308
rect 42107 13277 42119 13280
rect 42061 13271 42119 13277
rect 42613 13277 42625 13280
rect 42659 13277 42671 13311
rect 42613 13271 42671 13277
rect 42702 13268 42708 13320
rect 42760 13308 42766 13320
rect 43257 13311 43315 13317
rect 43257 13308 43269 13311
rect 42760 13280 43269 13308
rect 42760 13268 42766 13280
rect 43257 13277 43269 13280
rect 43303 13308 43315 13311
rect 45922 13308 45928 13320
rect 43303 13280 45928 13308
rect 43303 13277 43315 13280
rect 43257 13271 43315 13277
rect 45922 13268 45928 13280
rect 45980 13268 45986 13320
rect 46569 13311 46627 13317
rect 46569 13308 46581 13311
rect 46400 13280 46581 13308
rect 42426 13240 42432 13252
rect 39316 13212 42432 13240
rect 39316 13181 39344 13212
rect 42426 13200 42432 13212
rect 42484 13200 42490 13252
rect 43162 13240 43168 13252
rect 42628 13212 43168 13240
rect 38611 13144 38884 13172
rect 39301 13175 39359 13181
rect 38611 13141 38623 13144
rect 38565 13135 38623 13141
rect 39301 13141 39313 13175
rect 39347 13141 39359 13175
rect 39301 13135 39359 13141
rect 40037 13175 40095 13181
rect 40037 13141 40049 13175
rect 40083 13172 40095 13175
rect 40126 13172 40132 13184
rect 40083 13144 40132 13172
rect 40083 13141 40095 13144
rect 40037 13135 40095 13141
rect 40126 13132 40132 13144
rect 40184 13132 40190 13184
rect 41049 13175 41107 13181
rect 41049 13141 41061 13175
rect 41095 13172 41107 13175
rect 42628 13172 42656 13212
rect 43162 13200 43168 13212
rect 43220 13200 43226 13252
rect 43524 13243 43582 13249
rect 43524 13209 43536 13243
rect 43570 13240 43582 13243
rect 43714 13240 43720 13252
rect 43570 13212 43720 13240
rect 43570 13209 43582 13212
rect 43524 13203 43582 13209
rect 43714 13200 43720 13212
rect 43772 13200 43778 13252
rect 43806 13200 43812 13252
rect 43864 13240 43870 13252
rect 46302 13243 46360 13249
rect 46302 13240 46314 13243
rect 43864 13212 46314 13240
rect 43864 13200 43870 13212
rect 46302 13209 46314 13212
rect 46348 13209 46360 13243
rect 46302 13203 46360 13209
rect 42794 13172 42800 13184
rect 41095 13144 42656 13172
rect 42755 13144 42800 13172
rect 41095 13141 41107 13144
rect 41049 13135 41107 13141
rect 42794 13132 42800 13144
rect 42852 13132 42858 13184
rect 43622 13132 43628 13184
rect 43680 13172 43686 13184
rect 45189 13175 45247 13181
rect 45189 13172 45201 13175
rect 43680 13144 45201 13172
rect 43680 13132 43686 13144
rect 45189 13141 45201 13144
rect 45235 13141 45247 13175
rect 45189 13135 45247 13141
rect 45554 13132 45560 13184
rect 45612 13172 45618 13184
rect 46400 13172 46428 13280
rect 46569 13277 46581 13280
rect 46615 13308 46627 13311
rect 47210 13308 47216 13320
rect 46615 13280 47216 13308
rect 46615 13277 46627 13280
rect 46569 13271 46627 13277
rect 47210 13268 47216 13280
rect 47268 13268 47274 13320
rect 47949 13311 48007 13317
rect 47949 13277 47961 13311
rect 47995 13308 48007 13311
rect 49694 13308 49700 13320
rect 47995 13280 49700 13308
rect 47995 13277 48007 13280
rect 47949 13271 48007 13277
rect 49694 13268 49700 13280
rect 49752 13268 49758 13320
rect 49789 13311 49847 13317
rect 49789 13277 49801 13311
rect 49835 13308 49847 13311
rect 49878 13308 49884 13320
rect 49835 13280 49884 13308
rect 49835 13277 49847 13280
rect 49789 13271 49847 13277
rect 49878 13268 49884 13280
rect 49936 13268 49942 13320
rect 52365 13311 52423 13317
rect 52365 13308 52377 13311
rect 51046 13280 52377 13308
rect 48314 13200 48320 13252
rect 48372 13240 48378 13252
rect 49522 13243 49580 13249
rect 49522 13240 49534 13243
rect 48372 13212 49534 13240
rect 48372 13200 48378 13212
rect 49522 13209 49534 13212
rect 49568 13209 49580 13243
rect 49712 13240 49740 13268
rect 51046 13240 51074 13280
rect 52365 13277 52377 13280
rect 52411 13277 52423 13311
rect 53558 13308 53564 13320
rect 53519 13280 53564 13308
rect 52365 13271 52423 13277
rect 53558 13268 53564 13280
rect 53616 13268 53622 13320
rect 53668 13304 53696 13348
rect 55398 13308 55404 13320
rect 53760 13304 53880 13308
rect 53668 13280 53880 13304
rect 53668 13276 53788 13280
rect 53852 13249 53880 13280
rect 54404 13280 55404 13308
rect 49712 13212 51074 13240
rect 52120 13243 52178 13249
rect 49522 13203 49580 13209
rect 52120 13209 52132 13243
rect 52166 13240 52178 13243
rect 53828 13243 53886 13249
rect 52166 13212 52399 13240
rect 52166 13209 52178 13212
rect 52120 13203 52178 13209
rect 45612 13144 46428 13172
rect 47213 13175 47271 13181
rect 45612 13132 45618 13144
rect 47213 13141 47225 13175
rect 47259 13172 47271 13175
rect 49786 13172 49792 13184
rect 47259 13144 49792 13172
rect 47259 13141 47271 13144
rect 47213 13135 47271 13141
rect 49786 13132 49792 13144
rect 49844 13132 49850 13184
rect 50525 13175 50583 13181
rect 50525 13141 50537 13175
rect 50571 13172 50583 13175
rect 50706 13172 50712 13184
rect 50571 13144 50712 13172
rect 50571 13141 50583 13144
rect 50525 13135 50583 13141
rect 50706 13132 50712 13144
rect 50764 13132 50770 13184
rect 50798 13132 50804 13184
rect 50856 13172 50862 13184
rect 50985 13175 51043 13181
rect 50985 13172 50997 13175
rect 50856 13144 50997 13172
rect 50856 13132 50862 13144
rect 50985 13141 50997 13144
rect 51031 13141 51043 13175
rect 52371 13172 52399 13212
rect 53828 13209 53840 13243
rect 53874 13240 53886 13243
rect 54404 13240 54432 13280
rect 55398 13268 55404 13280
rect 55456 13268 55462 13320
rect 55493 13311 55551 13317
rect 55493 13277 55505 13311
rect 55539 13277 55551 13311
rect 55493 13271 55551 13277
rect 53874 13212 54432 13240
rect 55508 13240 55536 13271
rect 55582 13268 55588 13320
rect 55640 13308 55646 13320
rect 56137 13311 56195 13317
rect 56137 13308 56149 13311
rect 55640 13280 56149 13308
rect 55640 13268 55646 13280
rect 56137 13277 56149 13280
rect 56183 13277 56195 13311
rect 56244 13308 56272 13348
rect 57164 13348 58848 13376
rect 56393 13311 56451 13317
rect 56393 13308 56405 13311
rect 56244 13280 56405 13308
rect 56137 13271 56195 13277
rect 56393 13277 56405 13280
rect 56439 13277 56451 13311
rect 56393 13271 56451 13277
rect 56686 13268 56692 13320
rect 56744 13308 56750 13320
rect 57164 13308 57192 13348
rect 56744 13280 57192 13308
rect 56744 13268 56750 13280
rect 58618 13268 58624 13320
rect 58676 13308 58682 13320
rect 58713 13311 58771 13317
rect 58713 13308 58725 13311
rect 58676 13280 58725 13308
rect 58676 13268 58682 13280
rect 58713 13277 58725 13280
rect 58759 13277 58771 13311
rect 58820 13308 58848 13348
rect 61856 13348 65656 13376
rect 58820 13280 60504 13308
rect 58713 13271 58771 13277
rect 56042 13240 56048 13252
rect 55508 13212 56048 13240
rect 53874 13209 53886 13212
rect 53828 13203 53886 13209
rect 56042 13200 56048 13212
rect 56100 13200 56106 13252
rect 58958 13243 59016 13249
rect 58958 13240 58970 13243
rect 56612 13212 58970 13240
rect 53006 13172 53012 13184
rect 52371 13144 53012 13172
rect 50985 13135 51043 13141
rect 53006 13132 53012 13144
rect 53064 13132 53070 13184
rect 53101 13175 53159 13181
rect 53101 13141 53113 13175
rect 53147 13172 53159 13175
rect 56612 13172 56640 13212
rect 58958 13209 58970 13212
rect 59004 13240 59016 13243
rect 60366 13240 60372 13252
rect 59004 13212 60372 13240
rect 59004 13209 59016 13212
rect 58958 13203 59016 13209
rect 60366 13200 60372 13212
rect 60424 13200 60430 13252
rect 60476 13240 60504 13280
rect 60642 13268 60648 13320
rect 60700 13308 60706 13320
rect 60734 13308 60740 13320
rect 60700 13280 60740 13308
rect 60700 13268 60706 13280
rect 60734 13268 60740 13280
rect 60792 13268 60798 13320
rect 60826 13268 60832 13320
rect 60884 13308 60890 13320
rect 61856 13308 61884 13348
rect 65628 13320 65656 13348
rect 63402 13308 63408 13320
rect 60884 13280 60929 13308
rect 61028 13280 61884 13308
rect 63363 13280 63408 13308
rect 60884 13268 60890 13280
rect 61028 13240 61056 13280
rect 63402 13268 63408 13280
rect 63460 13268 63466 13320
rect 63497 13311 63555 13317
rect 63497 13277 63509 13311
rect 63543 13277 63555 13311
rect 63497 13271 63555 13277
rect 61102 13249 61108 13252
rect 60476 13212 61056 13240
rect 61096 13203 61108 13249
rect 61160 13240 61166 13252
rect 63512 13240 63540 13271
rect 63586 13268 63592 13320
rect 63644 13308 63650 13320
rect 65518 13308 65524 13320
rect 63644 13280 65524 13308
rect 63644 13268 63650 13280
rect 65518 13268 65524 13280
rect 65576 13268 65582 13320
rect 65610 13268 65616 13320
rect 65668 13268 65674 13320
rect 61160 13212 61196 13240
rect 62132 13212 63540 13240
rect 64325 13243 64383 13249
rect 61102 13200 61108 13203
rect 61160 13200 61166 13212
rect 57514 13172 57520 13184
rect 53147 13144 56640 13172
rect 57475 13144 57520 13172
rect 53147 13141 53159 13144
rect 53101 13135 53159 13141
rect 57514 13132 57520 13144
rect 57572 13132 57578 13184
rect 58253 13175 58311 13181
rect 58253 13141 58265 13175
rect 58299 13172 58311 13175
rect 58802 13172 58808 13184
rect 58299 13144 58808 13172
rect 58299 13141 58311 13144
rect 58253 13135 58311 13141
rect 58802 13132 58808 13144
rect 58860 13132 58866 13184
rect 60642 13132 60648 13184
rect 60700 13172 60706 13184
rect 62132 13172 62160 13212
rect 64325 13209 64337 13243
rect 64371 13240 64383 13243
rect 65150 13240 65156 13252
rect 64371 13212 65156 13240
rect 64371 13209 64383 13212
rect 64325 13203 64383 13209
rect 65150 13200 65156 13212
rect 65208 13200 65214 13252
rect 65720 13240 65748 13416
rect 65812 13317 65840 13484
rect 65981 13481 65993 13515
rect 66027 13512 66039 13515
rect 66438 13512 66444 13524
rect 66027 13484 66444 13512
rect 66027 13481 66039 13484
rect 65981 13475 66039 13481
rect 66438 13472 66444 13484
rect 66496 13472 66502 13524
rect 66622 13512 66628 13524
rect 66583 13484 66628 13512
rect 66622 13472 66628 13484
rect 66680 13472 66686 13524
rect 67637 13515 67695 13521
rect 67637 13481 67649 13515
rect 67683 13512 67695 13515
rect 68094 13512 68100 13524
rect 67683 13484 68100 13512
rect 67683 13481 67695 13484
rect 67637 13475 67695 13481
rect 68094 13472 68100 13484
rect 68152 13472 68158 13524
rect 68833 13515 68891 13521
rect 68833 13481 68845 13515
rect 68879 13512 68891 13515
rect 69198 13512 69204 13524
rect 68879 13484 69204 13512
rect 68879 13481 68891 13484
rect 68833 13475 68891 13481
rect 69198 13472 69204 13484
rect 69256 13472 69262 13524
rect 69477 13515 69535 13521
rect 69477 13481 69489 13515
rect 69523 13512 69535 13515
rect 69934 13512 69940 13524
rect 69523 13484 69940 13512
rect 69523 13481 69535 13484
rect 69477 13475 69535 13481
rect 69934 13472 69940 13484
rect 69992 13472 69998 13524
rect 70213 13515 70271 13521
rect 70213 13481 70225 13515
rect 70259 13512 70271 13515
rect 70854 13512 70860 13524
rect 70259 13484 70860 13512
rect 70259 13481 70271 13484
rect 70213 13475 70271 13481
rect 70854 13472 70860 13484
rect 70912 13472 70918 13524
rect 71314 13512 71320 13524
rect 71275 13484 71320 13512
rect 71314 13472 71320 13484
rect 71372 13472 71378 13524
rect 72050 13512 72056 13524
rect 72011 13484 72056 13512
rect 72050 13472 72056 13484
rect 72108 13472 72114 13524
rect 72786 13512 72792 13524
rect 72747 13484 72792 13512
rect 72786 13472 72792 13484
rect 72844 13472 72850 13524
rect 73890 13512 73896 13524
rect 73851 13484 73896 13512
rect 73890 13472 73896 13484
rect 73948 13472 73954 13524
rect 74626 13512 74632 13524
rect 74587 13484 74632 13512
rect 74626 13472 74632 13484
rect 74684 13472 74690 13524
rect 75454 13512 75460 13524
rect 75415 13484 75460 13512
rect 75454 13472 75460 13484
rect 75512 13472 75518 13524
rect 76193 13515 76251 13521
rect 76193 13481 76205 13515
rect 76239 13512 76251 13515
rect 76926 13512 76932 13524
rect 76239 13484 76932 13512
rect 76239 13481 76251 13484
rect 76193 13475 76251 13481
rect 76926 13472 76932 13484
rect 76984 13472 76990 13524
rect 78030 13512 78036 13524
rect 77991 13484 78036 13512
rect 78030 13472 78036 13484
rect 78088 13472 78094 13524
rect 78953 13515 79011 13521
rect 78953 13481 78965 13515
rect 78999 13512 79011 13515
rect 79134 13512 79140 13524
rect 78999 13484 79140 13512
rect 78999 13481 79011 13484
rect 78953 13475 79011 13481
rect 79134 13472 79140 13484
rect 79192 13472 79198 13524
rect 79778 13512 79784 13524
rect 79739 13484 79784 13512
rect 79778 13472 79784 13484
rect 79836 13472 79842 13524
rect 80238 13472 80244 13524
rect 80296 13512 80302 13524
rect 80425 13515 80483 13521
rect 80425 13512 80437 13515
rect 80296 13484 80437 13512
rect 80296 13472 80302 13484
rect 80425 13481 80437 13484
rect 80471 13481 80483 13515
rect 80425 13475 80483 13481
rect 80790 13472 80796 13524
rect 80848 13512 80854 13524
rect 81437 13515 81495 13521
rect 81437 13512 81449 13515
rect 80848 13484 81449 13512
rect 80848 13472 80854 13484
rect 81437 13481 81449 13484
rect 81483 13481 81495 13515
rect 81437 13475 81495 13481
rect 81894 13472 81900 13524
rect 81952 13512 81958 13524
rect 82817 13515 82875 13521
rect 82817 13512 82829 13515
rect 81952 13484 82829 13512
rect 81952 13472 81958 13484
rect 82817 13481 82829 13484
rect 82863 13481 82875 13515
rect 82817 13475 82875 13481
rect 82998 13472 83004 13524
rect 83056 13512 83062 13524
rect 83921 13515 83979 13521
rect 83921 13512 83933 13515
rect 83056 13484 83933 13512
rect 83056 13472 83062 13484
rect 83921 13481 83933 13484
rect 83967 13481 83979 13515
rect 83921 13475 83979 13481
rect 84102 13472 84108 13524
rect 84160 13512 84166 13524
rect 84562 13512 84568 13524
rect 84160 13484 84568 13512
rect 84160 13472 84166 13484
rect 84562 13472 84568 13484
rect 84620 13472 84626 13524
rect 84654 13472 84660 13524
rect 84712 13512 84718 13524
rect 85393 13515 85451 13521
rect 85393 13512 85405 13515
rect 84712 13484 85405 13512
rect 84712 13472 84718 13484
rect 85393 13481 85405 13484
rect 85439 13481 85451 13515
rect 88702 13512 88708 13524
rect 85393 13475 85451 13481
rect 87432 13484 88708 13512
rect 65886 13404 65892 13456
rect 65944 13444 65950 13456
rect 65944 13416 81296 13444
rect 65944 13404 65950 13416
rect 73982 13376 73988 13388
rect 66272 13348 73988 13376
rect 65797 13311 65855 13317
rect 65797 13277 65809 13311
rect 65843 13277 65855 13311
rect 65797 13271 65855 13277
rect 66272 13240 66300 13348
rect 73982 13336 73988 13348
rect 74040 13336 74046 13388
rect 79962 13376 79968 13388
rect 74092 13348 79968 13376
rect 67821 13311 67879 13317
rect 67821 13277 67833 13311
rect 67867 13277 67879 13311
rect 67821 13271 67879 13277
rect 68649 13311 68707 13317
rect 68649 13277 68661 13311
rect 68695 13308 68707 13311
rect 68830 13308 68836 13320
rect 68695 13280 68836 13308
rect 68695 13277 68707 13280
rect 68649 13271 68707 13277
rect 66898 13240 66904 13252
rect 65720 13212 66300 13240
rect 66859 13212 66904 13240
rect 66898 13200 66904 13212
rect 66956 13200 66962 13252
rect 67836 13240 67864 13271
rect 68830 13268 68836 13280
rect 68888 13268 68894 13320
rect 69658 13308 69664 13320
rect 69619 13280 69664 13308
rect 69658 13268 69664 13280
rect 69716 13268 69722 13320
rect 70397 13311 70455 13317
rect 70397 13277 70409 13311
rect 70443 13308 70455 13311
rect 71130 13308 71136 13320
rect 70443 13280 71136 13308
rect 70443 13277 70455 13280
rect 70397 13271 70455 13277
rect 71130 13268 71136 13280
rect 71188 13268 71194 13320
rect 71501 13311 71559 13317
rect 71501 13277 71513 13311
rect 71547 13308 71559 13311
rect 71682 13308 71688 13320
rect 71547 13280 71688 13308
rect 71547 13277 71559 13280
rect 71501 13271 71559 13277
rect 71682 13268 71688 13280
rect 71740 13268 71746 13320
rect 72237 13311 72295 13317
rect 72237 13277 72249 13311
rect 72283 13277 72295 13311
rect 72237 13271 72295 13277
rect 72973 13311 73031 13317
rect 72973 13277 72985 13311
rect 73019 13308 73031 13311
rect 73890 13308 73896 13320
rect 73019 13280 73896 13308
rect 73019 13277 73031 13280
rect 72973 13271 73031 13277
rect 70946 13240 70952 13252
rect 67836 13212 70952 13240
rect 70946 13200 70952 13212
rect 71004 13200 71010 13252
rect 72252 13240 72280 13271
rect 73890 13268 73896 13280
rect 73948 13268 73954 13320
rect 74092 13317 74120 13348
rect 79962 13336 79968 13348
rect 80020 13336 80026 13388
rect 81268 13376 81296 13416
rect 81342 13404 81348 13456
rect 81400 13444 81406 13456
rect 82081 13447 82139 13453
rect 82081 13444 82093 13447
rect 81400 13416 82093 13444
rect 81400 13404 81406 13416
rect 82081 13413 82093 13416
rect 82127 13413 82139 13447
rect 82081 13407 82139 13413
rect 83182 13404 83188 13456
rect 83240 13444 83246 13456
rect 87049 13447 87107 13453
rect 87049 13444 87061 13447
rect 83240 13416 87061 13444
rect 83240 13404 83246 13416
rect 87049 13413 87061 13416
rect 87095 13413 87107 13447
rect 87049 13407 87107 13413
rect 87432 13376 87460 13484
rect 88702 13472 88708 13484
rect 88760 13472 88766 13524
rect 88794 13472 88800 13524
rect 88852 13512 88858 13524
rect 90637 13515 90695 13521
rect 90637 13512 90649 13515
rect 88852 13484 90649 13512
rect 88852 13472 88858 13484
rect 90637 13481 90649 13484
rect 90683 13481 90695 13515
rect 90637 13475 90695 13481
rect 91002 13472 91008 13524
rect 91060 13512 91066 13524
rect 94225 13515 94283 13521
rect 94225 13512 94237 13515
rect 91060 13484 94237 13512
rect 91060 13472 91066 13484
rect 94225 13481 94237 13484
rect 94271 13481 94283 13515
rect 94225 13475 94283 13481
rect 95142 13472 95148 13524
rect 95200 13512 95206 13524
rect 97537 13515 97595 13521
rect 97537 13512 97549 13515
rect 95200 13484 97549 13512
rect 95200 13472 95206 13484
rect 97537 13481 97549 13484
rect 97583 13481 97595 13515
rect 97537 13475 97595 13481
rect 97994 13472 98000 13524
rect 98052 13512 98058 13524
rect 99377 13515 99435 13521
rect 99377 13512 99389 13515
rect 98052 13484 99389 13512
rect 98052 13472 98058 13484
rect 99377 13481 99389 13484
rect 99423 13481 99435 13515
rect 99377 13475 99435 13481
rect 102870 13472 102876 13524
rect 102928 13512 102934 13524
rect 104529 13515 104587 13521
rect 104529 13512 104541 13515
rect 102928 13484 104541 13512
rect 102928 13472 102934 13484
rect 104529 13481 104541 13484
rect 104575 13481 104587 13515
rect 104529 13475 104587 13481
rect 104802 13472 104808 13524
rect 104860 13512 104866 13524
rect 106093 13515 106151 13521
rect 106093 13512 106105 13515
rect 104860 13484 106105 13512
rect 104860 13472 104866 13484
rect 106093 13481 106105 13484
rect 106139 13481 106151 13515
rect 106093 13475 106151 13481
rect 106642 13472 106648 13524
rect 106700 13512 106706 13524
rect 107013 13515 107071 13521
rect 107013 13512 107025 13515
rect 106700 13484 107025 13512
rect 106700 13472 106706 13484
rect 107013 13481 107025 13484
rect 107059 13512 107071 13515
rect 107654 13512 107660 13524
rect 107059 13484 107660 13512
rect 107059 13481 107071 13484
rect 107013 13475 107071 13481
rect 107654 13472 107660 13484
rect 107712 13472 107718 13524
rect 107838 13472 107844 13524
rect 107896 13512 107902 13524
rect 107896 13484 108620 13512
rect 107896 13472 107902 13484
rect 88610 13404 88616 13456
rect 88668 13444 88674 13456
rect 91094 13444 91100 13456
rect 88668 13416 91100 13444
rect 88668 13404 88674 13416
rect 91094 13404 91100 13416
rect 91152 13404 91158 13456
rect 91741 13447 91799 13453
rect 91741 13413 91753 13447
rect 91787 13413 91799 13447
rect 91741 13407 91799 13413
rect 91756 13376 91784 13407
rect 93210 13404 93216 13456
rect 93268 13444 93274 13456
rect 95697 13447 95755 13453
rect 95697 13444 95709 13447
rect 93268 13416 95709 13444
rect 93268 13404 93274 13416
rect 95697 13413 95709 13416
rect 95743 13413 95755 13447
rect 95697 13407 95755 13413
rect 95786 13404 95792 13456
rect 95844 13444 95850 13456
rect 96801 13447 96859 13453
rect 96801 13444 96813 13447
rect 95844 13416 96813 13444
rect 95844 13404 95850 13416
rect 96801 13413 96813 13416
rect 96847 13413 96859 13447
rect 96801 13407 96859 13413
rect 97074 13404 97080 13456
rect 97132 13444 97138 13456
rect 98365 13447 98423 13453
rect 98365 13444 98377 13447
rect 97132 13416 98377 13444
rect 97132 13404 97138 13416
rect 98365 13413 98377 13416
rect 98411 13413 98423 13447
rect 98365 13407 98423 13413
rect 98454 13404 98460 13456
rect 98512 13444 98518 13456
rect 100205 13447 100263 13453
rect 100205 13444 100217 13447
rect 98512 13416 100217 13444
rect 98512 13404 98518 13416
rect 100205 13413 100217 13416
rect 100251 13413 100263 13447
rect 100205 13407 100263 13413
rect 101214 13404 101220 13456
rect 101272 13444 101278 13456
rect 103149 13447 103207 13453
rect 103149 13444 103161 13447
rect 101272 13416 103161 13444
rect 101272 13404 101278 13416
rect 103149 13413 103161 13416
rect 103195 13413 103207 13447
rect 103149 13407 103207 13413
rect 103514 13404 103520 13456
rect 103572 13444 103578 13456
rect 105265 13447 105323 13453
rect 105265 13444 105277 13447
rect 103572 13416 105277 13444
rect 103572 13404 103578 13416
rect 105265 13413 105277 13416
rect 105311 13413 105323 13447
rect 108592 13444 108620 13484
rect 108942 13472 108948 13524
rect 109000 13512 109006 13524
rect 110417 13515 110475 13521
rect 110417 13512 110429 13515
rect 109000 13484 110429 13512
rect 109000 13472 109006 13484
rect 110417 13481 110429 13484
rect 110463 13481 110475 13515
rect 110417 13475 110475 13481
rect 110598 13472 110604 13524
rect 110656 13512 110662 13524
rect 112257 13515 112315 13521
rect 112257 13512 112269 13515
rect 110656 13484 112269 13512
rect 110656 13472 110662 13484
rect 112257 13481 112269 13484
rect 112303 13481 112315 13515
rect 112257 13475 112315 13481
rect 112806 13472 112812 13524
rect 112864 13512 112870 13524
rect 113729 13515 113787 13521
rect 113729 13512 113741 13515
rect 112864 13484 113741 13512
rect 112864 13472 112870 13484
rect 113729 13481 113741 13484
rect 113775 13481 113787 13515
rect 113729 13475 113787 13481
rect 113910 13472 113916 13524
rect 113968 13512 113974 13524
rect 114925 13515 114983 13521
rect 114925 13512 114937 13515
rect 113968 13484 114937 13512
rect 113968 13472 113974 13484
rect 114925 13481 114937 13484
rect 114971 13481 114983 13515
rect 114925 13475 114983 13481
rect 115566 13472 115572 13524
rect 115624 13512 115630 13524
rect 115624 13484 116624 13512
rect 115624 13472 115630 13484
rect 109681 13447 109739 13453
rect 109681 13444 109693 13447
rect 108592 13416 109693 13444
rect 105265 13407 105323 13413
rect 109681 13413 109693 13416
rect 109727 13413 109739 13447
rect 109681 13407 109739 13413
rect 109770 13404 109776 13456
rect 109828 13444 109834 13456
rect 111153 13447 111211 13453
rect 111153 13444 111165 13447
rect 109828 13416 111165 13444
rect 109828 13404 109834 13416
rect 111153 13413 111165 13416
rect 111199 13413 111211 13447
rect 111153 13407 111211 13413
rect 111426 13404 111432 13456
rect 111484 13444 111490 13456
rect 113085 13447 113143 13453
rect 113085 13444 113097 13447
rect 111484 13416 113097 13444
rect 111484 13404 111490 13416
rect 113085 13413 113097 13416
rect 113131 13413 113143 13447
rect 113085 13407 113143 13413
rect 114462 13404 114468 13456
rect 114520 13444 114526 13456
rect 116397 13447 116455 13453
rect 116397 13444 116409 13447
rect 114520 13416 116409 13444
rect 114520 13404 114526 13416
rect 116397 13413 116409 13416
rect 116443 13413 116455 13447
rect 116596 13444 116624 13484
rect 116670 13472 116676 13524
rect 116728 13512 116734 13524
rect 118145 13515 118203 13521
rect 118145 13512 118157 13515
rect 116728 13484 118157 13512
rect 116728 13472 116734 13484
rect 118145 13481 118157 13484
rect 118191 13481 118203 13515
rect 118145 13475 118203 13481
rect 118326 13472 118332 13524
rect 118384 13512 118390 13524
rect 119985 13515 120043 13521
rect 119985 13512 119997 13515
rect 118384 13484 119997 13512
rect 118384 13472 118390 13484
rect 119985 13481 119997 13484
rect 120031 13481 120043 13515
rect 119985 13475 120043 13481
rect 120534 13472 120540 13524
rect 120592 13512 120598 13524
rect 121457 13515 121515 13521
rect 121457 13512 121469 13515
rect 120592 13484 121469 13512
rect 120592 13472 120598 13484
rect 121457 13481 121469 13484
rect 121503 13481 121515 13515
rect 121457 13475 121515 13481
rect 122742 13472 122748 13524
rect 122800 13512 122806 13524
rect 125137 13515 125195 13521
rect 125137 13512 125149 13515
rect 122800 13484 125149 13512
rect 122800 13472 122806 13484
rect 125137 13481 125149 13484
rect 125183 13481 125195 13515
rect 125137 13475 125195 13481
rect 125502 13472 125508 13524
rect 125560 13512 125566 13524
rect 126609 13515 126667 13521
rect 126609 13512 126621 13515
rect 125560 13484 126621 13512
rect 125560 13472 125566 13484
rect 126609 13481 126621 13484
rect 126655 13481 126667 13515
rect 126609 13475 126667 13481
rect 126882 13472 126888 13524
rect 126940 13512 126946 13524
rect 126940 13484 127848 13512
rect 126940 13472 126946 13484
rect 117501 13447 117559 13453
rect 117501 13444 117513 13447
rect 116596 13416 117513 13444
rect 116397 13407 116455 13413
rect 117501 13413 117513 13416
rect 117547 13413 117559 13447
rect 118881 13447 118939 13453
rect 118881 13444 118893 13447
rect 117501 13407 117559 13413
rect 117884 13416 118893 13444
rect 95050 13376 95056 13388
rect 81268 13348 83044 13376
rect 74077 13311 74135 13317
rect 74077 13277 74089 13311
rect 74123 13277 74135 13311
rect 74077 13271 74135 13277
rect 74813 13311 74871 13317
rect 74813 13277 74825 13311
rect 74859 13308 74871 13311
rect 75086 13308 75092 13320
rect 74859 13280 75092 13308
rect 74859 13277 74871 13280
rect 74813 13271 74871 13277
rect 75086 13268 75092 13280
rect 75144 13268 75150 13320
rect 75273 13311 75331 13317
rect 75273 13277 75285 13311
rect 75319 13308 75331 13311
rect 75362 13308 75368 13320
rect 75319 13280 75368 13308
rect 75319 13277 75331 13280
rect 75273 13271 75331 13277
rect 75362 13268 75368 13280
rect 75420 13268 75426 13320
rect 76377 13311 76435 13317
rect 76377 13277 76389 13311
rect 76423 13308 76435 13311
rect 77110 13308 77116 13320
rect 76423 13280 77116 13308
rect 76423 13277 76435 13280
rect 76377 13271 76435 13277
rect 77110 13268 77116 13280
rect 77168 13268 77174 13320
rect 77202 13268 77208 13320
rect 77260 13317 77266 13320
rect 77260 13311 77281 13317
rect 77269 13277 77281 13311
rect 77849 13311 77907 13317
rect 77849 13308 77861 13311
rect 77260 13271 77281 13277
rect 77404 13280 77861 13308
rect 77260 13268 77266 13271
rect 75730 13240 75736 13252
rect 72252 13212 75736 13240
rect 75730 13200 75736 13212
rect 75788 13200 75794 13252
rect 75822 13200 75828 13252
rect 75880 13240 75886 13252
rect 75880 13212 77064 13240
rect 75880 13200 75886 13212
rect 60700 13144 62160 13172
rect 63681 13175 63739 13181
rect 60700 13132 60706 13144
rect 63681 13141 63693 13175
rect 63727 13172 63739 13175
rect 64138 13172 64144 13184
rect 63727 13144 64144 13172
rect 63727 13141 63739 13144
rect 63681 13135 63739 13141
rect 64138 13132 64144 13144
rect 64196 13132 64202 13184
rect 65061 13175 65119 13181
rect 65061 13141 65073 13175
rect 65107 13172 65119 13175
rect 65886 13172 65892 13184
rect 65107 13144 65892 13172
rect 65107 13141 65119 13144
rect 65061 13135 65119 13141
rect 65886 13132 65892 13144
rect 65944 13132 65950 13184
rect 65978 13132 65984 13184
rect 66036 13172 66042 13184
rect 76929 13175 76987 13181
rect 76929 13172 76941 13175
rect 66036 13144 76941 13172
rect 66036 13132 66042 13144
rect 76929 13141 76941 13144
rect 76975 13141 76987 13175
rect 77036 13172 77064 13212
rect 77404 13172 77432 13280
rect 77849 13277 77861 13280
rect 77895 13277 77907 13311
rect 79134 13308 79140 13320
rect 79095 13280 79140 13308
rect 77849 13271 77907 13277
rect 79134 13268 79140 13280
rect 79192 13268 79198 13320
rect 79597 13311 79655 13317
rect 79597 13277 79609 13311
rect 79643 13277 79655 13311
rect 79597 13271 79655 13277
rect 80609 13311 80667 13317
rect 80609 13277 80621 13311
rect 80655 13308 80667 13311
rect 81066 13308 81072 13320
rect 80655 13280 81072 13308
rect 80655 13277 80667 13280
rect 80609 13271 80667 13277
rect 77036 13144 77432 13172
rect 76929 13135 76987 13141
rect 77570 13132 77576 13184
rect 77628 13172 77634 13184
rect 79612 13172 79640 13271
rect 81066 13268 81072 13280
rect 81124 13268 81130 13320
rect 81158 13268 81164 13320
rect 81216 13308 81222 13320
rect 81253 13311 81311 13317
rect 81253 13308 81265 13311
rect 81216 13280 81265 13308
rect 81216 13268 81222 13280
rect 81253 13277 81265 13280
rect 81299 13277 81311 13311
rect 82262 13308 82268 13320
rect 82223 13280 82268 13308
rect 81253 13271 81311 13277
rect 82262 13268 82268 13280
rect 82320 13268 82326 13320
rect 83016 13317 83044 13348
rect 84856 13348 87460 13376
rect 88352 13348 91784 13376
rect 94240 13348 95056 13376
rect 83001 13311 83059 13317
rect 83001 13277 83013 13311
rect 83047 13308 83059 13311
rect 84010 13308 84016 13320
rect 83047 13280 84016 13308
rect 83047 13277 83059 13280
rect 83001 13271 83059 13277
rect 84010 13268 84016 13280
rect 84068 13268 84074 13320
rect 84105 13311 84163 13317
rect 84105 13277 84117 13311
rect 84151 13308 84163 13311
rect 84286 13308 84292 13320
rect 84151 13280 84292 13308
rect 84151 13277 84163 13280
rect 84105 13271 84163 13277
rect 84286 13268 84292 13280
rect 84344 13268 84350 13320
rect 84856 13317 84884 13348
rect 84841 13311 84899 13317
rect 84841 13277 84853 13311
rect 84887 13277 84899 13311
rect 84841 13271 84899 13277
rect 85577 13311 85635 13317
rect 85577 13277 85589 13311
rect 85623 13308 85635 13311
rect 88352 13308 88380 13348
rect 85623 13280 88380 13308
rect 85623 13277 85635 13280
rect 85577 13271 85635 13277
rect 88426 13268 88432 13320
rect 88484 13308 88490 13320
rect 89438 13308 89444 13320
rect 88484 13280 89444 13308
rect 88484 13268 88490 13280
rect 89438 13268 89444 13280
rect 89496 13268 89502 13320
rect 89625 13311 89683 13317
rect 89625 13277 89637 13311
rect 89671 13308 89683 13311
rect 89714 13308 89720 13320
rect 89671 13280 89720 13308
rect 89671 13277 89683 13280
rect 89625 13271 89683 13277
rect 89714 13268 89720 13280
rect 89772 13308 89778 13320
rect 90542 13308 90548 13320
rect 89772 13280 90548 13308
rect 89772 13268 89778 13280
rect 90542 13268 90548 13280
rect 90600 13268 90606 13320
rect 90818 13308 90824 13320
rect 90779 13280 90824 13308
rect 90818 13268 90824 13280
rect 90876 13268 90882 13320
rect 91370 13268 91376 13320
rect 91428 13308 91434 13320
rect 93121 13311 93179 13317
rect 93121 13308 93133 13311
rect 91428 13280 93133 13308
rect 91428 13268 91434 13280
rect 93121 13277 93133 13280
rect 93167 13277 93179 13311
rect 93121 13271 93179 13277
rect 88058 13240 88064 13252
rect 86604 13212 88064 13240
rect 77628 13144 79640 13172
rect 77628 13132 77634 13144
rect 84562 13132 84568 13184
rect 84620 13172 84626 13184
rect 84657 13175 84715 13181
rect 84657 13172 84669 13175
rect 84620 13144 84669 13172
rect 84620 13132 84626 13144
rect 84657 13141 84669 13144
rect 84703 13141 84715 13175
rect 84657 13135 84715 13141
rect 85482 13132 85488 13184
rect 85540 13172 85546 13184
rect 86405 13175 86463 13181
rect 86405 13172 86417 13175
rect 85540 13144 86417 13172
rect 85540 13132 85546 13144
rect 86405 13141 86417 13144
rect 86451 13172 86463 13175
rect 86604 13172 86632 13212
rect 88058 13200 88064 13212
rect 88116 13200 88122 13252
rect 88184 13243 88242 13249
rect 88184 13209 88196 13243
rect 88230 13240 88242 13243
rect 88610 13240 88616 13252
rect 88230 13212 88616 13240
rect 88230 13209 88242 13212
rect 88184 13203 88242 13209
rect 88610 13200 88616 13212
rect 88668 13200 88674 13252
rect 89254 13200 89260 13252
rect 89312 13240 89318 13252
rect 89993 13243 90051 13249
rect 89993 13240 90005 13243
rect 89312 13212 90005 13240
rect 89312 13200 89318 13212
rect 89993 13209 90005 13212
rect 90039 13240 90051 13243
rect 92474 13240 92480 13252
rect 90039 13212 92480 13240
rect 90039 13209 90051 13212
rect 89993 13203 90051 13209
rect 92474 13200 92480 13212
rect 92532 13200 92538 13252
rect 92876 13243 92934 13249
rect 92876 13209 92888 13243
rect 92922 13240 92934 13243
rect 94240 13240 94268 13348
rect 95050 13336 95056 13348
rect 95108 13336 95114 13388
rect 104158 13376 104164 13388
rect 95712 13348 104164 13376
rect 94406 13308 94412 13320
rect 94367 13280 94412 13308
rect 94406 13268 94412 13280
rect 94464 13308 94470 13320
rect 95145 13311 95203 13317
rect 94464 13280 95096 13308
rect 94464 13268 94470 13280
rect 92922 13212 94268 13240
rect 95068 13240 95096 13280
rect 95145 13277 95157 13311
rect 95191 13308 95203 13311
rect 95418 13308 95424 13320
rect 95191 13280 95424 13308
rect 95191 13277 95203 13280
rect 95145 13271 95203 13277
rect 95418 13268 95424 13280
rect 95476 13268 95482 13320
rect 95602 13268 95608 13320
rect 95660 13308 95666 13320
rect 95712 13308 95740 13348
rect 104158 13336 104164 13348
rect 104216 13336 104222 13388
rect 104268 13348 105952 13376
rect 95878 13308 95884 13320
rect 95660 13280 95740 13308
rect 95839 13280 95884 13308
rect 95660 13268 95666 13280
rect 95878 13268 95884 13280
rect 95936 13268 95942 13320
rect 96982 13308 96988 13320
rect 96943 13280 96988 13308
rect 96982 13268 96988 13280
rect 97040 13268 97046 13320
rect 97718 13308 97724 13320
rect 97679 13280 97724 13308
rect 97718 13268 97724 13280
rect 97776 13268 97782 13320
rect 98181 13311 98239 13317
rect 98181 13277 98193 13311
rect 98227 13277 98239 13311
rect 98181 13271 98239 13277
rect 96614 13240 96620 13252
rect 95068 13212 96620 13240
rect 92922 13209 92934 13212
rect 92876 13203 92934 13209
rect 96614 13200 96620 13212
rect 96672 13200 96678 13252
rect 96890 13200 96896 13252
rect 96948 13240 96954 13252
rect 98196 13240 98224 13271
rect 99466 13268 99472 13320
rect 99524 13308 99530 13320
rect 99561 13311 99619 13317
rect 99561 13308 99573 13311
rect 99524 13280 99573 13308
rect 99524 13268 99530 13280
rect 99561 13277 99573 13280
rect 99607 13277 99619 13311
rect 100018 13308 100024 13320
rect 99979 13280 100024 13308
rect 99561 13271 99619 13277
rect 100018 13268 100024 13280
rect 100076 13268 100082 13320
rect 101033 13311 101091 13317
rect 100128 13280 100984 13308
rect 100128 13240 100156 13280
rect 96948 13212 98224 13240
rect 98288 13212 100156 13240
rect 100956 13240 100984 13280
rect 101033 13277 101045 13311
rect 101079 13308 101091 13311
rect 101858 13308 101864 13320
rect 101079 13280 101864 13308
rect 101079 13277 101091 13280
rect 101033 13271 101091 13277
rect 101858 13268 101864 13280
rect 101916 13268 101922 13320
rect 102318 13308 102324 13320
rect 102279 13280 102324 13308
rect 102318 13268 102324 13280
rect 102376 13268 102382 13320
rect 102413 13311 102471 13317
rect 102413 13277 102425 13311
rect 102459 13308 102471 13311
rect 102502 13308 102508 13320
rect 102459 13280 102508 13308
rect 102459 13277 102471 13280
rect 102413 13271 102471 13277
rect 102502 13268 102508 13280
rect 102560 13308 102566 13320
rect 103054 13308 103060 13320
rect 102560 13280 103060 13308
rect 102560 13268 102566 13280
rect 103054 13268 103060 13280
rect 103112 13268 103118 13320
rect 103333 13311 103391 13317
rect 103333 13277 103345 13311
rect 103379 13308 103391 13311
rect 104066 13308 104072 13320
rect 103379 13280 104072 13308
rect 103379 13277 103391 13280
rect 103333 13271 103391 13277
rect 104066 13268 104072 13280
rect 104124 13268 104130 13320
rect 104268 13240 104296 13348
rect 105924 13317 105952 13348
rect 110506 13336 110512 13388
rect 110564 13376 110570 13388
rect 110564 13348 112944 13376
rect 110564 13336 110570 13348
rect 104713 13311 104771 13317
rect 104713 13277 104725 13311
rect 104759 13277 104771 13311
rect 104713 13271 104771 13277
rect 105449 13311 105507 13317
rect 105449 13277 105461 13311
rect 105495 13277 105507 13311
rect 105449 13271 105507 13277
rect 105909 13311 105967 13317
rect 105909 13277 105921 13311
rect 105955 13277 105967 13311
rect 105909 13271 105967 13277
rect 100956 13212 104296 13240
rect 96948 13200 96954 13212
rect 86451 13144 86632 13172
rect 86451 13141 86463 13144
rect 86405 13135 86463 13141
rect 86678 13132 86684 13184
rect 86736 13172 86742 13184
rect 88886 13172 88892 13184
rect 86736 13144 88892 13172
rect 86736 13132 86742 13144
rect 88886 13132 88892 13144
rect 88944 13132 88950 13184
rect 88978 13132 88984 13184
rect 89036 13172 89042 13184
rect 89036 13144 89081 13172
rect 89036 13132 89042 13144
rect 91278 13132 91284 13184
rect 91336 13172 91342 13184
rect 94961 13175 95019 13181
rect 94961 13172 94973 13175
rect 91336 13144 94973 13172
rect 91336 13132 91342 13144
rect 94961 13141 94973 13144
rect 95007 13141 95019 13175
rect 94961 13135 95019 13141
rect 95050 13132 95056 13184
rect 95108 13172 95114 13184
rect 96706 13172 96712 13184
rect 95108 13144 96712 13172
rect 95108 13132 95114 13144
rect 96706 13132 96712 13144
rect 96764 13132 96770 13184
rect 96798 13132 96804 13184
rect 96856 13172 96862 13184
rect 98288 13172 98316 13212
rect 96856 13144 98316 13172
rect 96856 13132 96862 13144
rect 99006 13132 99012 13184
rect 99064 13172 99070 13184
rect 100849 13175 100907 13181
rect 100849 13172 100861 13175
rect 99064 13144 100861 13172
rect 99064 13132 99070 13144
rect 100849 13141 100861 13144
rect 100895 13141 100907 13175
rect 100849 13135 100907 13141
rect 102597 13175 102655 13181
rect 102597 13141 102609 13175
rect 102643 13172 102655 13175
rect 102962 13172 102968 13184
rect 102643 13144 102968 13172
rect 102643 13141 102655 13144
rect 102597 13135 102655 13141
rect 102962 13132 102968 13144
rect 103020 13132 103026 13184
rect 103054 13132 103060 13184
rect 103112 13172 103118 13184
rect 103793 13175 103851 13181
rect 103793 13172 103805 13175
rect 103112 13144 103805 13172
rect 103112 13132 103118 13144
rect 103793 13141 103805 13144
rect 103839 13141 103851 13175
rect 104728 13172 104756 13271
rect 105464 13240 105492 13271
rect 107010 13268 107016 13320
rect 107068 13308 107074 13320
rect 107657 13311 107715 13317
rect 107657 13308 107669 13311
rect 107068 13280 107669 13308
rect 107068 13268 107074 13280
rect 107657 13277 107669 13280
rect 107703 13277 107715 13311
rect 109034 13308 109040 13320
rect 107657 13271 107715 13277
rect 107764 13280 109040 13308
rect 107764 13240 107792 13280
rect 109034 13268 109040 13280
rect 109092 13308 109098 13320
rect 109678 13308 109684 13320
rect 109092 13280 109684 13308
rect 109092 13268 109098 13280
rect 109678 13268 109684 13280
rect 109736 13268 109742 13320
rect 109865 13311 109923 13317
rect 109865 13277 109877 13311
rect 109911 13308 109923 13311
rect 110046 13308 110052 13320
rect 109911 13280 110052 13308
rect 109911 13277 109923 13280
rect 109865 13271 109923 13277
rect 110046 13268 110052 13280
rect 110104 13268 110110 13320
rect 110601 13311 110659 13317
rect 110601 13277 110613 13311
rect 110647 13308 110659 13311
rect 111334 13308 111340 13320
rect 110647 13280 111196 13308
rect 111295 13280 111340 13308
rect 110647 13277 110659 13280
rect 110601 13271 110659 13277
rect 105464 13212 107792 13240
rect 107924 13243 107982 13249
rect 107924 13209 107936 13243
rect 107970 13240 107982 13243
rect 108574 13240 108580 13252
rect 107970 13212 108580 13240
rect 107970 13209 107982 13212
rect 107924 13203 107982 13209
rect 108574 13200 108580 13212
rect 108632 13200 108638 13252
rect 106366 13172 106372 13184
rect 104728 13144 106372 13172
rect 103793 13135 103851 13141
rect 106366 13132 106372 13144
rect 106424 13132 106430 13184
rect 109037 13175 109095 13181
rect 109037 13141 109049 13175
rect 109083 13172 109095 13175
rect 110414 13172 110420 13184
rect 109083 13144 110420 13172
rect 109083 13141 109095 13144
rect 109037 13135 109095 13141
rect 110414 13132 110420 13144
rect 110472 13132 110478 13184
rect 111168 13172 111196 13280
rect 111334 13268 111340 13280
rect 111392 13268 111398 13320
rect 112438 13308 112444 13320
rect 112399 13280 112444 13308
rect 112438 13268 112444 13280
rect 112496 13268 112502 13320
rect 112916 13317 112944 13348
rect 112990 13336 112996 13388
rect 113048 13376 113054 13388
rect 113048 13348 116256 13376
rect 113048 13336 113054 13348
rect 112907 13311 112965 13317
rect 112907 13277 112919 13311
rect 112953 13277 112965 13311
rect 112907 13271 112965 13277
rect 113913 13311 113971 13317
rect 113913 13277 113925 13311
rect 113959 13308 113971 13311
rect 114462 13308 114468 13320
rect 113959 13280 114468 13308
rect 113959 13277 113971 13280
rect 113913 13271 113971 13277
rect 114462 13268 114468 13280
rect 114520 13268 114526 13320
rect 114646 13268 114652 13320
rect 114704 13308 114710 13320
rect 114741 13311 114799 13317
rect 114741 13308 114753 13311
rect 114704 13280 114753 13308
rect 114704 13268 114710 13280
rect 114741 13277 114753 13280
rect 114787 13277 114799 13311
rect 114741 13271 114799 13277
rect 115658 13268 115664 13320
rect 115716 13308 115722 13320
rect 116228 13317 116256 13348
rect 117222 13336 117228 13388
rect 117280 13376 117286 13388
rect 117884 13376 117912 13416
rect 118881 13413 118893 13416
rect 118927 13413 118939 13447
rect 118881 13407 118939 13413
rect 119154 13404 119160 13456
rect 119212 13444 119218 13456
rect 120721 13447 120779 13453
rect 120721 13444 120733 13447
rect 119212 13416 120733 13444
rect 119212 13404 119218 13416
rect 120721 13413 120733 13416
rect 120767 13413 120779 13447
rect 120721 13407 120779 13413
rect 123849 13447 123907 13453
rect 123849 13413 123861 13447
rect 123895 13413 123907 13447
rect 123849 13407 123907 13413
rect 117280 13348 117912 13376
rect 117280 13336 117286 13348
rect 117958 13336 117964 13388
rect 118016 13376 118022 13388
rect 121362 13376 121368 13388
rect 118016 13348 121368 13376
rect 118016 13336 118022 13348
rect 121362 13336 121368 13348
rect 121420 13336 121426 13388
rect 122006 13336 122012 13388
rect 122064 13376 122070 13388
rect 122469 13379 122527 13385
rect 122469 13376 122481 13379
rect 122064 13348 122481 13376
rect 122064 13336 122070 13348
rect 122469 13345 122481 13348
rect 122515 13345 122527 13379
rect 122469 13339 122527 13345
rect 115753 13311 115811 13317
rect 115753 13308 115765 13311
rect 115716 13280 115765 13308
rect 115716 13268 115722 13280
rect 115753 13277 115765 13280
rect 115799 13277 115811 13311
rect 115753 13271 115811 13277
rect 116213 13311 116271 13317
rect 116213 13277 116225 13311
rect 116259 13277 116271 13311
rect 116213 13271 116271 13277
rect 116578 13268 116584 13320
rect 116636 13308 116642 13320
rect 116636 13280 117268 13308
rect 116636 13268 116642 13280
rect 112622 13200 112628 13252
rect 112680 13240 112686 13252
rect 112990 13240 112996 13252
rect 112680 13212 112996 13240
rect 112680 13200 112686 13212
rect 112990 13200 112996 13212
rect 113048 13200 113054 13252
rect 113082 13200 113088 13252
rect 113140 13240 113146 13252
rect 117130 13240 117136 13252
rect 113140 13212 117136 13240
rect 113140 13200 113146 13212
rect 117130 13200 117136 13212
rect 117188 13200 117194 13252
rect 117240 13240 117268 13280
rect 117314 13268 117320 13320
rect 117372 13308 117378 13320
rect 118329 13311 118387 13317
rect 117372 13280 117417 13308
rect 117372 13268 117378 13280
rect 118329 13277 118341 13311
rect 118375 13308 118387 13311
rect 119065 13311 119123 13317
rect 118375 13280 118694 13308
rect 118375 13277 118387 13280
rect 118329 13271 118387 13277
rect 118666 13240 118694 13280
rect 119065 13277 119077 13311
rect 119111 13308 119123 13311
rect 119890 13308 119896 13320
rect 119111 13280 119896 13308
rect 119111 13277 119123 13280
rect 119065 13271 119123 13277
rect 119890 13268 119896 13280
rect 119948 13268 119954 13320
rect 120169 13311 120227 13317
rect 120169 13277 120181 13311
rect 120215 13308 120227 13311
rect 120810 13308 120816 13320
rect 120215 13280 120816 13308
rect 120215 13277 120227 13280
rect 120169 13271 120227 13277
rect 120810 13268 120816 13280
rect 120868 13268 120874 13320
rect 120902 13268 120908 13320
rect 120960 13308 120966 13320
rect 121641 13311 121699 13317
rect 120960 13280 121005 13308
rect 120960 13268 120966 13280
rect 121641 13277 121653 13311
rect 121687 13308 121699 13311
rect 122098 13308 122104 13320
rect 121687 13280 122104 13308
rect 121687 13277 121699 13280
rect 121641 13271 121699 13277
rect 122098 13268 122104 13280
rect 122156 13268 122162 13320
rect 122736 13243 122794 13249
rect 117240 13212 117452 13240
rect 118666 13212 121408 13240
rect 113174 13172 113180 13184
rect 111168 13144 113180 13172
rect 113174 13132 113180 13144
rect 113232 13132 113238 13184
rect 114738 13132 114744 13184
rect 114796 13172 114802 13184
rect 115569 13175 115627 13181
rect 115569 13172 115581 13175
rect 114796 13144 115581 13172
rect 114796 13132 114802 13144
rect 115569 13141 115581 13144
rect 115615 13172 115627 13175
rect 117314 13172 117320 13184
rect 115615 13144 117320 13172
rect 115615 13141 115627 13144
rect 115569 13135 115627 13141
rect 117314 13132 117320 13144
rect 117372 13132 117378 13184
rect 117424 13172 117452 13212
rect 119154 13172 119160 13184
rect 117424 13144 119160 13172
rect 119154 13132 119160 13144
rect 119212 13132 119218 13184
rect 121380 13172 121408 13212
rect 122736 13209 122748 13243
rect 122782 13240 122794 13243
rect 123478 13240 123484 13252
rect 122782 13212 123484 13240
rect 122782 13209 122794 13212
rect 122736 13203 122794 13209
rect 123478 13200 123484 13212
rect 123536 13200 123542 13252
rect 123864 13240 123892 13407
rect 124674 13404 124680 13456
rect 124732 13444 124738 13456
rect 125873 13447 125931 13453
rect 125873 13444 125885 13447
rect 124732 13416 125885 13444
rect 124732 13404 124738 13416
rect 125873 13413 125885 13416
rect 125919 13413 125931 13447
rect 125873 13407 125931 13413
rect 126054 13404 126060 13456
rect 126112 13444 126118 13456
rect 127713 13447 127771 13453
rect 127713 13444 127725 13447
rect 126112 13416 127725 13444
rect 126112 13404 126118 13416
rect 127713 13413 127725 13416
rect 127759 13413 127771 13447
rect 127820 13444 127848 13484
rect 127986 13472 127992 13524
rect 128044 13512 128050 13524
rect 129185 13515 129243 13521
rect 129185 13512 129197 13515
rect 128044 13484 129197 13512
rect 128044 13472 128050 13484
rect 129185 13481 129197 13484
rect 129231 13481 129243 13515
rect 129185 13475 129243 13481
rect 129918 13472 129924 13524
rect 129976 13512 129982 13524
rect 131025 13515 131083 13521
rect 131025 13512 131037 13515
rect 129976 13484 131037 13512
rect 129976 13472 129982 13484
rect 131025 13481 131037 13484
rect 131071 13481 131083 13515
rect 131025 13475 131083 13481
rect 131114 13472 131120 13524
rect 131172 13512 131178 13524
rect 131761 13515 131819 13521
rect 131761 13512 131773 13515
rect 131172 13484 131773 13512
rect 131172 13472 131178 13484
rect 131761 13481 131773 13484
rect 131807 13481 131819 13515
rect 131761 13475 131819 13481
rect 132494 13472 132500 13524
rect 132552 13512 132558 13524
rect 132957 13515 133015 13521
rect 132957 13512 132969 13515
rect 132552 13484 132969 13512
rect 132552 13472 132558 13484
rect 132957 13481 132969 13484
rect 133003 13481 133015 13515
rect 132957 13475 133015 13481
rect 133230 13472 133236 13524
rect 133288 13512 133294 13524
rect 133288 13484 133920 13512
rect 133288 13472 133294 13484
rect 128449 13447 128507 13453
rect 128449 13444 128461 13447
rect 127820 13416 128461 13444
rect 127713 13407 127771 13413
rect 128449 13413 128461 13416
rect 128495 13413 128507 13447
rect 128449 13407 128507 13413
rect 128814 13404 128820 13456
rect 128872 13444 128878 13456
rect 130289 13447 130347 13453
rect 130289 13444 130301 13447
rect 128872 13416 130301 13444
rect 128872 13404 128878 13416
rect 130289 13413 130301 13416
rect 130335 13413 130347 13447
rect 130289 13407 130347 13413
rect 130488 13416 132632 13444
rect 124766 13336 124772 13388
rect 124824 13376 124830 13388
rect 125594 13376 125600 13388
rect 124824 13348 125600 13376
rect 124824 13336 124830 13348
rect 125594 13336 125600 13348
rect 125652 13336 125658 13388
rect 127434 13376 127440 13388
rect 126072 13348 127440 13376
rect 125318 13308 125324 13320
rect 125279 13280 125324 13308
rect 125318 13268 125324 13280
rect 125376 13268 125382 13320
rect 126072 13317 126100 13348
rect 127434 13336 127440 13348
rect 127492 13336 127498 13388
rect 127526 13336 127532 13388
rect 127584 13376 127590 13388
rect 130378 13376 130384 13388
rect 127584 13348 130384 13376
rect 127584 13336 127590 13348
rect 130378 13336 130384 13348
rect 130436 13336 130442 13388
rect 126057 13311 126115 13317
rect 126057 13277 126069 13311
rect 126103 13277 126115 13311
rect 126057 13271 126115 13277
rect 126793 13311 126851 13317
rect 126793 13277 126805 13311
rect 126839 13308 126851 13311
rect 127710 13308 127716 13320
rect 126839 13280 127716 13308
rect 126839 13277 126851 13280
rect 126793 13271 126851 13277
rect 127710 13268 127716 13280
rect 127768 13268 127774 13320
rect 127894 13308 127900 13320
rect 127855 13280 127900 13308
rect 127894 13268 127900 13280
rect 127952 13268 127958 13320
rect 128633 13311 128691 13317
rect 128633 13277 128645 13311
rect 128679 13308 128691 13311
rect 128722 13308 128728 13320
rect 128679 13280 128728 13308
rect 128679 13277 128691 13280
rect 128633 13271 128691 13277
rect 128722 13268 128728 13280
rect 128780 13268 128786 13320
rect 129369 13311 129427 13317
rect 129369 13277 129381 13311
rect 129415 13308 129427 13311
rect 130102 13308 130108 13320
rect 129415 13280 130108 13308
rect 129415 13277 129427 13280
rect 129369 13271 129427 13277
rect 130102 13268 130108 13280
rect 130160 13268 130166 13320
rect 130488 13317 130516 13416
rect 132604 13376 132632 13416
rect 132678 13404 132684 13456
rect 132736 13444 132742 13456
rect 133693 13447 133751 13453
rect 133693 13444 133705 13447
rect 132736 13416 133705 13444
rect 132736 13404 132742 13416
rect 133693 13413 133705 13416
rect 133739 13413 133751 13447
rect 133892 13444 133920 13484
rect 134334 13472 134340 13524
rect 134392 13512 134398 13524
rect 135441 13515 135499 13521
rect 135441 13512 135453 13515
rect 134392 13484 135453 13512
rect 134392 13472 134398 13484
rect 135441 13481 135453 13484
rect 135487 13481 135499 13515
rect 135441 13475 135499 13481
rect 135714 13472 135720 13524
rect 135772 13512 135778 13524
rect 136269 13515 136327 13521
rect 136269 13512 136281 13515
rect 135772 13484 136281 13512
rect 135772 13472 135778 13484
rect 136269 13481 136281 13484
rect 136315 13481 136327 13515
rect 136269 13475 136327 13481
rect 136358 13472 136364 13524
rect 136416 13512 136422 13524
rect 137005 13515 137063 13521
rect 137005 13512 137017 13515
rect 136416 13484 137017 13512
rect 136416 13472 136422 13484
rect 137005 13481 137017 13484
rect 137051 13481 137063 13515
rect 137005 13475 137063 13481
rect 137094 13472 137100 13524
rect 137152 13512 137158 13524
rect 138017 13515 138075 13521
rect 138017 13512 138029 13515
rect 137152 13484 138029 13512
rect 137152 13472 137158 13484
rect 138017 13481 138029 13484
rect 138063 13481 138075 13515
rect 138017 13475 138075 13481
rect 138198 13472 138204 13524
rect 138256 13512 138262 13524
rect 138753 13515 138811 13521
rect 138753 13512 138765 13515
rect 138256 13484 138765 13512
rect 138256 13472 138262 13484
rect 138753 13481 138765 13484
rect 138799 13481 138811 13515
rect 138753 13475 138811 13481
rect 138842 13472 138848 13524
rect 138900 13512 138906 13524
rect 139581 13515 139639 13521
rect 139581 13512 139593 13515
rect 138900 13484 139593 13512
rect 138900 13472 138906 13484
rect 139581 13481 139593 13484
rect 139627 13481 139639 13515
rect 139581 13475 139639 13481
rect 139854 13472 139860 13524
rect 139912 13512 139918 13524
rect 140593 13515 140651 13521
rect 140593 13512 140605 13515
rect 139912 13484 140605 13512
rect 139912 13472 139918 13484
rect 140593 13481 140605 13484
rect 140639 13481 140651 13515
rect 140593 13475 140651 13481
rect 140682 13472 140688 13524
rect 140740 13512 140746 13524
rect 141421 13515 141479 13521
rect 141421 13512 141433 13515
rect 140740 13484 141433 13512
rect 140740 13472 140746 13484
rect 141421 13481 141433 13484
rect 141467 13481 141479 13515
rect 141421 13475 141479 13481
rect 141510 13472 141516 13524
rect 141568 13512 141574 13524
rect 141568 13484 142292 13512
rect 141568 13472 141574 13484
rect 134429 13447 134487 13453
rect 134429 13444 134441 13447
rect 133892 13416 134441 13444
rect 133693 13407 133751 13413
rect 134429 13413 134441 13416
rect 134475 13413 134487 13447
rect 138382 13444 138388 13456
rect 134429 13407 134487 13413
rect 135226 13416 138388 13444
rect 135226 13376 135254 13416
rect 138382 13404 138388 13416
rect 138440 13404 138446 13456
rect 138566 13404 138572 13456
rect 138624 13444 138630 13456
rect 141142 13444 141148 13456
rect 138624 13416 141148 13444
rect 138624 13404 138630 13416
rect 141142 13404 141148 13416
rect 141200 13404 141206 13456
rect 141234 13404 141240 13456
rect 141292 13444 141298 13456
rect 142157 13447 142215 13453
rect 142157 13444 142169 13447
rect 141292 13416 142169 13444
rect 141292 13404 141298 13416
rect 142157 13413 142169 13416
rect 142203 13413 142215 13447
rect 142264 13444 142292 13484
rect 142522 13472 142528 13524
rect 142580 13512 142586 13524
rect 147309 13515 147367 13521
rect 142580 13484 147260 13512
rect 142580 13472 142586 13484
rect 147232 13444 147260 13484
rect 147309 13481 147321 13515
rect 147355 13512 147367 13515
rect 148042 13512 148048 13524
rect 147355 13484 148048 13512
rect 147355 13481 147367 13484
rect 147309 13475 147367 13481
rect 148042 13472 148048 13484
rect 148100 13472 148106 13524
rect 148594 13472 148600 13524
rect 148652 13512 148658 13524
rect 149882 13512 149888 13524
rect 148652 13484 149888 13512
rect 148652 13472 148658 13484
rect 149882 13472 149888 13484
rect 149940 13472 149946 13524
rect 151262 13512 151268 13524
rect 149992 13484 151268 13512
rect 147398 13444 147404 13456
rect 142264 13416 143212 13444
rect 147232 13416 147404 13444
rect 142157 13407 142215 13413
rect 131868 13348 132356 13376
rect 132604 13348 135254 13376
rect 130473 13311 130531 13317
rect 130473 13277 130485 13311
rect 130519 13277 130531 13311
rect 130473 13271 130531 13277
rect 131209 13311 131267 13317
rect 131209 13277 131221 13311
rect 131255 13308 131267 13311
rect 131868 13308 131896 13348
rect 131255 13280 131896 13308
rect 131255 13277 131267 13280
rect 131209 13271 131267 13277
rect 131942 13268 131948 13320
rect 132000 13308 132006 13320
rect 132328 13308 132356 13348
rect 135346 13336 135352 13388
rect 135404 13376 135410 13388
rect 135404 13348 136220 13376
rect 135404 13336 135410 13348
rect 132402 13308 132408 13320
rect 132000 13280 132045 13308
rect 132328 13280 132408 13308
rect 132000 13268 132006 13280
rect 132402 13268 132408 13280
rect 132460 13268 132466 13320
rect 132773 13311 132831 13317
rect 132773 13277 132785 13311
rect 132819 13277 132831 13311
rect 133509 13311 133567 13317
rect 133509 13308 133521 13311
rect 132773 13271 132831 13277
rect 132880 13280 133521 13308
rect 132788 13240 132816 13271
rect 123864 13212 132816 13240
rect 124306 13172 124312 13184
rect 121380 13144 124312 13172
rect 124306 13132 124312 13144
rect 124364 13132 124370 13184
rect 124398 13132 124404 13184
rect 124456 13172 124462 13184
rect 128630 13172 128636 13184
rect 124456 13144 128636 13172
rect 124456 13132 124462 13144
rect 128630 13132 128636 13144
rect 128688 13132 128694 13184
rect 128814 13132 128820 13184
rect 128872 13172 128878 13184
rect 129090 13172 129096 13184
rect 128872 13144 129096 13172
rect 128872 13132 128878 13144
rect 129090 13132 129096 13144
rect 129148 13132 129154 13184
rect 131206 13132 131212 13184
rect 131264 13172 131270 13184
rect 132880 13172 132908 13280
rect 133509 13277 133521 13280
rect 133555 13277 133567 13311
rect 133509 13271 133567 13277
rect 133874 13268 133880 13320
rect 133932 13308 133938 13320
rect 134245 13311 134303 13317
rect 134245 13308 134257 13311
rect 133932 13280 134257 13308
rect 133932 13268 133938 13280
rect 134245 13277 134257 13280
rect 134291 13277 134303 13311
rect 135622 13308 135628 13320
rect 135583 13280 135628 13308
rect 134245 13271 134303 13277
rect 135622 13268 135628 13280
rect 135680 13268 135686 13320
rect 136082 13308 136088 13320
rect 136043 13280 136088 13308
rect 136082 13268 136088 13280
rect 136140 13268 136146 13320
rect 136192 13308 136220 13348
rect 136726 13336 136732 13388
rect 136784 13376 136790 13388
rect 143077 13379 143135 13385
rect 143077 13376 143089 13379
rect 136784 13348 143089 13376
rect 136784 13336 136790 13348
rect 136821 13311 136879 13317
rect 136821 13308 136833 13311
rect 136192 13280 136833 13308
rect 136821 13277 136833 13280
rect 136867 13277 136879 13311
rect 136821 13271 136879 13277
rect 138106 13268 138112 13320
rect 138164 13308 138170 13320
rect 138952 13317 138980 13348
rect 143077 13345 143089 13348
rect 143123 13345 143135 13379
rect 143077 13339 143135 13345
rect 138201 13311 138259 13317
rect 138201 13308 138213 13311
rect 138164 13280 138213 13308
rect 138164 13268 138170 13280
rect 138201 13277 138213 13280
rect 138247 13277 138259 13311
rect 138201 13271 138259 13277
rect 138937 13311 138995 13317
rect 138937 13277 138949 13311
rect 138983 13277 138995 13311
rect 139394 13308 139400 13320
rect 139355 13280 139400 13308
rect 138937 13271 138995 13277
rect 139394 13268 139400 13280
rect 139452 13268 139458 13320
rect 140774 13308 140780 13320
rect 140735 13280 140780 13308
rect 140774 13268 140780 13280
rect 140832 13268 140838 13320
rect 140866 13268 140872 13320
rect 140924 13308 140930 13320
rect 141237 13311 141295 13317
rect 141237 13308 141249 13311
rect 140924 13280 141249 13308
rect 140924 13268 140930 13280
rect 141237 13277 141249 13280
rect 141283 13277 141295 13311
rect 141237 13271 141295 13277
rect 141973 13311 142031 13317
rect 141973 13277 141985 13311
rect 142019 13277 142031 13311
rect 141973 13271 142031 13277
rect 133598 13200 133604 13252
rect 133656 13240 133662 13252
rect 139578 13240 139584 13252
rect 133656 13212 139584 13240
rect 133656 13200 133662 13212
rect 139578 13200 139584 13212
rect 139636 13200 139642 13252
rect 139670 13200 139676 13252
rect 139728 13240 139734 13252
rect 141988 13240 142016 13271
rect 139728 13212 142016 13240
rect 143184 13240 143212 13416
rect 147398 13404 147404 13416
rect 147456 13404 147462 13456
rect 148134 13444 148140 13456
rect 147646 13416 148140 13444
rect 146938 13336 146944 13388
rect 146996 13376 147002 13388
rect 147646 13376 147674 13416
rect 148134 13404 148140 13416
rect 148192 13404 148198 13456
rect 149609 13447 149667 13453
rect 149609 13413 149621 13447
rect 149655 13444 149667 13447
rect 149992 13444 150020 13484
rect 151262 13472 151268 13484
rect 151320 13472 151326 13524
rect 151814 13472 151820 13524
rect 151872 13512 151878 13524
rect 151872 13484 152228 13512
rect 151872 13472 151878 13484
rect 149655 13416 150020 13444
rect 150069 13447 150127 13453
rect 149655 13413 149667 13416
rect 149609 13407 149667 13413
rect 150069 13413 150081 13447
rect 150115 13413 150127 13447
rect 150802 13444 150808 13456
rect 150763 13416 150808 13444
rect 150069 13407 150127 13413
rect 146996 13348 147674 13376
rect 146996 13336 147002 13348
rect 149238 13336 149244 13388
rect 149296 13376 149302 13388
rect 150084 13376 150112 13407
rect 150802 13404 150808 13416
rect 150860 13404 150866 13456
rect 152200 13444 152228 13484
rect 153562 13472 153568 13524
rect 153620 13512 153626 13524
rect 154298 13512 154304 13524
rect 153620 13484 153665 13512
rect 154259 13484 154304 13512
rect 153620 13472 153626 13484
rect 154298 13472 154304 13484
rect 154356 13472 154362 13524
rect 155862 13472 155868 13524
rect 155920 13512 155926 13524
rect 156141 13515 156199 13521
rect 156141 13512 156153 13515
rect 155920 13484 156153 13512
rect 155920 13472 155926 13484
rect 156141 13481 156153 13484
rect 156187 13481 156199 13515
rect 156141 13475 156199 13481
rect 155678 13444 155684 13456
rect 152200 13416 155684 13444
rect 155678 13404 155684 13416
rect 155736 13404 155742 13456
rect 155770 13404 155776 13456
rect 155828 13444 155834 13456
rect 156877 13447 156935 13453
rect 156877 13444 156889 13447
rect 155828 13416 156889 13444
rect 155828 13404 155834 13416
rect 156877 13413 156889 13416
rect 156923 13413 156935 13447
rect 156877 13407 156935 13413
rect 149296 13348 150112 13376
rect 149296 13336 149302 13348
rect 152366 13336 152372 13388
rect 152424 13376 152430 13388
rect 156782 13376 156788 13388
rect 152424 13348 156788 13376
rect 152424 13336 152430 13348
rect 156782 13336 156788 13348
rect 156840 13336 156846 13388
rect 143350 13268 143356 13320
rect 143408 13308 143414 13320
rect 143721 13311 143779 13317
rect 143721 13308 143733 13311
rect 143408 13280 143733 13308
rect 143408 13268 143414 13280
rect 143721 13277 143733 13280
rect 143767 13308 143779 13311
rect 145929 13311 145987 13317
rect 145929 13308 145941 13311
rect 143767 13280 145941 13308
rect 143767 13277 143779 13280
rect 143721 13271 143779 13277
rect 145929 13277 145941 13280
rect 145975 13308 145987 13311
rect 147490 13308 147496 13320
rect 145975 13280 147496 13308
rect 145975 13277 145987 13280
rect 145929 13271 145987 13277
rect 147490 13268 147496 13280
rect 147548 13308 147554 13320
rect 148229 13311 148287 13317
rect 148229 13308 148241 13311
rect 147548 13280 148241 13308
rect 147548 13268 147554 13280
rect 148229 13277 148241 13280
rect 148275 13308 148287 13311
rect 150253 13311 150311 13317
rect 148275 13280 149376 13308
rect 148275 13277 148287 13280
rect 148229 13271 148287 13277
rect 143994 13249 144000 13252
rect 143988 13240 144000 13249
rect 143184 13212 144000 13240
rect 139728 13200 139734 13212
rect 143988 13203 144000 13212
rect 143994 13200 144000 13203
rect 144052 13200 144058 13252
rect 145834 13240 145840 13252
rect 144104 13212 145840 13240
rect 131264 13144 132908 13172
rect 131264 13132 131270 13144
rect 133138 13132 133144 13184
rect 133196 13172 133202 13184
rect 135162 13172 135168 13184
rect 133196 13144 135168 13172
rect 133196 13132 133202 13144
rect 135162 13132 135168 13144
rect 135220 13132 135226 13184
rect 135530 13132 135536 13184
rect 135588 13172 135594 13184
rect 142706 13172 142712 13184
rect 135588 13144 142712 13172
rect 135588 13132 135594 13144
rect 142706 13132 142712 13144
rect 142764 13132 142770 13184
rect 143810 13132 143816 13184
rect 143868 13172 143874 13184
rect 144104 13172 144132 13212
rect 145834 13200 145840 13212
rect 145892 13200 145898 13252
rect 146202 13249 146208 13252
rect 146196 13240 146208 13249
rect 146163 13212 146208 13240
rect 146196 13203 146208 13212
rect 146202 13200 146208 13203
rect 146260 13200 146266 13252
rect 146478 13200 146484 13252
rect 146536 13240 146542 13252
rect 148496 13243 148554 13249
rect 146536 13212 148456 13240
rect 146536 13200 146542 13212
rect 145098 13172 145104 13184
rect 143868 13144 144132 13172
rect 145059 13144 145104 13172
rect 143868 13132 143874 13144
rect 145098 13132 145104 13144
rect 145156 13132 145162 13184
rect 148428 13172 148456 13212
rect 148496 13209 148508 13243
rect 148542 13240 148554 13243
rect 148594 13240 148600 13252
rect 148542 13212 148600 13240
rect 148542 13209 148554 13212
rect 148496 13203 148554 13209
rect 148594 13200 148600 13212
rect 148652 13200 148658 13252
rect 149238 13240 149244 13252
rect 148704 13212 149244 13240
rect 148704 13172 148732 13212
rect 149238 13200 149244 13212
rect 149296 13200 149302 13252
rect 149348 13240 149376 13280
rect 150253 13277 150265 13311
rect 150299 13308 150311 13311
rect 150894 13308 150900 13320
rect 150299 13280 150900 13308
rect 150299 13277 150311 13280
rect 150253 13271 150311 13277
rect 150894 13268 150900 13280
rect 150952 13268 150958 13320
rect 152185 13311 152243 13317
rect 151004 13280 152044 13308
rect 151004 13240 151032 13280
rect 149348 13212 151032 13240
rect 151918 13243 151976 13249
rect 151918 13209 151930 13243
rect 151964 13209 151976 13243
rect 152016 13240 152044 13280
rect 152185 13277 152197 13311
rect 152231 13308 152243 13311
rect 152458 13308 152464 13320
rect 152231 13280 152464 13308
rect 152231 13277 152243 13280
rect 152185 13271 152243 13277
rect 152458 13268 152464 13280
rect 152516 13268 152522 13320
rect 152826 13308 152832 13320
rect 152787 13280 152832 13308
rect 152826 13268 152832 13280
rect 152884 13268 152890 13320
rect 153378 13308 153384 13320
rect 153339 13280 153384 13308
rect 153378 13268 153384 13280
rect 153436 13268 153442 13320
rect 153470 13268 153476 13320
rect 153528 13308 153534 13320
rect 154117 13311 154175 13317
rect 154117 13308 154129 13311
rect 153528 13280 154129 13308
rect 153528 13268 153534 13280
rect 154117 13277 154129 13280
rect 154163 13277 154175 13311
rect 154850 13308 154856 13320
rect 154811 13280 154856 13308
rect 154117 13271 154175 13277
rect 154850 13268 154856 13280
rect 154908 13268 154914 13320
rect 155954 13308 155960 13320
rect 155915 13280 155960 13308
rect 155954 13268 155960 13280
rect 156012 13268 156018 13320
rect 156690 13308 156696 13320
rect 156651 13280 156696 13308
rect 156690 13268 156696 13280
rect 156748 13268 156754 13320
rect 157426 13308 157432 13320
rect 157387 13280 157432 13308
rect 157426 13268 157432 13280
rect 157484 13268 157490 13320
rect 152734 13240 152740 13252
rect 152016 13212 152740 13240
rect 151918 13203 151976 13209
rect 148428 13144 148732 13172
rect 149146 13132 149152 13184
rect 149204 13172 149210 13184
rect 151814 13172 151820 13184
rect 149204 13144 151820 13172
rect 149204 13132 149210 13144
rect 151814 13132 151820 13144
rect 151872 13172 151878 13184
rect 151933 13172 151961 13203
rect 152734 13200 152740 13212
rect 152792 13200 152798 13252
rect 153286 13200 153292 13252
rect 153344 13240 153350 13252
rect 153344 13212 157656 13240
rect 153344 13200 153350 13212
rect 151872 13144 151961 13172
rect 151872 13132 151878 13144
rect 152366 13132 152372 13184
rect 152424 13172 152430 13184
rect 152645 13175 152703 13181
rect 152645 13172 152657 13175
rect 152424 13144 152657 13172
rect 152424 13132 152430 13144
rect 152645 13141 152657 13144
rect 152691 13141 152703 13175
rect 152645 13135 152703 13141
rect 153194 13132 153200 13184
rect 153252 13172 153258 13184
rect 153746 13172 153752 13184
rect 153252 13144 153752 13172
rect 153252 13132 153258 13144
rect 153746 13132 153752 13144
rect 153804 13172 153810 13184
rect 154206 13172 154212 13184
rect 153804 13144 154212 13172
rect 153804 13132 153810 13144
rect 154206 13132 154212 13144
rect 154264 13132 154270 13184
rect 154390 13132 154396 13184
rect 154448 13172 154454 13184
rect 157628 13181 157656 13212
rect 155037 13175 155095 13181
rect 155037 13172 155049 13175
rect 154448 13144 155049 13172
rect 154448 13132 154454 13144
rect 155037 13141 155049 13144
rect 155083 13141 155095 13175
rect 155037 13135 155095 13141
rect 157613 13175 157671 13181
rect 157613 13141 157625 13175
rect 157659 13141 157671 13175
rect 157613 13135 157671 13141
rect 1104 13082 159043 13104
rect 1104 13030 40394 13082
rect 40446 13030 40458 13082
rect 40510 13030 40522 13082
rect 40574 13030 40586 13082
rect 40638 13030 40650 13082
rect 40702 13030 79839 13082
rect 79891 13030 79903 13082
rect 79955 13030 79967 13082
rect 80019 13030 80031 13082
rect 80083 13030 80095 13082
rect 80147 13030 119284 13082
rect 119336 13030 119348 13082
rect 119400 13030 119412 13082
rect 119464 13030 119476 13082
rect 119528 13030 119540 13082
rect 119592 13030 158729 13082
rect 158781 13030 158793 13082
rect 158845 13030 158857 13082
rect 158909 13030 158921 13082
rect 158973 13030 158985 13082
rect 159037 13030 159043 13082
rect 1104 13008 159043 13030
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 9398 12968 9404 12980
rect 7331 12940 9404 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 10134 12968 10140 12980
rect 9539 12940 10140 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 11790 12968 11796 12980
rect 10275 12940 11796 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12032 12940 13584 12968
rect 12032 12928 12038 12940
rect 13556 12900 13584 12940
rect 13906 12928 13912 12980
rect 13964 12968 13970 12980
rect 15010 12968 15016 12980
rect 13964 12940 15016 12968
rect 13964 12928 13970 12940
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15562 12968 15568 12980
rect 15475 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12968 15626 12980
rect 15746 12968 15752 12980
rect 15620 12940 15752 12968
rect 15620 12928 15626 12940
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12968 16175 12971
rect 16758 12968 16764 12980
rect 16163 12940 16764 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 18690 12968 18696 12980
rect 18651 12940 18696 12968
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 19429 12971 19487 12977
rect 19429 12937 19441 12971
rect 19475 12968 19487 12971
rect 20070 12968 20076 12980
rect 19475 12940 20076 12968
rect 19475 12937 19487 12940
rect 19429 12931 19487 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 22649 12971 22707 12977
rect 20220 12940 22600 12968
rect 20220 12928 20226 12940
rect 14746 12903 14804 12909
rect 14746 12900 14758 12903
rect 9692 12872 12940 12900
rect 13556 12872 14758 12900
rect 9692 12841 9720 12872
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 9677 12795 9735 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10870 12832 10876 12844
rect 10831 12804 10876 12832
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 11974 12832 11980 12844
rect 11931 12804 11980 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 10778 12764 10784 12776
rect 8987 12736 10784 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 10962 12724 10968 12776
rect 11020 12764 11026 12776
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 11020 12736 11713 12764
rect 11020 12724 11026 12736
rect 11701 12733 11713 12736
rect 11747 12764 11759 12767
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 11747 12736 12817 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12912 12764 12940 12872
rect 14746 12869 14758 12872
rect 14792 12869 14804 12903
rect 15838 12900 15844 12912
rect 14746 12863 14804 12869
rect 14844 12872 15844 12900
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 14844 12832 14872 12872
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 22572 12900 22600 12940
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 23382 12968 23388 12980
rect 22695 12940 23388 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 23477 12971 23535 12977
rect 23477 12937 23489 12971
rect 23523 12968 23535 12971
rect 24762 12968 24768 12980
rect 23523 12940 24768 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 26234 12968 26240 12980
rect 25096 12940 26240 12968
rect 25096 12928 25102 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 26418 12968 26424 12980
rect 26379 12940 26424 12968
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 26786 12968 26792 12980
rect 26528 12940 26792 12968
rect 26528 12900 26556 12940
rect 26786 12928 26792 12940
rect 26844 12928 26850 12980
rect 31386 12968 31392 12980
rect 27540 12940 31392 12968
rect 16316 12872 18828 12900
rect 16316 12841 16344 12872
rect 13035 12804 14872 12832
rect 16301 12835 16359 12841
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 16301 12801 16313 12835
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 17736 12804 17781 12832
rect 17736 12792 17742 12804
rect 15010 12764 15016 12776
rect 12912 12736 13768 12764
rect 14971 12736 15016 12764
rect 12805 12727 12863 12733
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12696 8447 12699
rect 10042 12696 10048 12708
rect 8435 12668 10048 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 11057 12699 11115 12705
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 13446 12696 13452 12708
rect 11103 12668 13452 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 7837 12631 7895 12637
rect 7837 12597 7849 12631
rect 7883 12628 7895 12631
rect 11882 12628 11888 12640
rect 7883 12600 11888 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12342 12628 12348 12640
rect 12115 12600 12348 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 13136 12600 13185 12628
rect 13136 12588 13142 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 13173 12591 13231 12597
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13633 12631 13691 12637
rect 13633 12628 13645 12631
rect 13412 12600 13645 12628
rect 13412 12588 13418 12600
rect 13633 12597 13645 12600
rect 13679 12597 13691 12631
rect 13740 12628 13768 12736
rect 15010 12724 15016 12736
rect 15068 12764 15074 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15068 12736 16865 12764
rect 15068 12724 15074 12736
rect 16853 12733 16865 12736
rect 16899 12764 16911 12767
rect 17218 12764 17224 12776
rect 16899 12736 17224 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 17696 12696 17724 12792
rect 18800 12764 18828 12872
rect 18892 12872 19564 12900
rect 18892 12841 18920 12872
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19150 12764 19156 12776
rect 18800 12736 19156 12764
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19536 12764 19564 12872
rect 19628 12872 22508 12900
rect 22572 12872 26556 12900
rect 19628 12841 19656 12872
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 21197 12835 21255 12841
rect 21197 12801 21209 12835
rect 21243 12832 21255 12835
rect 22186 12832 22192 12844
rect 21243 12804 22192 12832
rect 21243 12801 21255 12804
rect 21197 12795 21255 12801
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 22480 12832 22508 12872
rect 22738 12832 22744 12844
rect 22480 12804 22744 12832
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23014 12832 23020 12844
rect 22879 12804 23020 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 25153 12835 25211 12841
rect 25153 12801 25165 12835
rect 25199 12832 25211 12835
rect 25682 12832 25688 12844
rect 25199 12804 25688 12832
rect 25199 12801 25211 12804
rect 25153 12795 25211 12801
rect 19794 12764 19800 12776
rect 19536 12736 19800 12764
rect 19794 12724 19800 12736
rect 19852 12724 19858 12776
rect 21450 12764 21456 12776
rect 21411 12736 21456 12764
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 23308 12764 23336 12795
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 27540 12832 27568 12940
rect 31386 12928 31392 12940
rect 31444 12928 31450 12980
rect 32306 12968 32312 12980
rect 31516 12940 32312 12968
rect 26651 12804 27568 12832
rect 27724 12872 28764 12900
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 22152 12736 23336 12764
rect 22152 12724 22158 12736
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 26142 12764 26148 12776
rect 25464 12736 26148 12764
rect 25464 12724 25470 12736
rect 26142 12724 26148 12736
rect 26200 12764 26206 12776
rect 27724 12764 27752 12872
rect 28638 12835 28696 12841
rect 28638 12832 28650 12835
rect 26200 12736 27752 12764
rect 27908 12804 28650 12832
rect 26200 12724 26206 12736
rect 22370 12696 22376 12708
rect 17696 12668 20208 12696
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 13740 12600 20085 12628
rect 13633 12591 13691 12597
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 20180 12628 20208 12668
rect 21468 12668 22376 12696
rect 21468 12628 21496 12668
rect 22370 12656 22376 12668
rect 22428 12656 22434 12708
rect 24026 12696 24032 12708
rect 23987 12668 24032 12696
rect 24026 12656 24032 12668
rect 24084 12656 24090 12708
rect 25590 12656 25596 12708
rect 25648 12696 25654 12708
rect 25648 12668 27660 12696
rect 25648 12656 25654 12668
rect 20180 12600 21496 12628
rect 22097 12631 22155 12637
rect 20073 12591 20131 12597
rect 22097 12597 22109 12631
rect 22143 12628 22155 12631
rect 23750 12628 23756 12640
rect 22143 12600 23756 12628
rect 22143 12597 22155 12600
rect 22097 12591 22155 12597
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 27430 12588 27436 12640
rect 27488 12628 27494 12640
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 27488 12600 27537 12628
rect 27488 12588 27494 12600
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27632 12628 27660 12668
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 27908 12696 27936 12804
rect 28638 12801 28650 12804
rect 28684 12801 28696 12835
rect 28736 12832 28764 12872
rect 28810 12860 28816 12912
rect 28868 12900 28874 12912
rect 31516 12909 31544 12940
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 32490 12968 32496 12980
rect 32451 12940 32496 12968
rect 32490 12928 32496 12940
rect 32548 12928 32554 12980
rect 33502 12968 33508 12980
rect 33463 12940 33508 12968
rect 33502 12928 33508 12940
rect 33560 12928 33566 12980
rect 36538 12968 36544 12980
rect 33980 12940 36544 12968
rect 31512 12903 31570 12909
rect 28868 12872 29868 12900
rect 28868 12860 28874 12872
rect 28905 12835 28963 12841
rect 28905 12832 28917 12835
rect 28736 12804 28917 12832
rect 28638 12795 28696 12801
rect 28905 12801 28917 12804
rect 28951 12832 28963 12835
rect 28994 12832 29000 12844
rect 28951 12804 29000 12832
rect 28951 12801 28963 12804
rect 28905 12795 28963 12801
rect 28994 12792 29000 12804
rect 29052 12792 29058 12844
rect 29641 12835 29699 12841
rect 29641 12801 29653 12835
rect 29687 12801 29699 12835
rect 29840 12832 29868 12872
rect 31512 12869 31524 12903
rect 31558 12869 31570 12903
rect 31512 12863 31570 12869
rect 31754 12860 31760 12912
rect 31812 12900 31818 12912
rect 31812 12872 32352 12900
rect 31812 12860 31818 12872
rect 32324 12841 32352 12872
rect 32309 12835 32367 12841
rect 29840 12804 32260 12832
rect 29641 12795 29699 12801
rect 27764 12668 27936 12696
rect 27764 12656 27770 12668
rect 29656 12628 29684 12795
rect 31757 12767 31815 12773
rect 31757 12733 31769 12767
rect 31803 12764 31815 12767
rect 32030 12764 32036 12776
rect 31803 12736 32036 12764
rect 31803 12733 31815 12736
rect 31757 12727 31815 12733
rect 32030 12724 32036 12736
rect 32088 12724 32094 12776
rect 32232 12764 32260 12804
rect 32309 12801 32321 12835
rect 32355 12801 32367 12835
rect 33686 12832 33692 12844
rect 33647 12804 33692 12832
rect 32309 12795 32367 12801
rect 33686 12792 33692 12804
rect 33744 12792 33750 12844
rect 33980 12764 34008 12940
rect 36538 12928 36544 12940
rect 36596 12928 36602 12980
rect 36630 12928 36636 12980
rect 36688 12968 36694 12980
rect 36817 12971 36875 12977
rect 36817 12968 36829 12971
rect 36688 12940 36829 12968
rect 36688 12928 36694 12940
rect 36817 12937 36829 12940
rect 36863 12937 36875 12971
rect 36817 12931 36875 12937
rect 37734 12928 37740 12980
rect 37792 12968 37798 12980
rect 37921 12971 37979 12977
rect 37921 12968 37933 12971
rect 37792 12940 37933 12968
rect 37792 12928 37798 12940
rect 37921 12937 37933 12940
rect 37967 12937 37979 12971
rect 37921 12931 37979 12937
rect 38565 12971 38623 12977
rect 38565 12937 38577 12971
rect 38611 12968 38623 12971
rect 38838 12968 38844 12980
rect 38611 12940 38844 12968
rect 38611 12937 38623 12940
rect 38565 12931 38623 12937
rect 38838 12928 38844 12940
rect 38896 12928 38902 12980
rect 39393 12971 39451 12977
rect 39393 12937 39405 12971
rect 39439 12968 39451 12971
rect 41598 12968 41604 12980
rect 39439 12940 41604 12968
rect 39439 12937 39451 12940
rect 39393 12931 39451 12937
rect 41598 12928 41604 12940
rect 41656 12928 41662 12980
rect 43806 12968 43812 12980
rect 41892 12940 43812 12968
rect 34146 12860 34152 12912
rect 34204 12900 34210 12912
rect 34394 12903 34452 12909
rect 34394 12900 34406 12903
rect 34204 12872 34406 12900
rect 34204 12860 34210 12872
rect 34394 12869 34406 12872
rect 34440 12869 34452 12903
rect 34394 12863 34452 12869
rect 35434 12860 35440 12912
rect 35492 12900 35498 12912
rect 35492 12872 39252 12900
rect 35492 12860 35498 12872
rect 36633 12835 36691 12841
rect 36633 12832 36645 12835
rect 32232 12736 34008 12764
rect 34072 12804 36645 12832
rect 29730 12656 29736 12708
rect 29788 12696 29794 12708
rect 30377 12699 30435 12705
rect 30377 12696 30389 12699
rect 29788 12668 30389 12696
rect 29788 12656 29794 12668
rect 30377 12665 30389 12668
rect 30423 12665 30435 12699
rect 30377 12659 30435 12665
rect 29822 12628 29828 12640
rect 27632 12600 29684 12628
rect 29783 12600 29828 12628
rect 27525 12591 27583 12597
rect 29822 12588 29828 12600
rect 29880 12588 29886 12640
rect 31386 12588 31392 12640
rect 31444 12628 31450 12640
rect 34072 12628 34100 12804
rect 36633 12801 36645 12804
rect 36679 12801 36691 12835
rect 36633 12795 36691 12801
rect 36722 12792 36728 12844
rect 36780 12832 36786 12844
rect 37737 12835 37795 12841
rect 37737 12832 37749 12835
rect 36780 12804 37749 12832
rect 36780 12792 36786 12804
rect 37737 12801 37749 12804
rect 37783 12801 37795 12835
rect 37737 12795 37795 12801
rect 37826 12792 37832 12844
rect 37884 12832 37890 12844
rect 39224 12841 39252 12872
rect 39960 12872 41414 12900
rect 38749 12835 38807 12841
rect 37884 12804 38700 12832
rect 37884 12792 37890 12804
rect 34149 12767 34207 12773
rect 34149 12733 34161 12767
rect 34195 12733 34207 12767
rect 34149 12727 34207 12733
rect 31444 12600 34100 12628
rect 34164 12628 34192 12727
rect 35342 12724 35348 12776
rect 35400 12764 35406 12776
rect 35400 12736 38516 12764
rect 35400 12724 35406 12736
rect 35529 12699 35587 12705
rect 35529 12665 35541 12699
rect 35575 12696 35587 12699
rect 38378 12696 38384 12708
rect 35575 12668 38384 12696
rect 35575 12665 35587 12668
rect 35529 12659 35587 12665
rect 38378 12656 38384 12668
rect 38436 12656 38442 12708
rect 34422 12628 34428 12640
rect 34164 12600 34428 12628
rect 31444 12588 31450 12600
rect 34422 12588 34428 12600
rect 34480 12588 34486 12640
rect 36173 12631 36231 12637
rect 36173 12597 36185 12631
rect 36219 12628 36231 12631
rect 36262 12628 36268 12640
rect 36219 12600 36268 12628
rect 36219 12597 36231 12600
rect 36173 12591 36231 12597
rect 36262 12588 36268 12600
rect 36320 12588 36326 12640
rect 38488 12628 38516 12736
rect 38672 12696 38700 12804
rect 38749 12801 38761 12835
rect 38795 12801 38807 12835
rect 38749 12795 38807 12801
rect 39209 12835 39267 12841
rect 39209 12801 39221 12835
rect 39255 12801 39267 12835
rect 39209 12795 39267 12801
rect 38764 12764 38792 12795
rect 39850 12764 39856 12776
rect 38764 12736 39856 12764
rect 39850 12724 39856 12736
rect 39908 12724 39914 12776
rect 39960 12696 39988 12872
rect 40218 12832 40224 12844
rect 40179 12804 40224 12832
rect 40218 12792 40224 12804
rect 40276 12792 40282 12844
rect 41386 12832 41414 12872
rect 41690 12860 41696 12912
rect 41748 12900 41754 12912
rect 41794 12903 41852 12909
rect 41794 12900 41806 12903
rect 41748 12872 41806 12900
rect 41748 12860 41754 12872
rect 41794 12869 41806 12872
rect 41840 12869 41852 12903
rect 41794 12863 41852 12869
rect 41892 12832 41920 12940
rect 43806 12928 43812 12940
rect 43864 12928 43870 12980
rect 43990 12968 43996 12980
rect 43951 12940 43996 12968
rect 43990 12928 43996 12940
rect 44048 12928 44054 12980
rect 48958 12968 48964 12980
rect 45020 12940 48964 12968
rect 42242 12860 42248 12912
rect 42300 12900 42306 12912
rect 42858 12903 42916 12909
rect 42858 12900 42870 12903
rect 42300 12872 42870 12900
rect 42300 12860 42306 12872
rect 42858 12869 42870 12872
rect 42904 12869 42916 12903
rect 42858 12863 42916 12869
rect 43714 12860 43720 12912
rect 43772 12900 43778 12912
rect 45020 12900 45048 12940
rect 48958 12928 48964 12940
rect 49016 12928 49022 12980
rect 50341 12971 50399 12977
rect 50341 12937 50353 12971
rect 50387 12968 50399 12971
rect 54294 12968 54300 12980
rect 50387 12940 54300 12968
rect 50387 12937 50399 12940
rect 50341 12931 50399 12937
rect 54294 12928 54300 12940
rect 54352 12928 54358 12980
rect 54386 12928 54392 12980
rect 54444 12968 54450 12980
rect 57422 12968 57428 12980
rect 54444 12940 57428 12968
rect 54444 12928 54450 12940
rect 57422 12928 57428 12940
rect 57480 12928 57486 12980
rect 57517 12971 57575 12977
rect 57517 12937 57529 12971
rect 57563 12937 57575 12971
rect 57517 12931 57575 12937
rect 58897 12971 58955 12977
rect 58897 12937 58909 12971
rect 58943 12968 58955 12971
rect 61470 12968 61476 12980
rect 58943 12940 61476 12968
rect 58943 12937 58955 12940
rect 58897 12931 58955 12937
rect 53466 12900 53472 12912
rect 43772 12872 45048 12900
rect 45112 12872 53472 12900
rect 43772 12860 43778 12872
rect 41386 12804 41920 12832
rect 42613 12835 42671 12841
rect 42613 12801 42625 12835
rect 42659 12832 42671 12835
rect 42702 12832 42708 12844
rect 42659 12804 42708 12832
rect 42659 12801 42671 12804
rect 42613 12795 42671 12801
rect 42702 12792 42708 12804
rect 42760 12792 42766 12844
rect 45112 12841 45140 12872
rect 53466 12860 53472 12872
rect 53524 12860 53530 12912
rect 55674 12900 55680 12912
rect 54036 12872 55680 12900
rect 45097 12835 45155 12841
rect 45097 12801 45109 12835
rect 45143 12801 45155 12835
rect 45097 12795 45155 12801
rect 45824 12835 45882 12841
rect 45824 12801 45836 12835
rect 45870 12832 45882 12835
rect 47854 12832 47860 12844
rect 45870 12804 47860 12832
rect 45870 12801 45882 12804
rect 45824 12795 45882 12801
rect 47854 12792 47860 12804
rect 47912 12792 47918 12844
rect 48038 12841 48044 12844
rect 48032 12795 48044 12841
rect 48096 12832 48102 12844
rect 50522 12832 50528 12844
rect 48096 12804 49004 12832
rect 50483 12804 50528 12832
rect 48038 12792 48044 12795
rect 48096 12792 48102 12804
rect 42061 12767 42119 12773
rect 42061 12733 42073 12767
rect 42107 12733 42119 12767
rect 42061 12727 42119 12733
rect 38672 12668 39988 12696
rect 40037 12699 40095 12705
rect 40037 12665 40049 12699
rect 40083 12696 40095 12699
rect 40083 12668 40816 12696
rect 40083 12665 40095 12668
rect 40037 12659 40095 12665
rect 40681 12631 40739 12637
rect 40681 12628 40693 12631
rect 38488 12600 40693 12628
rect 40681 12597 40693 12600
rect 40727 12597 40739 12631
rect 40788 12628 40816 12668
rect 41782 12628 41788 12640
rect 40788 12600 41788 12628
rect 40681 12591 40739 12597
rect 41782 12588 41788 12600
rect 41840 12588 41846 12640
rect 42076 12628 42104 12727
rect 44266 12724 44272 12776
rect 44324 12764 44330 12776
rect 45554 12764 45560 12776
rect 44324 12736 45560 12764
rect 44324 12724 44330 12736
rect 45554 12724 45560 12736
rect 45612 12724 45618 12776
rect 47210 12724 47216 12776
rect 47268 12764 47274 12776
rect 47765 12767 47823 12773
rect 47765 12764 47777 12767
rect 47268 12736 47777 12764
rect 47268 12724 47274 12736
rect 47765 12733 47777 12736
rect 47811 12733 47823 12767
rect 48976 12764 49004 12804
rect 50522 12792 50528 12804
rect 50580 12792 50586 12844
rect 51166 12792 51172 12844
rect 51224 12832 51230 12844
rect 52098 12835 52156 12841
rect 52098 12832 52110 12835
rect 51224 12804 52110 12832
rect 51224 12792 51230 12804
rect 52098 12801 52110 12804
rect 52144 12832 52156 12835
rect 53190 12832 53196 12844
rect 52144 12804 53196 12832
rect 52144 12801 52156 12804
rect 52098 12795 52156 12801
rect 53190 12792 53196 12804
rect 53248 12792 53254 12844
rect 53561 12835 53619 12841
rect 53561 12801 53573 12835
rect 53607 12801 53619 12835
rect 53561 12795 53619 12801
rect 50798 12764 50804 12776
rect 48976 12736 50804 12764
rect 47765 12727 47823 12733
rect 50798 12724 50804 12736
rect 50856 12724 50862 12776
rect 52362 12764 52368 12776
rect 52323 12736 52368 12764
rect 52362 12724 52368 12736
rect 52420 12724 52426 12776
rect 53576 12764 53604 12795
rect 53650 12792 53656 12844
rect 53708 12832 53714 12844
rect 54036 12841 54064 12872
rect 55674 12860 55680 12872
rect 55732 12860 55738 12912
rect 56962 12900 56968 12912
rect 55968 12872 56968 12900
rect 54021 12835 54079 12841
rect 54021 12832 54033 12835
rect 53708 12804 54033 12832
rect 53708 12792 53714 12804
rect 54021 12801 54033 12804
rect 54067 12801 54079 12835
rect 54021 12795 54079 12801
rect 54110 12792 54116 12844
rect 54168 12792 54174 12844
rect 54288 12835 54346 12841
rect 54288 12801 54300 12835
rect 54334 12832 54346 12835
rect 54754 12832 54760 12844
rect 54334 12804 54760 12832
rect 54334 12801 54346 12804
rect 54288 12795 54346 12801
rect 54754 12792 54760 12804
rect 54812 12792 54818 12844
rect 55968 12832 55996 12872
rect 56962 12860 56968 12872
rect 57020 12860 57026 12912
rect 57532 12900 57560 12931
rect 61470 12928 61476 12940
rect 61528 12928 61534 12980
rect 63862 12968 63868 12980
rect 63823 12940 63868 12968
rect 63862 12928 63868 12940
rect 63920 12928 63926 12980
rect 64601 12971 64659 12977
rect 64601 12937 64613 12971
rect 64647 12937 64659 12971
rect 65426 12968 65432 12980
rect 65387 12940 65432 12968
rect 64601 12931 64659 12937
rect 57532 12872 60964 12900
rect 55048 12804 55996 12832
rect 54128 12764 54156 12792
rect 53576 12736 54156 12764
rect 46934 12696 46940 12708
rect 46895 12668 46940 12696
rect 46934 12656 46940 12668
rect 46992 12656 46998 12708
rect 49602 12696 49608 12708
rect 48700 12668 49608 12696
rect 42886 12628 42892 12640
rect 42076 12600 42892 12628
rect 42886 12588 42892 12600
rect 42944 12588 42950 12640
rect 44913 12631 44971 12637
rect 44913 12597 44925 12631
rect 44959 12628 44971 12631
rect 48700 12628 48728 12668
rect 49602 12656 49608 12668
rect 49660 12656 49666 12708
rect 53006 12656 53012 12708
rect 53064 12696 53070 12708
rect 54018 12696 54024 12708
rect 53064 12668 54024 12696
rect 53064 12656 53070 12668
rect 54018 12656 54024 12668
rect 54076 12656 54082 12708
rect 49142 12628 49148 12640
rect 44959 12600 48728 12628
rect 49103 12600 49148 12628
rect 44959 12597 44971 12600
rect 44913 12591 44971 12597
rect 49142 12588 49148 12600
rect 49200 12588 49206 12640
rect 49789 12631 49847 12637
rect 49789 12597 49801 12631
rect 49835 12628 49847 12631
rect 50890 12628 50896 12640
rect 49835 12600 50896 12628
rect 49835 12597 49847 12600
rect 49789 12591 49847 12597
rect 50890 12588 50896 12600
rect 50948 12588 50954 12640
rect 50985 12631 51043 12637
rect 50985 12597 50997 12631
rect 51031 12628 51043 12631
rect 51626 12628 51632 12640
rect 51031 12600 51632 12628
rect 51031 12597 51043 12600
rect 50985 12591 51043 12597
rect 51626 12588 51632 12600
rect 51684 12588 51690 12640
rect 53377 12631 53435 12637
rect 53377 12597 53389 12631
rect 53423 12628 53435 12631
rect 54294 12628 54300 12640
rect 53423 12600 54300 12628
rect 53423 12597 53435 12600
rect 53377 12591 53435 12597
rect 54294 12588 54300 12600
rect 54352 12588 54358 12640
rect 54386 12588 54392 12640
rect 54444 12628 54450 12640
rect 55048 12628 55076 12804
rect 56042 12792 56048 12844
rect 56100 12832 56106 12844
rect 56393 12835 56451 12841
rect 56393 12832 56405 12835
rect 56100 12804 56405 12832
rect 56100 12792 56106 12804
rect 56393 12801 56405 12804
rect 56439 12801 56451 12835
rect 56393 12795 56451 12801
rect 56870 12792 56876 12844
rect 56928 12832 56934 12844
rect 58250 12832 58256 12844
rect 56928 12804 57974 12832
rect 58211 12804 58256 12832
rect 56928 12792 56934 12804
rect 55674 12724 55680 12776
rect 55732 12764 55738 12776
rect 56137 12767 56195 12773
rect 56137 12764 56149 12767
rect 55732 12736 56149 12764
rect 55732 12724 55738 12736
rect 56137 12733 56149 12736
rect 56183 12733 56195 12767
rect 57946 12764 57974 12804
rect 58250 12792 58256 12804
rect 58308 12792 58314 12844
rect 58713 12835 58771 12841
rect 58713 12801 58725 12835
rect 58759 12801 58771 12835
rect 58713 12795 58771 12801
rect 58728 12764 58756 12795
rect 60550 12792 60556 12844
rect 60608 12841 60614 12844
rect 60608 12832 60620 12841
rect 60826 12832 60832 12844
rect 60608 12804 60653 12832
rect 60787 12804 60832 12832
rect 60608 12795 60620 12804
rect 60608 12792 60614 12795
rect 60826 12792 60832 12804
rect 60884 12792 60890 12844
rect 60936 12832 60964 12872
rect 63402 12860 63408 12912
rect 63460 12900 63466 12912
rect 64616 12900 64644 12931
rect 65426 12928 65432 12940
rect 65484 12928 65490 12980
rect 66070 12968 66076 12980
rect 66031 12940 66076 12968
rect 66070 12928 66076 12940
rect 66128 12928 66134 12980
rect 66990 12968 66996 12980
rect 66951 12940 66996 12968
rect 66990 12928 66996 12940
rect 67048 12928 67054 12980
rect 67542 12928 67548 12980
rect 67600 12968 67606 12980
rect 67637 12971 67695 12977
rect 67637 12968 67649 12971
rect 67600 12940 67649 12968
rect 67600 12928 67606 12940
rect 67637 12937 67649 12940
rect 67683 12937 67695 12971
rect 67637 12931 67695 12937
rect 68373 12971 68431 12977
rect 68373 12937 68385 12971
rect 68419 12937 68431 12971
rect 71774 12968 71780 12980
rect 68373 12931 68431 12937
rect 68480 12940 71780 12968
rect 65150 12900 65156 12912
rect 63460 12872 64644 12900
rect 64800 12872 65156 12900
rect 63460 12860 63466 12872
rect 61378 12832 61384 12844
rect 60936 12804 61384 12832
rect 61378 12792 61384 12804
rect 61436 12792 61442 12844
rect 61556 12835 61614 12841
rect 61556 12801 61568 12835
rect 61602 12832 61614 12835
rect 63313 12835 63371 12841
rect 61602 12804 63172 12832
rect 61602 12801 61614 12804
rect 61556 12795 61614 12801
rect 57946 12736 58756 12764
rect 56137 12727 56195 12733
rect 58802 12724 58808 12776
rect 58860 12764 58866 12776
rect 59170 12764 59176 12776
rect 58860 12736 59176 12764
rect 58860 12724 58866 12736
rect 59170 12724 59176 12736
rect 59228 12764 59234 12776
rect 59538 12764 59544 12776
rect 59228 12736 59544 12764
rect 59228 12724 59234 12736
rect 59538 12724 59544 12736
rect 59596 12724 59602 12776
rect 61010 12724 61016 12776
rect 61068 12764 61074 12776
rect 61289 12767 61347 12773
rect 61289 12764 61301 12767
rect 61068 12736 61301 12764
rect 61068 12724 61074 12736
rect 61289 12733 61301 12736
rect 61335 12733 61347 12767
rect 61289 12727 61347 12733
rect 57440 12668 59584 12696
rect 54444 12600 55076 12628
rect 55401 12631 55459 12637
rect 54444 12588 54450 12600
rect 55401 12597 55413 12631
rect 55447 12628 55459 12631
rect 57440 12628 57468 12668
rect 55447 12600 57468 12628
rect 55447 12597 55459 12600
rect 55401 12591 55459 12597
rect 57974 12588 57980 12640
rect 58032 12628 58038 12640
rect 58069 12631 58127 12637
rect 58069 12628 58081 12631
rect 58032 12600 58081 12628
rect 58032 12588 58038 12600
rect 58069 12597 58081 12600
rect 58115 12597 58127 12631
rect 58069 12591 58127 12597
rect 58158 12588 58164 12640
rect 58216 12628 58222 12640
rect 59449 12631 59507 12637
rect 59449 12628 59461 12631
rect 58216 12600 59461 12628
rect 58216 12588 58222 12600
rect 59449 12597 59461 12600
rect 59495 12597 59507 12631
rect 59556 12628 59584 12668
rect 61930 12628 61936 12640
rect 59556 12600 61936 12628
rect 59449 12591 59507 12597
rect 61930 12588 61936 12600
rect 61988 12588 61994 12640
rect 62669 12631 62727 12637
rect 62669 12597 62681 12631
rect 62715 12628 62727 12631
rect 62758 12628 62764 12640
rect 62715 12600 62764 12628
rect 62715 12597 62727 12600
rect 62669 12591 62727 12597
rect 62758 12588 62764 12600
rect 62816 12588 62822 12640
rect 63144 12628 63172 12804
rect 63313 12801 63325 12835
rect 63359 12832 63371 12835
rect 64049 12835 64107 12841
rect 63359 12804 64000 12832
rect 63359 12801 63371 12804
rect 63313 12795 63371 12801
rect 63972 12764 64000 12804
rect 64049 12801 64061 12835
rect 64095 12832 64107 12835
rect 64414 12832 64420 12844
rect 64095 12804 64420 12832
rect 64095 12801 64107 12804
rect 64049 12795 64107 12801
rect 64414 12792 64420 12804
rect 64472 12792 64478 12844
rect 64800 12841 64828 12872
rect 65150 12860 65156 12872
rect 65208 12900 65214 12912
rect 66898 12900 66904 12912
rect 65208 12872 66904 12900
rect 65208 12860 65214 12872
rect 66898 12860 66904 12872
rect 66956 12860 66962 12912
rect 64785 12835 64843 12841
rect 64785 12801 64797 12835
rect 64831 12801 64843 12835
rect 64785 12795 64843 12801
rect 65245 12835 65303 12841
rect 65245 12801 65257 12835
rect 65291 12801 65303 12835
rect 66254 12832 66260 12844
rect 66215 12804 66260 12832
rect 65245 12795 65303 12801
rect 64800 12764 64828 12795
rect 63972 12736 64828 12764
rect 64046 12656 64052 12708
rect 64104 12696 64110 12708
rect 65260 12696 65288 12795
rect 66254 12792 66260 12804
rect 66312 12792 66318 12844
rect 66806 12832 66812 12844
rect 66767 12804 66812 12832
rect 66806 12792 66812 12804
rect 66864 12792 66870 12844
rect 67821 12835 67879 12841
rect 67821 12801 67833 12835
rect 67867 12832 67879 12835
rect 68388 12832 68416 12931
rect 67867 12804 68416 12832
rect 67867 12801 67879 12804
rect 67821 12795 67879 12801
rect 66898 12724 66904 12776
rect 66956 12764 66962 12776
rect 68480 12764 68508 12940
rect 71774 12928 71780 12940
rect 71832 12928 71838 12980
rect 72237 12971 72295 12977
rect 72237 12937 72249 12971
rect 72283 12937 72295 12971
rect 72237 12931 72295 12937
rect 72252 12900 72280 12931
rect 72510 12928 72516 12980
rect 72568 12968 72574 12980
rect 72789 12971 72847 12977
rect 72789 12968 72801 12971
rect 72568 12940 72801 12968
rect 72568 12928 72574 12940
rect 72789 12937 72801 12940
rect 72835 12937 72847 12971
rect 72789 12931 72847 12937
rect 73614 12928 73620 12980
rect 73672 12968 73678 12980
rect 74629 12971 74687 12977
rect 74629 12968 74641 12971
rect 73672 12940 74641 12968
rect 73672 12928 73678 12940
rect 74629 12937 74641 12940
rect 74675 12937 74687 12971
rect 74629 12931 74687 12937
rect 75270 12928 75276 12980
rect 75328 12968 75334 12980
rect 75549 12971 75607 12977
rect 75549 12968 75561 12971
rect 75328 12940 75561 12968
rect 75328 12928 75334 12940
rect 75549 12937 75561 12940
rect 75595 12937 75607 12971
rect 75549 12931 75607 12937
rect 76374 12928 76380 12980
rect 76432 12968 76438 12980
rect 76561 12971 76619 12977
rect 76561 12968 76573 12971
rect 76432 12940 76573 12968
rect 76432 12928 76438 12940
rect 76561 12937 76573 12940
rect 76607 12937 76619 12971
rect 76561 12931 76619 12937
rect 76650 12928 76656 12980
rect 76708 12968 76714 12980
rect 77202 12968 77208 12980
rect 76708 12940 77208 12968
rect 76708 12928 76714 12940
rect 77202 12928 77208 12940
rect 77260 12968 77266 12980
rect 77386 12968 77392 12980
rect 77260 12940 77392 12968
rect 77260 12928 77266 12940
rect 77386 12928 77392 12940
rect 77444 12928 77450 12980
rect 77665 12971 77723 12977
rect 77665 12937 77677 12971
rect 77711 12968 77723 12971
rect 77754 12968 77760 12980
rect 77711 12940 77760 12968
rect 77711 12937 77723 12940
rect 77665 12931 77723 12937
rect 77754 12928 77760 12940
rect 77812 12928 77818 12980
rect 78766 12968 78772 12980
rect 78727 12940 78772 12968
rect 78766 12928 78772 12940
rect 78824 12928 78830 12980
rect 79502 12968 79508 12980
rect 79415 12940 79508 12968
rect 79502 12928 79508 12940
rect 79560 12968 79566 12980
rect 80238 12968 80244 12980
rect 79560 12940 80244 12968
rect 79560 12928 79566 12940
rect 80238 12928 80244 12940
rect 80296 12928 80302 12980
rect 81084 12940 81296 12968
rect 77570 12900 77576 12912
rect 72252 12872 77576 12900
rect 77570 12860 77576 12872
rect 77628 12860 77634 12912
rect 81084 12900 81112 12940
rect 77864 12872 81112 12900
rect 81268 12900 81296 12940
rect 82446 12928 82452 12980
rect 82504 12968 82510 12980
rect 83001 12971 83059 12977
rect 83001 12968 83013 12971
rect 82504 12940 83013 12968
rect 82504 12928 82510 12940
rect 83001 12937 83013 12940
rect 83047 12937 83059 12971
rect 83001 12931 83059 12937
rect 83550 12928 83556 12980
rect 83608 12968 83614 12980
rect 83921 12971 83979 12977
rect 83921 12968 83933 12971
rect 83608 12940 83933 12968
rect 83608 12928 83614 12940
rect 83921 12937 83933 12940
rect 83967 12937 83979 12971
rect 83921 12931 83979 12937
rect 84010 12928 84016 12980
rect 84068 12968 84074 12980
rect 84565 12971 84623 12977
rect 84565 12968 84577 12971
rect 84068 12940 84577 12968
rect 84068 12928 84074 12940
rect 84565 12937 84577 12940
rect 84611 12937 84623 12971
rect 84565 12931 84623 12937
rect 86586 12928 86592 12980
rect 86644 12968 86650 12980
rect 88061 12971 88119 12977
rect 88061 12968 88073 12971
rect 86644 12940 88073 12968
rect 86644 12928 86650 12940
rect 88061 12937 88073 12940
rect 88107 12937 88119 12971
rect 88061 12931 88119 12937
rect 89073 12971 89131 12977
rect 89073 12937 89085 12971
rect 89119 12937 89131 12971
rect 89073 12931 89131 12937
rect 89180 12940 90680 12968
rect 87322 12900 87328 12912
rect 81268 12872 87328 12900
rect 69474 12832 69480 12844
rect 69532 12841 69538 12844
rect 69444 12804 69480 12832
rect 69474 12792 69480 12804
rect 69532 12795 69544 12841
rect 71124 12835 71182 12841
rect 71124 12801 71136 12835
rect 71170 12832 71182 12835
rect 72326 12832 72332 12844
rect 71170 12804 72332 12832
rect 71170 12801 71182 12804
rect 71124 12795 71182 12801
rect 69532 12792 69538 12795
rect 72326 12792 72332 12804
rect 72384 12792 72390 12844
rect 72973 12835 73031 12841
rect 72973 12801 72985 12835
rect 73019 12801 73031 12835
rect 72973 12795 73031 12801
rect 66956 12736 68508 12764
rect 69753 12767 69811 12773
rect 66956 12724 66962 12736
rect 69753 12733 69765 12767
rect 69799 12764 69811 12767
rect 69934 12764 69940 12776
rect 69799 12736 69940 12764
rect 69799 12733 69811 12736
rect 69753 12727 69811 12733
rect 69934 12724 69940 12736
rect 69992 12764 69998 12776
rect 70305 12767 70363 12773
rect 70305 12764 70317 12767
rect 69992 12736 70317 12764
rect 69992 12724 69998 12736
rect 70305 12733 70317 12736
rect 70351 12764 70363 12767
rect 70857 12767 70915 12773
rect 70857 12764 70869 12767
rect 70351 12736 70869 12764
rect 70351 12733 70363 12736
rect 70305 12727 70363 12733
rect 70857 12733 70869 12736
rect 70903 12733 70915 12767
rect 72988 12764 73016 12795
rect 73062 12792 73068 12844
rect 73120 12832 73126 12844
rect 74077 12835 74135 12841
rect 74077 12832 74089 12835
rect 73120 12804 74089 12832
rect 73120 12792 73126 12804
rect 74077 12801 74089 12804
rect 74123 12832 74135 12835
rect 74626 12832 74632 12844
rect 74123 12804 74632 12832
rect 74123 12801 74135 12804
rect 74077 12795 74135 12801
rect 74626 12792 74632 12804
rect 74684 12792 74690 12844
rect 74810 12832 74816 12844
rect 74771 12804 74816 12832
rect 74810 12792 74816 12804
rect 74868 12792 74874 12844
rect 75365 12835 75423 12841
rect 75365 12801 75377 12835
rect 75411 12801 75423 12835
rect 75365 12795 75423 12801
rect 76745 12835 76803 12841
rect 76745 12801 76757 12835
rect 76791 12801 76803 12835
rect 76745 12795 76803 12801
rect 74166 12764 74172 12776
rect 72988 12736 74172 12764
rect 70857 12727 70915 12733
rect 74166 12724 74172 12736
rect 74224 12724 74230 12776
rect 74994 12724 75000 12776
rect 75052 12764 75058 12776
rect 75386 12764 75414 12795
rect 76650 12764 76656 12776
rect 75052 12736 75414 12764
rect 75472 12736 76656 12764
rect 75052 12724 75058 12736
rect 64104 12668 65288 12696
rect 64104 12656 64110 12668
rect 66438 12656 66444 12708
rect 66496 12696 66502 12708
rect 73338 12696 73344 12708
rect 66496 12668 68324 12696
rect 66496 12656 66502 12668
rect 67634 12628 67640 12640
rect 63144 12600 67640 12628
rect 67634 12588 67640 12600
rect 67692 12588 67698 12640
rect 68296 12628 68324 12668
rect 71884 12668 73344 12696
rect 71884 12628 71912 12668
rect 73338 12656 73344 12668
rect 73396 12656 73402 12708
rect 74626 12656 74632 12708
rect 74684 12696 74690 12708
rect 75472 12696 75500 12736
rect 76650 12724 76656 12736
rect 76708 12724 76714 12776
rect 76753 12764 76781 12795
rect 76834 12792 76840 12844
rect 76892 12832 76898 12844
rect 77386 12832 77392 12844
rect 76892 12804 77392 12832
rect 76892 12792 76898 12804
rect 77386 12792 77392 12804
rect 77444 12792 77450 12844
rect 77864 12841 77892 12872
rect 87322 12860 87328 12872
rect 87380 12860 87386 12912
rect 87414 12860 87420 12912
rect 87472 12900 87478 12912
rect 89088 12900 89116 12931
rect 87472 12872 89116 12900
rect 87472 12860 87478 12872
rect 77849 12835 77907 12841
rect 77496 12822 77616 12832
rect 77496 12804 77800 12822
rect 77294 12764 77300 12776
rect 76753 12736 77300 12764
rect 77294 12724 77300 12736
rect 77352 12724 77358 12776
rect 74684 12668 75500 12696
rect 74684 12656 74690 12668
rect 75730 12656 75736 12708
rect 75788 12696 75794 12708
rect 77496 12696 77524 12804
rect 77588 12794 77800 12804
rect 77849 12801 77861 12835
rect 77895 12801 77907 12835
rect 78950 12832 78956 12844
rect 78911 12804 78956 12832
rect 77849 12795 77907 12801
rect 77772 12764 77800 12794
rect 78950 12792 78956 12804
rect 79008 12792 79014 12844
rect 81342 12841 81348 12844
rect 81336 12832 81348 12841
rect 81303 12804 81348 12832
rect 81336 12795 81348 12804
rect 81342 12792 81348 12795
rect 81400 12792 81406 12844
rect 83182 12832 83188 12844
rect 83143 12804 83188 12832
rect 83182 12792 83188 12804
rect 83240 12792 83246 12844
rect 84102 12832 84108 12844
rect 84063 12804 84108 12832
rect 84102 12792 84108 12804
rect 84160 12792 84166 12844
rect 84470 12792 84476 12844
rect 84528 12832 84534 12844
rect 85301 12835 85359 12841
rect 85301 12832 85313 12835
rect 84528 12804 85313 12832
rect 84528 12792 84534 12804
rect 85301 12801 85313 12804
rect 85347 12832 85359 12835
rect 87150 12835 87208 12841
rect 87150 12832 87162 12835
rect 85347 12804 87162 12832
rect 85347 12801 85359 12804
rect 85301 12795 85359 12801
rect 87150 12801 87162 12804
rect 87196 12801 87208 12835
rect 87874 12832 87880 12844
rect 87835 12804 87880 12832
rect 87150 12795 87208 12801
rect 87874 12792 87880 12804
rect 87932 12792 87938 12844
rect 88150 12792 88156 12844
rect 88208 12832 88214 12844
rect 89180 12832 89208 12940
rect 89438 12860 89444 12912
rect 89496 12900 89502 12912
rect 90652 12900 90680 12940
rect 92382 12928 92388 12980
rect 92440 12968 92446 12980
rect 94225 12971 94283 12977
rect 94225 12968 94237 12971
rect 92440 12940 94237 12968
rect 92440 12928 92446 12940
rect 94225 12937 94237 12940
rect 94271 12937 94283 12971
rect 94225 12931 94283 12937
rect 94314 12928 94320 12980
rect 94372 12968 94378 12980
rect 96798 12968 96804 12980
rect 94372 12940 96804 12968
rect 94372 12928 94378 12940
rect 96798 12928 96804 12940
rect 96856 12928 96862 12980
rect 97353 12971 97411 12977
rect 97353 12937 97365 12971
rect 97399 12937 97411 12971
rect 97353 12931 97411 12937
rect 91646 12900 91652 12912
rect 89496 12872 90588 12900
rect 89496 12860 89502 12872
rect 88208 12804 89208 12832
rect 89257 12835 89315 12841
rect 88208 12792 88214 12804
rect 89257 12801 89269 12835
rect 89303 12801 89315 12835
rect 89257 12795 89315 12801
rect 81069 12767 81127 12773
rect 81069 12764 81081 12767
rect 77772 12736 80376 12764
rect 75788 12668 77524 12696
rect 75788 12656 75794 12668
rect 68296 12600 71912 12628
rect 73893 12631 73951 12637
rect 73893 12597 73905 12631
rect 73939 12628 73951 12631
rect 74258 12628 74264 12640
rect 73939 12600 74264 12628
rect 73939 12597 73951 12600
rect 73893 12591 73951 12597
rect 74258 12588 74264 12600
rect 74316 12588 74322 12640
rect 75638 12588 75644 12640
rect 75696 12628 75702 12640
rect 77478 12628 77484 12640
rect 75696 12600 77484 12628
rect 75696 12588 75702 12600
rect 77478 12588 77484 12600
rect 77536 12588 77542 12640
rect 80057 12631 80115 12637
rect 80057 12597 80069 12631
rect 80103 12628 80115 12631
rect 80238 12628 80244 12640
rect 80103 12600 80244 12628
rect 80103 12597 80115 12600
rect 80057 12591 80115 12597
rect 80238 12588 80244 12600
rect 80296 12588 80302 12640
rect 80348 12628 80376 12736
rect 80532 12736 81081 12764
rect 80532 12708 80560 12736
rect 81069 12733 81081 12736
rect 81115 12733 81127 12767
rect 81069 12727 81127 12733
rect 82078 12724 82084 12776
rect 82136 12764 82142 12776
rect 85390 12764 85396 12776
rect 82136 12736 85396 12764
rect 82136 12724 82142 12736
rect 85390 12724 85396 12736
rect 85448 12724 85454 12776
rect 85482 12724 85488 12776
rect 85540 12764 85546 12776
rect 87417 12767 87475 12773
rect 85540 12736 85585 12764
rect 85540 12724 85546 12736
rect 87417 12733 87429 12767
rect 87463 12764 87475 12767
rect 88426 12764 88432 12776
rect 87463 12736 88432 12764
rect 87463 12733 87475 12736
rect 87417 12727 87475 12733
rect 80514 12696 80520 12708
rect 80475 12668 80520 12696
rect 80514 12656 80520 12668
rect 80572 12656 80578 12708
rect 86037 12699 86095 12705
rect 86037 12696 86049 12699
rect 82004 12668 86049 12696
rect 82004 12628 82032 12668
rect 86037 12665 86049 12668
rect 86083 12665 86095 12699
rect 86037 12659 86095 12665
rect 82446 12628 82452 12640
rect 80348 12600 82032 12628
rect 82407 12600 82452 12628
rect 82446 12588 82452 12600
rect 82504 12588 82510 12640
rect 84654 12588 84660 12640
rect 84712 12628 84718 12640
rect 85117 12631 85175 12637
rect 85117 12628 85129 12631
rect 84712 12600 85129 12628
rect 84712 12588 84718 12600
rect 85117 12597 85129 12600
rect 85163 12597 85175 12631
rect 85117 12591 85175 12597
rect 86770 12588 86776 12640
rect 86828 12628 86834 12640
rect 87432 12628 87460 12727
rect 88426 12724 88432 12736
rect 88484 12724 88490 12776
rect 89272 12764 89300 12795
rect 89346 12792 89352 12844
rect 89404 12832 89410 12844
rect 89717 12835 89775 12841
rect 89717 12832 89729 12835
rect 89404 12804 89729 12832
rect 89404 12792 89410 12804
rect 89717 12801 89729 12804
rect 89763 12801 89775 12835
rect 89717 12795 89775 12801
rect 89806 12764 89812 12776
rect 89272 12736 89812 12764
rect 89806 12724 89812 12736
rect 89864 12724 89870 12776
rect 90453 12767 90511 12773
rect 90453 12733 90465 12767
rect 90499 12733 90511 12767
rect 90560 12764 90588 12872
rect 90652 12872 91652 12900
rect 90652 12841 90680 12872
rect 91646 12860 91652 12872
rect 91704 12860 91710 12912
rect 95326 12900 95332 12912
rect 94424 12872 95332 12900
rect 90637 12835 90695 12841
rect 90637 12801 90649 12835
rect 90683 12801 90695 12835
rect 90637 12795 90695 12801
rect 91281 12835 91339 12841
rect 91281 12801 91293 12835
rect 91327 12832 91339 12835
rect 91370 12832 91376 12844
rect 91327 12804 91376 12832
rect 91327 12801 91339 12804
rect 91281 12795 91339 12801
rect 91296 12764 91324 12795
rect 91370 12792 91376 12804
rect 91428 12792 91434 12844
rect 91548 12835 91606 12841
rect 91548 12801 91560 12835
rect 91594 12832 91606 12835
rect 91594 12804 93348 12832
rect 91594 12801 91606 12804
rect 91548 12795 91606 12801
rect 90560 12736 91324 12764
rect 93320 12764 93348 12804
rect 93394 12792 93400 12844
rect 93452 12832 93458 12844
rect 94424 12841 94452 12872
rect 95326 12860 95332 12872
rect 95384 12860 95390 12912
rect 95970 12860 95976 12912
rect 96028 12900 96034 12912
rect 97368 12900 97396 12931
rect 97626 12928 97632 12980
rect 97684 12968 97690 12980
rect 98181 12971 98239 12977
rect 98181 12968 98193 12971
rect 97684 12940 98193 12968
rect 97684 12928 97690 12940
rect 98181 12937 98193 12940
rect 98227 12937 98239 12971
rect 98181 12931 98239 12937
rect 98546 12928 98552 12980
rect 98604 12968 98610 12980
rect 100018 12968 100024 12980
rect 98604 12940 100024 12968
rect 98604 12928 98610 12940
rect 100018 12928 100024 12940
rect 100076 12928 100082 12980
rect 100110 12928 100116 12980
rect 100168 12968 100174 12980
rect 100941 12971 100999 12977
rect 100941 12968 100953 12971
rect 100168 12940 100953 12968
rect 100168 12928 100174 12940
rect 100941 12937 100953 12940
rect 100987 12937 100999 12971
rect 100941 12931 100999 12937
rect 101766 12928 101772 12980
rect 101824 12968 101830 12980
rect 102413 12971 102471 12977
rect 102413 12968 102425 12971
rect 101824 12940 102425 12968
rect 101824 12928 101830 12940
rect 102413 12937 102425 12940
rect 102459 12937 102471 12971
rect 102413 12931 102471 12937
rect 102594 12928 102600 12980
rect 102652 12968 102658 12980
rect 103149 12971 103207 12977
rect 103149 12968 103161 12971
rect 102652 12940 103161 12968
rect 102652 12928 102658 12940
rect 103149 12937 103161 12940
rect 103195 12937 103207 12971
rect 103149 12931 103207 12937
rect 103974 12928 103980 12980
rect 104032 12968 104038 12980
rect 104529 12971 104587 12977
rect 104529 12968 104541 12971
rect 104032 12940 104541 12968
rect 104032 12928 104038 12940
rect 104529 12937 104541 12940
rect 104575 12937 104587 12971
rect 104529 12931 104587 12937
rect 104802 12928 104808 12980
rect 104860 12968 104866 12980
rect 107010 12968 107016 12980
rect 104860 12940 107016 12968
rect 104860 12928 104866 12940
rect 107010 12928 107016 12940
rect 107068 12928 107074 12980
rect 107286 12928 107292 12980
rect 107344 12968 107350 12980
rect 108301 12971 108359 12977
rect 108301 12968 108313 12971
rect 107344 12940 108313 12968
rect 107344 12928 107350 12940
rect 108301 12937 108313 12940
rect 108347 12937 108359 12971
rect 108301 12931 108359 12937
rect 108390 12928 108396 12980
rect 108448 12968 108454 12980
rect 109681 12971 109739 12977
rect 109681 12968 109693 12971
rect 108448 12940 109693 12968
rect 108448 12928 108454 12940
rect 109681 12937 109693 12940
rect 109727 12937 109739 12971
rect 109681 12931 109739 12937
rect 112254 12928 112260 12980
rect 112312 12968 112318 12980
rect 112901 12971 112959 12977
rect 112901 12968 112913 12971
rect 112312 12940 112913 12968
rect 112312 12928 112318 12940
rect 112901 12937 112913 12940
rect 112947 12937 112959 12971
rect 113634 12968 113640 12980
rect 113595 12940 113640 12968
rect 112901 12931 112959 12937
rect 113634 12928 113640 12940
rect 113692 12928 113698 12980
rect 117682 12968 117688 12980
rect 113744 12940 117688 12968
rect 98454 12900 98460 12912
rect 96028 12872 97396 12900
rect 97460 12872 98460 12900
rect 96028 12860 96034 12872
rect 94409 12835 94467 12841
rect 93452 12804 93497 12832
rect 93452 12792 93458 12804
rect 94409 12801 94421 12835
rect 94455 12801 94467 12835
rect 94409 12795 94467 12801
rect 95421 12835 95479 12841
rect 95421 12801 95433 12835
rect 95467 12832 95479 12835
rect 95510 12832 95516 12844
rect 95467 12804 95516 12832
rect 95467 12801 95479 12804
rect 95421 12795 95479 12801
rect 95510 12792 95516 12804
rect 95568 12792 95574 12844
rect 95688 12835 95746 12841
rect 95688 12801 95700 12835
rect 95734 12832 95746 12835
rect 97460 12832 97488 12872
rect 98454 12860 98460 12872
rect 98512 12860 98518 12912
rect 100386 12900 100392 12912
rect 99484 12872 100392 12900
rect 95734 12804 97488 12832
rect 97537 12835 97595 12841
rect 95734 12801 95746 12804
rect 95688 12795 95746 12801
rect 97537 12801 97549 12835
rect 97583 12801 97595 12835
rect 97994 12832 98000 12844
rect 97955 12804 98000 12832
rect 97537 12795 97595 12801
rect 94222 12764 94228 12776
rect 93320 12736 94228 12764
rect 90453 12727 90511 12733
rect 87966 12656 87972 12708
rect 88024 12696 88030 12708
rect 89901 12699 89959 12705
rect 89901 12696 89913 12699
rect 88024 12668 89913 12696
rect 88024 12656 88030 12668
rect 89901 12665 89913 12668
rect 89947 12665 89959 12699
rect 90468 12696 90496 12727
rect 94222 12724 94228 12736
rect 94280 12724 94286 12776
rect 95234 12764 95240 12776
rect 94608 12736 95240 12764
rect 90542 12696 90548 12708
rect 90468 12668 90548 12696
rect 89901 12659 89959 12665
rect 90542 12656 90548 12668
rect 90600 12656 90606 12708
rect 92661 12699 92719 12705
rect 92661 12665 92673 12699
rect 92707 12696 92719 12699
rect 94314 12696 94320 12708
rect 92707 12668 94320 12696
rect 92707 12665 92719 12668
rect 92661 12659 92719 12665
rect 94314 12656 94320 12668
rect 94372 12656 94378 12708
rect 86828 12600 87460 12628
rect 86828 12588 86834 12600
rect 88886 12588 88892 12640
rect 88944 12628 88950 12640
rect 89530 12628 89536 12640
rect 88944 12600 89536 12628
rect 88944 12588 88950 12600
rect 89530 12588 89536 12600
rect 89588 12588 89594 12640
rect 90821 12631 90879 12637
rect 90821 12597 90833 12631
rect 90867 12628 90879 12631
rect 92382 12628 92388 12640
rect 90867 12600 92388 12628
rect 90867 12597 90879 12600
rect 90821 12591 90879 12597
rect 92382 12588 92388 12600
rect 92440 12588 92446 12640
rect 93210 12628 93216 12640
rect 93171 12600 93216 12628
rect 93210 12588 93216 12600
rect 93268 12588 93274 12640
rect 93394 12588 93400 12640
rect 93452 12628 93458 12640
rect 94608 12628 94636 12736
rect 95234 12724 95240 12736
rect 95292 12724 95298 12776
rect 97552 12764 97580 12795
rect 97994 12792 98000 12804
rect 98052 12792 98058 12844
rect 99484 12841 99512 12872
rect 100386 12860 100392 12872
rect 100444 12860 100450 12912
rect 103882 12900 103888 12912
rect 101876 12872 103888 12900
rect 99469 12835 99527 12841
rect 99469 12801 99481 12835
rect 99515 12801 99527 12835
rect 100110 12832 100116 12844
rect 100071 12804 100116 12832
rect 99469 12795 99527 12801
rect 100110 12792 100116 12804
rect 100168 12792 100174 12844
rect 101125 12835 101183 12841
rect 101125 12801 101137 12835
rect 101171 12832 101183 12835
rect 101306 12832 101312 12844
rect 101171 12804 101312 12832
rect 101171 12801 101183 12804
rect 101125 12795 101183 12801
rect 101306 12792 101312 12804
rect 101364 12792 101370 12844
rect 101876 12841 101904 12872
rect 103882 12860 103888 12872
rect 103940 12860 103946 12912
rect 104066 12860 104072 12912
rect 104124 12900 104130 12912
rect 106768 12903 106826 12909
rect 104124 12872 106274 12900
rect 104124 12860 104130 12872
rect 101861 12835 101919 12841
rect 101861 12801 101873 12835
rect 101907 12801 101919 12835
rect 101861 12795 101919 12801
rect 102597 12835 102655 12841
rect 102597 12801 102609 12835
rect 102643 12801 102655 12835
rect 102597 12795 102655 12801
rect 103333 12835 103391 12841
rect 103333 12801 103345 12835
rect 103379 12832 103391 12835
rect 104713 12835 104771 12841
rect 103379 12804 104664 12832
rect 103379 12801 103391 12804
rect 103333 12795 103391 12801
rect 99374 12764 99380 12776
rect 97552 12736 99380 12764
rect 99374 12724 99380 12736
rect 99432 12724 99438 12776
rect 99653 12767 99711 12773
rect 99653 12733 99665 12767
rect 99699 12764 99711 12767
rect 100202 12764 100208 12776
rect 99699 12736 100208 12764
rect 99699 12733 99711 12736
rect 99653 12727 99711 12733
rect 100202 12724 100208 12736
rect 100260 12724 100266 12776
rect 102612 12764 102640 12795
rect 103606 12764 103612 12776
rect 102612 12736 103612 12764
rect 103606 12724 103612 12736
rect 103664 12724 103670 12776
rect 103882 12764 103888 12776
rect 103843 12736 103888 12764
rect 103882 12724 103888 12736
rect 103940 12724 103946 12776
rect 104636 12764 104664 12804
rect 104713 12801 104725 12835
rect 104759 12832 104771 12835
rect 104894 12832 104900 12844
rect 104759 12804 104900 12832
rect 104759 12801 104771 12804
rect 104713 12795 104771 12801
rect 104894 12792 104900 12804
rect 104952 12792 104958 12844
rect 106246 12832 106274 12872
rect 106768 12869 106780 12903
rect 106814 12900 106826 12903
rect 109402 12900 109408 12912
rect 106814 12872 109408 12900
rect 106814 12869 106826 12872
rect 106768 12863 106826 12869
rect 109402 12860 109408 12872
rect 109460 12860 109466 12912
rect 112104 12903 112162 12909
rect 112104 12869 112116 12903
rect 112150 12900 112162 12903
rect 113266 12900 113272 12912
rect 112150 12872 113272 12900
rect 112150 12869 112162 12872
rect 112104 12863 112162 12869
rect 113266 12860 113272 12872
rect 113324 12860 113330 12912
rect 106918 12832 106924 12844
rect 106246 12804 106924 12832
rect 106918 12792 106924 12804
rect 106976 12792 106982 12844
rect 107749 12835 107807 12841
rect 107749 12801 107761 12835
rect 107795 12832 107807 12835
rect 108114 12832 108120 12844
rect 107795 12804 108120 12832
rect 107795 12801 107807 12804
rect 107749 12795 107807 12801
rect 108114 12792 108120 12804
rect 108172 12792 108178 12844
rect 108485 12835 108543 12841
rect 108485 12801 108497 12835
rect 108531 12801 108543 12835
rect 108485 12795 108543 12801
rect 105722 12764 105728 12776
rect 104636 12736 105728 12764
rect 105722 12724 105728 12736
rect 105780 12724 105786 12776
rect 107010 12764 107016 12776
rect 106971 12736 107016 12764
rect 107010 12724 107016 12736
rect 107068 12724 107074 12776
rect 108500 12764 108528 12795
rect 109034 12792 109040 12844
rect 109092 12832 109098 12844
rect 109865 12835 109923 12841
rect 109092 12804 109137 12832
rect 109092 12792 109098 12804
rect 109865 12801 109877 12835
rect 109911 12832 109923 12835
rect 113085 12835 113143 12841
rect 109911 12804 113036 12832
rect 109911 12801 109923 12804
rect 109865 12795 109923 12801
rect 112349 12767 112407 12773
rect 108500 12736 109457 12764
rect 94682 12656 94688 12708
rect 94740 12696 94746 12708
rect 96801 12699 96859 12705
rect 94740 12668 95004 12696
rect 94740 12656 94746 12668
rect 94866 12628 94872 12640
rect 93452 12600 94636 12628
rect 94827 12600 94872 12628
rect 93452 12588 93458 12600
rect 94866 12588 94872 12600
rect 94924 12588 94930 12640
rect 94976 12628 95004 12668
rect 96801 12665 96813 12699
rect 96847 12696 96859 12699
rect 96890 12696 96896 12708
rect 96847 12668 96896 12696
rect 96847 12665 96859 12668
rect 96801 12659 96859 12665
rect 96890 12656 96896 12668
rect 96948 12656 96954 12708
rect 96982 12656 96988 12708
rect 97040 12696 97046 12708
rect 97040 12668 99512 12696
rect 97040 12656 97046 12668
rect 97994 12628 98000 12640
rect 94976 12600 98000 12628
rect 97994 12588 98000 12600
rect 98052 12588 98058 12640
rect 99282 12628 99288 12640
rect 99243 12600 99288 12628
rect 99282 12588 99288 12600
rect 99340 12588 99346 12640
rect 99484 12628 99512 12668
rect 99558 12656 99564 12708
rect 99616 12696 99622 12708
rect 100297 12699 100355 12705
rect 100297 12696 100309 12699
rect 99616 12668 100309 12696
rect 99616 12656 99622 12668
rect 100297 12665 100309 12668
rect 100343 12665 100355 12699
rect 100297 12659 100355 12665
rect 100662 12656 100668 12708
rect 100720 12696 100726 12708
rect 101677 12699 101735 12705
rect 101677 12696 101689 12699
rect 100720 12668 101689 12696
rect 100720 12656 100726 12668
rect 101677 12665 101689 12668
rect 101723 12665 101735 12699
rect 105633 12699 105691 12705
rect 105633 12696 105645 12699
rect 101677 12659 101735 12665
rect 101784 12668 105645 12696
rect 101784 12628 101812 12668
rect 105633 12665 105645 12668
rect 105679 12665 105691 12699
rect 107028 12696 107056 12724
rect 108942 12696 108948 12708
rect 107028 12668 108948 12696
rect 105633 12659 105691 12665
rect 108942 12656 108948 12668
rect 109000 12656 109006 12708
rect 109429 12696 109457 12736
rect 112349 12733 112361 12767
rect 112395 12764 112407 12767
rect 112438 12764 112444 12776
rect 112395 12736 112444 12764
rect 112395 12733 112407 12736
rect 112349 12727 112407 12733
rect 112438 12724 112444 12736
rect 112496 12724 112502 12776
rect 113008 12764 113036 12804
rect 113085 12801 113097 12835
rect 113131 12832 113143 12835
rect 113744 12832 113772 12940
rect 117682 12928 117688 12940
rect 117740 12928 117746 12980
rect 117774 12928 117780 12980
rect 117832 12968 117838 12980
rect 118513 12971 118571 12977
rect 118513 12968 118525 12971
rect 117832 12940 118525 12968
rect 117832 12928 117838 12940
rect 118513 12937 118525 12940
rect 118559 12937 118571 12971
rect 118513 12931 118571 12937
rect 119706 12928 119712 12980
rect 119764 12968 119770 12980
rect 119985 12971 120043 12977
rect 119985 12968 119997 12971
rect 119764 12940 119997 12968
rect 119764 12928 119770 12940
rect 119985 12937 119997 12940
rect 120031 12937 120043 12971
rect 119985 12931 120043 12937
rect 120074 12928 120080 12980
rect 120132 12968 120138 12980
rect 120721 12971 120779 12977
rect 120721 12968 120733 12971
rect 120132 12940 120733 12968
rect 120132 12928 120138 12940
rect 120721 12937 120733 12940
rect 120767 12937 120779 12971
rect 120721 12931 120779 12937
rect 121086 12928 121092 12980
rect 121144 12968 121150 12980
rect 121457 12971 121515 12977
rect 121457 12968 121469 12971
rect 121144 12940 121469 12968
rect 121144 12928 121150 12940
rect 121457 12937 121469 12940
rect 121503 12937 121515 12971
rect 123202 12968 123208 12980
rect 121457 12931 121515 12937
rect 121564 12940 123208 12968
rect 115008 12903 115066 12909
rect 115008 12869 115020 12903
rect 115054 12900 115066 12903
rect 120626 12900 120632 12912
rect 115054 12872 120632 12900
rect 115054 12869 115066 12872
rect 115008 12863 115066 12869
rect 120626 12860 120632 12872
rect 120684 12860 120690 12912
rect 113131 12804 113772 12832
rect 113821 12835 113879 12841
rect 113131 12801 113143 12804
rect 113085 12795 113143 12801
rect 113821 12801 113833 12835
rect 113867 12832 113879 12835
rect 115750 12832 115756 12844
rect 113867 12804 115756 12832
rect 113867 12801 113879 12804
rect 113821 12795 113879 12801
rect 115750 12792 115756 12804
rect 115808 12792 115814 12844
rect 115842 12792 115848 12844
rect 115900 12832 115906 12844
rect 116578 12832 116584 12844
rect 115900 12804 116584 12832
rect 115900 12792 115906 12804
rect 116578 12792 116584 12804
rect 116636 12792 116642 12844
rect 116848 12835 116906 12841
rect 116848 12801 116860 12835
rect 116894 12832 116906 12835
rect 118697 12835 118755 12841
rect 116894 12804 118648 12832
rect 116894 12801 116906 12804
rect 116848 12795 116906 12801
rect 113542 12764 113548 12776
rect 113008 12736 113548 12764
rect 113542 12724 113548 12736
rect 113600 12724 113606 12776
rect 114738 12764 114744 12776
rect 114699 12736 114744 12764
rect 114738 12724 114744 12736
rect 114796 12724 114802 12776
rect 110322 12696 110328 12708
rect 109429 12668 110328 12696
rect 110322 12656 110328 12668
rect 110380 12656 110386 12708
rect 114462 12656 114468 12708
rect 114520 12696 114526 12708
rect 117958 12696 117964 12708
rect 114520 12668 114784 12696
rect 114520 12656 114526 12668
rect 99484 12600 101812 12628
rect 103790 12588 103796 12640
rect 103848 12628 103854 12640
rect 104802 12628 104808 12640
rect 103848 12600 104808 12628
rect 103848 12588 103854 12600
rect 104802 12588 104808 12600
rect 104860 12588 104866 12640
rect 106274 12588 106280 12640
rect 106332 12628 106338 12640
rect 107565 12631 107623 12637
rect 107565 12628 107577 12631
rect 106332 12600 107577 12628
rect 106332 12588 106338 12600
rect 107565 12597 107577 12600
rect 107611 12597 107623 12631
rect 107565 12591 107623 12597
rect 107654 12588 107660 12640
rect 107712 12628 107718 12640
rect 109126 12628 109132 12640
rect 107712 12600 109132 12628
rect 107712 12588 107718 12600
rect 109126 12588 109132 12600
rect 109184 12588 109190 12640
rect 109402 12588 109408 12640
rect 109460 12628 109466 12640
rect 110414 12628 110420 12640
rect 109460 12600 110420 12628
rect 109460 12588 109466 12600
rect 110414 12588 110420 12600
rect 110472 12588 110478 12640
rect 110966 12628 110972 12640
rect 110927 12600 110972 12628
rect 110966 12588 110972 12600
rect 111024 12588 111030 12640
rect 111334 12588 111340 12640
rect 111392 12628 111398 12640
rect 114554 12628 114560 12640
rect 111392 12600 114560 12628
rect 111392 12588 111398 12600
rect 114554 12588 114560 12600
rect 114612 12588 114618 12640
rect 114756 12628 114784 12668
rect 115952 12668 116624 12696
rect 117919 12668 117964 12696
rect 115952 12628 115980 12668
rect 116118 12628 116124 12640
rect 114756 12600 115980 12628
rect 116079 12600 116124 12628
rect 116118 12588 116124 12600
rect 116176 12588 116182 12640
rect 116596 12628 116624 12668
rect 117958 12656 117964 12668
rect 118016 12656 118022 12708
rect 118620 12696 118648 12804
rect 118697 12801 118709 12835
rect 118743 12801 118755 12835
rect 118697 12795 118755 12801
rect 118712 12764 118740 12795
rect 118786 12792 118792 12844
rect 118844 12832 118850 12844
rect 119246 12832 119252 12844
rect 118844 12804 119252 12832
rect 118844 12792 118850 12804
rect 119246 12792 119252 12804
rect 119304 12792 119310 12844
rect 120166 12832 120172 12844
rect 120127 12804 120172 12832
rect 120166 12792 120172 12804
rect 120224 12792 120230 12844
rect 120905 12835 120963 12841
rect 120905 12801 120917 12835
rect 120951 12832 120963 12835
rect 121454 12832 121460 12844
rect 120951 12804 121460 12832
rect 120951 12801 120963 12804
rect 120905 12795 120963 12801
rect 121454 12792 121460 12804
rect 121512 12792 121518 12844
rect 121564 12764 121592 12940
rect 123202 12928 123208 12940
rect 123260 12928 123266 12980
rect 123294 12928 123300 12980
rect 123352 12968 123358 12980
rect 125137 12971 125195 12977
rect 125137 12968 125149 12971
rect 123352 12940 125149 12968
rect 123352 12928 123358 12940
rect 125137 12937 125149 12940
rect 125183 12937 125195 12971
rect 125137 12931 125195 12937
rect 125318 12928 125324 12980
rect 125376 12968 125382 12980
rect 126882 12968 126888 12980
rect 125376 12940 126888 12968
rect 125376 12928 125382 12940
rect 126882 12928 126888 12940
rect 126940 12928 126946 12980
rect 128262 12928 128268 12980
rect 128320 12968 128326 12980
rect 128817 12971 128875 12977
rect 128817 12968 128829 12971
rect 128320 12940 128829 12968
rect 128320 12928 128326 12940
rect 128817 12937 128829 12940
rect 128863 12937 128875 12971
rect 129550 12968 129556 12980
rect 129511 12940 129556 12968
rect 128817 12931 128875 12937
rect 129550 12928 129556 12940
rect 129608 12928 129614 12980
rect 129734 12928 129740 12980
rect 129792 12968 129798 12980
rect 130289 12971 130347 12977
rect 130289 12968 130301 12971
rect 129792 12940 130301 12968
rect 129792 12928 129798 12940
rect 130289 12937 130301 12940
rect 130335 12937 130347 12971
rect 130289 12931 130347 12937
rect 130470 12928 130476 12980
rect 130528 12968 130534 12980
rect 131025 12971 131083 12977
rect 131025 12968 131037 12971
rect 130528 12940 131037 12968
rect 130528 12928 130534 12940
rect 131025 12937 131037 12940
rect 131071 12937 131083 12971
rect 131206 12968 131212 12980
rect 131025 12931 131083 12937
rect 131132 12940 131212 12968
rect 123386 12900 123392 12912
rect 121656 12872 123392 12900
rect 121656 12841 121684 12872
rect 123386 12860 123392 12872
rect 123444 12860 123450 12912
rect 125962 12900 125968 12912
rect 124140 12872 125968 12900
rect 121641 12835 121699 12841
rect 121641 12801 121653 12835
rect 121687 12801 121699 12835
rect 121641 12795 121699 12801
rect 122460 12835 122518 12841
rect 122460 12801 122472 12835
rect 122506 12832 122518 12835
rect 124140 12832 124168 12872
rect 125962 12860 125968 12872
rect 126020 12860 126026 12912
rect 126974 12900 126980 12912
rect 126072 12872 126980 12900
rect 124306 12832 124312 12844
rect 122506 12804 124168 12832
rect 124267 12804 124312 12832
rect 122506 12801 122518 12804
rect 122460 12795 122518 12801
rect 124306 12792 124312 12804
rect 124364 12792 124370 12844
rect 126072 12841 126100 12872
rect 126974 12860 126980 12872
rect 127032 12860 127038 12912
rect 127152 12903 127210 12909
rect 127152 12869 127164 12903
rect 127198 12900 127210 12903
rect 127342 12900 127348 12912
rect 127198 12872 127348 12900
rect 127198 12869 127210 12872
rect 127152 12863 127210 12869
rect 127342 12860 127348 12872
rect 127400 12860 127406 12912
rect 127434 12860 127440 12912
rect 127492 12900 127498 12912
rect 130010 12900 130016 12912
rect 127492 12872 130016 12900
rect 127492 12860 127498 12872
rect 130010 12860 130016 12872
rect 130068 12860 130074 12912
rect 131132 12900 131160 12940
rect 131206 12928 131212 12940
rect 131264 12928 131270 12980
rect 131850 12968 131856 12980
rect 131811 12940 131856 12968
rect 131850 12928 131856 12940
rect 131908 12928 131914 12980
rect 131942 12928 131948 12980
rect 132000 12968 132006 12980
rect 133598 12968 133604 12980
rect 132000 12940 133604 12968
rect 132000 12928 132006 12940
rect 133598 12928 133604 12940
rect 133656 12928 133662 12980
rect 133782 12928 133788 12980
rect 133840 12968 133846 12980
rect 134153 12971 134211 12977
rect 134153 12968 134165 12971
rect 133840 12940 134165 12968
rect 133840 12928 133846 12940
rect 134153 12937 134165 12940
rect 134199 12937 134211 12971
rect 134153 12931 134211 12937
rect 134886 12928 134892 12980
rect 134944 12968 134950 12980
rect 135533 12971 135591 12977
rect 135533 12968 135545 12971
rect 134944 12940 135545 12968
rect 134944 12928 134950 12940
rect 135533 12937 135545 12940
rect 135579 12937 135591 12971
rect 135533 12931 135591 12937
rect 136542 12928 136548 12980
rect 136600 12968 136606 12980
rect 136821 12971 136879 12977
rect 136821 12968 136833 12971
rect 136600 12940 136833 12968
rect 136600 12928 136606 12940
rect 136821 12937 136833 12940
rect 136867 12937 136879 12971
rect 137922 12968 137928 12980
rect 137883 12940 137928 12968
rect 136821 12931 136879 12937
rect 137922 12928 137928 12940
rect 137980 12928 137986 12980
rect 139486 12928 139492 12980
rect 139544 12968 139550 12980
rect 139581 12971 139639 12977
rect 139581 12968 139593 12971
rect 139544 12940 139593 12968
rect 139544 12928 139550 12940
rect 139581 12937 139593 12940
rect 139627 12937 139639 12971
rect 139581 12931 139639 12937
rect 140590 12928 140596 12980
rect 140648 12968 140654 12980
rect 140869 12971 140927 12977
rect 140869 12968 140881 12971
rect 140648 12940 140881 12968
rect 140648 12928 140654 12940
rect 140869 12937 140881 12940
rect 140915 12937 140927 12971
rect 140869 12931 140927 12937
rect 142154 12928 142160 12980
rect 142212 12968 142218 12980
rect 142893 12971 142951 12977
rect 142893 12968 142905 12971
rect 142212 12940 142905 12968
rect 142212 12928 142218 12940
rect 142893 12937 142905 12940
rect 142939 12937 142951 12971
rect 146294 12968 146300 12980
rect 142893 12931 142951 12937
rect 143276 12940 146300 12968
rect 130120 12872 131160 12900
rect 131224 12872 133092 12900
rect 125321 12835 125379 12841
rect 125321 12801 125333 12835
rect 125367 12801 125379 12835
rect 125321 12795 125379 12801
rect 126057 12835 126115 12841
rect 126057 12801 126069 12835
rect 126103 12801 126115 12835
rect 128814 12832 128820 12844
rect 126057 12795 126115 12801
rect 126808 12804 128820 12832
rect 118712 12736 121592 12764
rect 122006 12724 122012 12776
rect 122064 12764 122070 12776
rect 122193 12767 122251 12773
rect 122193 12764 122205 12767
rect 122064 12736 122205 12764
rect 122064 12724 122070 12736
rect 122193 12733 122205 12736
rect 122239 12733 122251 12767
rect 125336 12764 125364 12795
rect 126808 12764 126836 12804
rect 128814 12792 128820 12804
rect 128872 12792 128878 12844
rect 128998 12832 129004 12844
rect 128959 12804 129004 12832
rect 128998 12792 129004 12804
rect 129056 12792 129062 12844
rect 129918 12832 129924 12844
rect 129200 12804 129924 12832
rect 125336 12736 126836 12764
rect 122193 12727 122251 12733
rect 126882 12724 126888 12776
rect 126940 12764 126946 12776
rect 126940 12736 126985 12764
rect 126940 12724 126946 12736
rect 127986 12724 127992 12776
rect 128044 12764 128050 12776
rect 129200 12764 129228 12804
rect 129918 12792 129924 12804
rect 129976 12792 129982 12844
rect 130120 12764 130148 12872
rect 130470 12832 130476 12844
rect 130431 12804 130476 12832
rect 130470 12792 130476 12804
rect 130528 12792 130534 12844
rect 131224 12841 131252 12872
rect 131209 12835 131267 12841
rect 131209 12801 131221 12835
rect 131255 12801 131267 12835
rect 131209 12795 131267 12801
rect 131669 12835 131727 12841
rect 131669 12801 131681 12835
rect 131715 12801 131727 12835
rect 133064 12832 133092 12872
rect 133138 12860 133144 12912
rect 133196 12900 133202 12912
rect 138566 12900 138572 12912
rect 133196 12872 138572 12900
rect 133196 12860 133202 12872
rect 138566 12860 138572 12872
rect 138624 12860 138630 12912
rect 143276 12900 143304 12940
rect 146294 12928 146300 12940
rect 146352 12928 146358 12980
rect 149425 12971 149483 12977
rect 149425 12968 149437 12971
rect 149256 12940 149437 12968
rect 138952 12872 143304 12900
rect 134150 12832 134156 12844
rect 133064 12804 134156 12832
rect 131669 12795 131727 12801
rect 128044 12736 129228 12764
rect 129752 12736 130148 12764
rect 128044 12724 128050 12736
rect 120166 12696 120172 12708
rect 118620 12668 120172 12696
rect 120166 12656 120172 12668
rect 120224 12656 120230 12708
rect 123573 12699 123631 12705
rect 123573 12665 123585 12699
rect 123619 12696 123631 12699
rect 129752 12696 129780 12736
rect 130562 12724 130568 12776
rect 130620 12764 130626 12776
rect 131684 12764 131712 12795
rect 134150 12792 134156 12804
rect 134208 12792 134214 12844
rect 134334 12832 134340 12844
rect 134295 12804 134340 12832
rect 134334 12792 134340 12804
rect 134392 12792 134398 12844
rect 135374 12835 135432 12841
rect 135374 12832 135386 12835
rect 135370 12801 135386 12832
rect 135420 12801 135432 12835
rect 136634 12832 136640 12844
rect 136595 12804 136640 12832
rect 135370 12795 135432 12801
rect 132770 12764 132776 12776
rect 130620 12736 131712 12764
rect 132731 12736 132776 12764
rect 130620 12724 130626 12736
rect 132770 12724 132776 12736
rect 132828 12724 132834 12776
rect 133046 12764 133052 12776
rect 133007 12736 133052 12764
rect 133046 12724 133052 12736
rect 133104 12724 133110 12776
rect 135370 12696 135398 12795
rect 136634 12792 136640 12804
rect 136692 12792 136698 12844
rect 137738 12832 137744 12844
rect 137699 12804 137744 12832
rect 137738 12792 137744 12804
rect 137796 12792 137802 12844
rect 138952 12841 138980 12872
rect 143350 12860 143356 12912
rect 143408 12900 143414 12912
rect 146788 12903 146846 12909
rect 143408 12872 145144 12900
rect 143408 12860 143414 12872
rect 138937 12835 138995 12841
rect 138937 12801 138949 12835
rect 138983 12801 138995 12835
rect 138937 12795 138995 12801
rect 139397 12835 139455 12841
rect 139397 12801 139409 12835
rect 139443 12801 139455 12835
rect 139397 12795 139455 12801
rect 135714 12724 135720 12776
rect 135772 12764 135778 12776
rect 136085 12767 136143 12773
rect 136085 12764 136097 12767
rect 135772 12736 136097 12764
rect 135772 12724 135778 12736
rect 136085 12733 136097 12736
rect 136131 12733 136143 12767
rect 136085 12727 136143 12733
rect 136174 12724 136180 12776
rect 136232 12764 136238 12776
rect 139412 12764 139440 12795
rect 139578 12792 139584 12844
rect 139636 12832 139642 12844
rect 141510 12832 141516 12844
rect 139636 12804 141516 12832
rect 139636 12792 139642 12804
rect 141510 12792 141516 12804
rect 141568 12792 141574 12844
rect 141993 12835 142051 12841
rect 141993 12801 142005 12835
rect 142039 12832 142051 12835
rect 142522 12832 142528 12844
rect 142039 12804 142528 12832
rect 142039 12801 142051 12804
rect 141993 12795 142051 12801
rect 142522 12792 142528 12804
rect 142580 12792 142586 12844
rect 142706 12832 142712 12844
rect 142667 12804 142712 12832
rect 142706 12792 142712 12804
rect 142764 12792 142770 12844
rect 145116 12841 145144 12872
rect 146788 12869 146800 12903
rect 146834 12900 146846 12903
rect 148502 12900 148508 12912
rect 146834 12872 148508 12900
rect 146834 12869 146846 12872
rect 146788 12863 146846 12869
rect 148502 12860 148508 12872
rect 148560 12860 148566 12912
rect 148778 12860 148784 12912
rect 148836 12900 148842 12912
rect 149256 12900 149284 12940
rect 149425 12937 149437 12940
rect 149471 12937 149483 12971
rect 149425 12931 149483 12937
rect 150894 12928 150900 12980
rect 150952 12968 150958 12980
rect 151998 12968 152004 12980
rect 150952 12940 152004 12968
rect 150952 12928 150958 12940
rect 151998 12928 152004 12940
rect 152056 12928 152062 12980
rect 152918 12928 152924 12980
rect 152976 12968 152982 12980
rect 153470 12968 153476 12980
rect 152976 12940 153476 12968
rect 152976 12928 152982 12940
rect 153470 12928 153476 12940
rect 153528 12928 153534 12980
rect 156138 12968 156144 12980
rect 156099 12940 156144 12968
rect 156138 12928 156144 12940
rect 156196 12928 156202 12980
rect 156782 12928 156788 12980
rect 156840 12968 156846 12980
rect 156877 12971 156935 12977
rect 156877 12968 156889 12971
rect 156840 12940 156889 12968
rect 156840 12928 156846 12940
rect 156877 12937 156889 12940
rect 156923 12937 156935 12971
rect 158070 12968 158076 12980
rect 158031 12940 158076 12968
rect 156877 12931 156935 12937
rect 158070 12928 158076 12940
rect 158128 12928 158134 12980
rect 148836 12872 149284 12900
rect 148836 12860 148842 12872
rect 151354 12860 151360 12912
rect 151412 12900 151418 12912
rect 152458 12900 152464 12912
rect 151412 12872 152464 12900
rect 151412 12860 151418 12872
rect 144845 12835 144903 12841
rect 144845 12801 144857 12835
rect 144891 12832 144903 12835
rect 145101 12835 145159 12841
rect 144891 12804 145052 12832
rect 144891 12801 144903 12804
rect 144845 12795 144903 12801
rect 136232 12736 139440 12764
rect 142249 12767 142307 12773
rect 136232 12724 136238 12736
rect 142249 12733 142261 12767
rect 142295 12764 142307 12767
rect 145024 12764 145052 12804
rect 145101 12801 145113 12835
rect 145147 12801 145159 12835
rect 145101 12795 145159 12801
rect 147033 12835 147091 12841
rect 147033 12801 147045 12835
rect 147079 12832 147091 12835
rect 147490 12832 147496 12844
rect 147079 12804 147496 12832
rect 147079 12801 147091 12804
rect 147033 12795 147091 12801
rect 147490 12792 147496 12804
rect 147548 12792 147554 12844
rect 147760 12835 147818 12841
rect 147760 12801 147772 12835
rect 147806 12832 147818 12835
rect 148870 12832 148876 12844
rect 147806 12804 148876 12832
rect 147806 12801 147818 12804
rect 147760 12795 147818 12801
rect 148870 12792 148876 12804
rect 148928 12792 148934 12844
rect 149514 12792 149520 12844
rect 149572 12832 149578 12844
rect 149609 12835 149667 12841
rect 149609 12832 149621 12835
rect 149572 12804 149621 12832
rect 149572 12792 149578 12804
rect 149609 12801 149621 12804
rect 149655 12801 149667 12835
rect 149609 12795 149667 12801
rect 149698 12792 149704 12844
rect 149756 12832 149762 12844
rect 152200 12841 152228 12872
rect 152458 12860 152464 12872
rect 152516 12900 152522 12912
rect 155402 12900 155408 12912
rect 152516 12872 154068 12900
rect 152516 12860 152522 12872
rect 150253 12835 150311 12841
rect 150253 12832 150265 12835
rect 149756 12804 150265 12832
rect 149756 12792 149762 12804
rect 150253 12801 150265 12804
rect 150299 12801 150311 12835
rect 151918 12835 151976 12841
rect 151918 12832 151930 12835
rect 150253 12795 150311 12801
rect 150360 12804 151930 12832
rect 145834 12764 145840 12776
rect 142295 12736 144132 12764
rect 145024 12736 145840 12764
rect 142295 12733 142307 12736
rect 142249 12727 142307 12733
rect 123619 12668 126928 12696
rect 123619 12665 123631 12668
rect 123573 12659 123631 12665
rect 118142 12628 118148 12640
rect 116596 12600 118148 12628
rect 118142 12588 118148 12600
rect 118200 12588 118206 12640
rect 119154 12628 119160 12640
rect 119115 12600 119160 12628
rect 119154 12588 119160 12600
rect 119212 12588 119218 12640
rect 119246 12588 119252 12640
rect 119304 12628 119310 12640
rect 122374 12628 122380 12640
rect 119304 12600 122380 12628
rect 119304 12588 119310 12600
rect 122374 12588 122380 12600
rect 122432 12588 122438 12640
rect 122466 12588 122472 12640
rect 122524 12628 122530 12640
rect 124125 12631 124183 12637
rect 124125 12628 124137 12631
rect 122524 12600 124137 12628
rect 122524 12588 122530 12600
rect 124125 12597 124137 12600
rect 124171 12597 124183 12631
rect 124125 12591 124183 12597
rect 125226 12588 125232 12640
rect 125284 12628 125290 12640
rect 125873 12631 125931 12637
rect 125873 12628 125885 12631
rect 125284 12600 125885 12628
rect 125284 12588 125290 12600
rect 125873 12597 125885 12600
rect 125919 12597 125931 12631
rect 125873 12591 125931 12597
rect 125962 12588 125968 12640
rect 126020 12628 126026 12640
rect 126698 12628 126704 12640
rect 126020 12600 126704 12628
rect 126020 12588 126026 12600
rect 126698 12588 126704 12600
rect 126756 12588 126762 12640
rect 126900 12628 126928 12668
rect 127820 12668 129780 12696
rect 129844 12668 135398 12696
rect 127820 12628 127848 12668
rect 126900 12600 127848 12628
rect 128265 12631 128323 12637
rect 128265 12597 128277 12631
rect 128311 12628 128323 12631
rect 129844 12628 129872 12668
rect 142338 12656 142344 12708
rect 142396 12696 142402 12708
rect 143721 12699 143779 12705
rect 143721 12696 143733 12699
rect 142396 12668 143733 12696
rect 142396 12656 142402 12668
rect 143721 12665 143733 12668
rect 143767 12696 143779 12699
rect 143902 12696 143908 12708
rect 143767 12668 143908 12696
rect 143767 12665 143779 12668
rect 143721 12659 143779 12665
rect 143902 12656 143908 12668
rect 143960 12656 143966 12708
rect 128311 12600 129872 12628
rect 128311 12597 128323 12600
rect 128265 12591 128323 12597
rect 129918 12588 129924 12640
rect 129976 12628 129982 12640
rect 135346 12628 135352 12640
rect 129976 12600 135352 12628
rect 129976 12588 129982 12600
rect 135346 12588 135352 12600
rect 135404 12588 135410 12640
rect 138753 12631 138811 12637
rect 138753 12597 138765 12631
rect 138799 12628 138811 12631
rect 142614 12628 142620 12640
rect 138799 12600 142620 12628
rect 138799 12597 138811 12600
rect 138753 12591 138811 12597
rect 142614 12588 142620 12600
rect 142672 12588 142678 12640
rect 144104 12628 144132 12736
rect 145834 12724 145840 12736
rect 145892 12724 145898 12776
rect 150360 12764 150388 12804
rect 151918 12801 151930 12804
rect 151964 12801 151976 12835
rect 151918 12795 151976 12801
rect 152185 12835 152243 12841
rect 152185 12801 152197 12835
rect 152231 12801 152243 12835
rect 153378 12832 153384 12844
rect 152185 12795 152243 12801
rect 152292 12804 153384 12832
rect 149348 12736 150388 12764
rect 148873 12699 148931 12705
rect 148873 12665 148885 12699
rect 148919 12696 148931 12699
rect 149146 12696 149152 12708
rect 148919 12668 149152 12696
rect 148919 12665 148931 12668
rect 148873 12659 148931 12665
rect 149146 12656 149152 12668
rect 149204 12656 149210 12708
rect 149348 12696 149376 12736
rect 150066 12696 150072 12708
rect 149256 12668 149376 12696
rect 150027 12668 150072 12696
rect 144730 12628 144736 12640
rect 144104 12600 144736 12628
rect 144730 12588 144736 12600
rect 144788 12588 144794 12640
rect 145558 12588 145564 12640
rect 145616 12628 145622 12640
rect 145653 12631 145711 12637
rect 145653 12628 145665 12631
rect 145616 12600 145665 12628
rect 145616 12588 145622 12600
rect 145653 12597 145665 12600
rect 145699 12597 145711 12631
rect 145653 12591 145711 12597
rect 147030 12588 147036 12640
rect 147088 12628 147094 12640
rect 149256 12628 149284 12668
rect 150066 12656 150072 12668
rect 150124 12656 150130 12708
rect 150802 12696 150808 12708
rect 150763 12668 150808 12696
rect 150802 12656 150808 12668
rect 150860 12656 150866 12708
rect 147088 12600 149284 12628
rect 147088 12588 147094 12600
rect 150342 12588 150348 12640
rect 150400 12628 150406 12640
rect 152292 12628 152320 12804
rect 153378 12792 153384 12804
rect 153436 12792 153442 12844
rect 153746 12792 153752 12844
rect 153804 12841 153810 12844
rect 154040 12841 154068 12872
rect 154592 12872 155408 12900
rect 154592 12841 154620 12872
rect 155402 12860 155408 12872
rect 155460 12860 155466 12912
rect 155586 12860 155592 12912
rect 155644 12900 155650 12912
rect 155644 12872 158300 12900
rect 155644 12860 155650 12872
rect 153804 12832 153816 12841
rect 154025 12835 154083 12841
rect 153804 12804 153849 12832
rect 153804 12795 153816 12804
rect 154025 12801 154037 12835
rect 154071 12801 154083 12835
rect 154025 12795 154083 12801
rect 154577 12835 154635 12841
rect 154577 12801 154589 12835
rect 154623 12801 154635 12835
rect 154577 12795 154635 12801
rect 154669 12835 154727 12841
rect 154669 12801 154681 12835
rect 154715 12801 154727 12835
rect 154669 12795 154727 12801
rect 155957 12835 156015 12841
rect 155957 12801 155969 12835
rect 156003 12832 156015 12835
rect 156046 12832 156052 12844
rect 156003 12804 156052 12832
rect 156003 12801 156015 12804
rect 155957 12795 156015 12801
rect 153804 12792 153810 12795
rect 154114 12724 154120 12776
rect 154172 12764 154178 12776
rect 154684 12764 154712 12795
rect 156046 12792 156052 12804
rect 156104 12792 156110 12844
rect 156690 12832 156696 12844
rect 156651 12804 156696 12832
rect 156690 12792 156696 12804
rect 156748 12792 156754 12844
rect 158272 12841 158300 12872
rect 157613 12835 157671 12841
rect 157613 12801 157625 12835
rect 157659 12801 157671 12835
rect 157613 12795 157671 12801
rect 158257 12835 158315 12841
rect 158257 12801 158269 12835
rect 158303 12801 158315 12835
rect 158257 12795 158315 12801
rect 154172 12736 154712 12764
rect 154853 12767 154911 12773
rect 154172 12724 154178 12736
rect 154853 12733 154865 12767
rect 154899 12764 154911 12767
rect 157628 12764 157656 12795
rect 158346 12764 158352 12776
rect 154899 12736 157564 12764
rect 157628 12736 158352 12764
rect 154899 12733 154911 12736
rect 154853 12727 154911 12733
rect 152642 12696 152648 12708
rect 152603 12668 152648 12696
rect 152642 12656 152648 12668
rect 152700 12656 152706 12708
rect 155313 12699 155371 12705
rect 155313 12696 155325 12699
rect 154040 12668 155325 12696
rect 150400 12600 152320 12628
rect 150400 12588 150406 12600
rect 152734 12588 152740 12640
rect 152792 12628 152798 12640
rect 154040 12628 154068 12668
rect 155313 12665 155325 12668
rect 155359 12665 155371 12699
rect 157429 12699 157487 12705
rect 157429 12696 157441 12699
rect 155313 12659 155371 12665
rect 155972 12668 157441 12696
rect 152792 12600 154068 12628
rect 152792 12588 152798 12600
rect 154298 12588 154304 12640
rect 154356 12628 154362 12640
rect 155972 12628 156000 12668
rect 157429 12665 157441 12668
rect 157475 12665 157487 12699
rect 157536 12696 157564 12736
rect 158346 12724 158352 12736
rect 158404 12724 158410 12776
rect 158162 12696 158168 12708
rect 157536 12668 158168 12696
rect 157429 12659 157487 12665
rect 158162 12656 158168 12668
rect 158220 12656 158226 12708
rect 154356 12600 156000 12628
rect 154356 12588 154362 12600
rect 1104 12538 158884 12560
rect 1104 12486 20672 12538
rect 20724 12486 20736 12538
rect 20788 12486 20800 12538
rect 20852 12486 20864 12538
rect 20916 12486 20928 12538
rect 20980 12486 60117 12538
rect 60169 12486 60181 12538
rect 60233 12486 60245 12538
rect 60297 12486 60309 12538
rect 60361 12486 60373 12538
rect 60425 12486 99562 12538
rect 99614 12486 99626 12538
rect 99678 12486 99690 12538
rect 99742 12486 99754 12538
rect 99806 12486 99818 12538
rect 99870 12486 139007 12538
rect 139059 12486 139071 12538
rect 139123 12486 139135 12538
rect 139187 12486 139199 12538
rect 139251 12486 139263 12538
rect 139315 12486 158884 12538
rect 1104 12464 158884 12486
rect 10502 12424 10508 12436
rect 10463 12396 10508 12424
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 12066 12424 12072 12436
rect 11072 12396 12072 12424
rect 7745 12359 7803 12365
rect 7745 12325 7757 12359
rect 7791 12356 7803 12359
rect 11072 12356 11100 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13998 12424 14004 12436
rect 13679 12396 14004 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14148 12396 21680 12424
rect 14148 12384 14154 12396
rect 7791 12328 11100 12356
rect 12084 12328 13032 12356
rect 7791 12325 7803 12328
rect 7745 12319 7803 12325
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10962 12288 10968 12300
rect 10100 12260 10968 12288
rect 10100 12248 10106 12260
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 4430 12180 4436 12232
rect 4488 12220 4494 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4488 12192 4629 12220
rect 4488 12180 4494 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 5776 12192 6377 12220
rect 5776 12180 5782 12192
rect 6365 12189 6377 12192
rect 6411 12220 6423 12223
rect 9858 12220 9864 12232
rect 6411 12192 9352 12220
rect 9819 12192 9864 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6632 12155 6690 12161
rect 6632 12121 6644 12155
rect 6678 12152 6690 12155
rect 6822 12152 6828 12164
rect 6678 12124 6828 12152
rect 6678 12121 6690 12124
rect 6632 12115 6690 12121
rect 6822 12112 6828 12124
rect 6880 12112 6886 12164
rect 9324 12161 9352 12192
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11054 12220 11060 12232
rect 10967 12192 11060 12220
rect 11054 12180 11060 12192
rect 11112 12220 11118 12232
rect 12084 12220 12112 12328
rect 11112 12192 12112 12220
rect 11112 12180 11118 12192
rect 9309 12155 9367 12161
rect 9309 12121 9321 12155
rect 9355 12152 9367 12155
rect 11072 12152 11100 12180
rect 9355 12124 11100 12152
rect 11324 12155 11382 12161
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 11324 12121 11336 12155
rect 11370 12152 11382 12155
rect 11698 12152 11704 12164
rect 11370 12124 11704 12152
rect 11370 12121 11382 12124
rect 11324 12115 11382 12121
rect 11698 12112 11704 12124
rect 11756 12112 11762 12164
rect 13004 12161 13032 12328
rect 19886 12316 19892 12368
rect 19944 12356 19950 12368
rect 20622 12356 20628 12368
rect 19944 12328 20628 12356
rect 19944 12316 19950 12328
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 21652 12356 21680 12396
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22152 12396 22197 12424
rect 22152 12384 22158 12396
rect 22830 12384 22836 12436
rect 22888 12424 22894 12436
rect 23017 12427 23075 12433
rect 23017 12424 23029 12427
rect 22888 12396 23029 12424
rect 22888 12384 22894 12396
rect 23017 12393 23029 12396
rect 23063 12393 23075 12427
rect 23017 12387 23075 12393
rect 23845 12427 23903 12433
rect 23845 12393 23857 12427
rect 23891 12424 23903 12427
rect 24486 12424 24492 12436
rect 23891 12396 24492 12424
rect 23891 12393 23903 12396
rect 23845 12387 23903 12393
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 27246 12424 27252 12436
rect 24596 12396 27108 12424
rect 27207 12396 27252 12424
rect 24394 12356 24400 12368
rect 21652 12328 24400 12356
rect 24394 12316 24400 12328
rect 24452 12316 24458 12368
rect 24596 12288 24624 12396
rect 26142 12316 26148 12368
rect 26200 12356 26206 12368
rect 26421 12359 26479 12365
rect 26421 12356 26433 12359
rect 26200 12328 26433 12356
rect 26200 12316 26206 12328
rect 26421 12325 26433 12328
rect 26467 12325 26479 12359
rect 27080 12356 27108 12396
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 27798 12384 27804 12436
rect 27856 12424 27862 12436
rect 27985 12427 28043 12433
rect 27985 12424 27997 12427
rect 27856 12396 27997 12424
rect 27856 12384 27862 12396
rect 27985 12393 27997 12396
rect 28031 12393 28043 12427
rect 27985 12387 28043 12393
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 29917 12427 29975 12433
rect 29917 12424 29929 12427
rect 29512 12396 29929 12424
rect 29512 12384 29518 12396
rect 29917 12393 29929 12396
rect 29963 12393 29975 12427
rect 30650 12424 30656 12436
rect 30611 12396 30656 12424
rect 29917 12387 29975 12393
rect 30650 12384 30656 12396
rect 30708 12384 30714 12436
rect 31294 12424 31300 12436
rect 31128 12396 31300 12424
rect 31128 12356 31156 12396
rect 31294 12384 31300 12396
rect 31352 12384 31358 12436
rect 31662 12384 31668 12436
rect 31720 12424 31726 12436
rect 32677 12427 32735 12433
rect 32677 12424 32689 12427
rect 31720 12396 32689 12424
rect 31720 12384 31726 12396
rect 32677 12393 32689 12396
rect 32723 12393 32735 12427
rect 32677 12387 32735 12393
rect 33870 12384 33876 12436
rect 33928 12424 33934 12436
rect 34057 12427 34115 12433
rect 34057 12424 34069 12427
rect 33928 12396 34069 12424
rect 33928 12384 33934 12396
rect 34057 12393 34069 12396
rect 34103 12393 34115 12427
rect 35158 12424 35164 12436
rect 35119 12396 35164 12424
rect 34057 12387 34115 12393
rect 35158 12384 35164 12396
rect 35216 12384 35222 12436
rect 36078 12384 36084 12436
rect 36136 12424 36142 12436
rect 36357 12427 36415 12433
rect 36357 12424 36369 12427
rect 36136 12396 36369 12424
rect 36136 12384 36142 12396
rect 36357 12393 36369 12396
rect 36403 12393 36415 12427
rect 36357 12387 36415 12393
rect 37182 12384 37188 12436
rect 37240 12424 37246 12436
rect 37369 12427 37427 12433
rect 37369 12424 37381 12427
rect 37240 12396 37381 12424
rect 37240 12384 37246 12396
rect 37369 12393 37381 12396
rect 37415 12393 37427 12427
rect 37369 12387 37427 12393
rect 38286 12384 38292 12436
rect 38344 12424 38350 12436
rect 38565 12427 38623 12433
rect 38565 12424 38577 12427
rect 38344 12396 38577 12424
rect 38344 12384 38350 12396
rect 38565 12393 38577 12396
rect 38611 12393 38623 12427
rect 38565 12387 38623 12393
rect 39393 12427 39451 12433
rect 39393 12393 39405 12427
rect 39439 12424 39451 12427
rect 39942 12424 39948 12436
rect 39439 12396 39948 12424
rect 39439 12393 39451 12396
rect 39393 12387 39451 12393
rect 39942 12384 39948 12396
rect 40000 12384 40006 12436
rect 40052 12396 41414 12424
rect 38102 12356 38108 12368
rect 27080 12328 31156 12356
rect 32232 12328 38108 12356
rect 26421 12319 26479 12325
rect 32030 12288 32036 12300
rect 23216 12260 24624 12288
rect 28184 12260 29868 12288
rect 31991 12260 32036 12288
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13228 12192 13461 12220
rect 13228 12180 13234 12192
rect 13449 12189 13461 12192
rect 13495 12220 13507 12223
rect 13538 12220 13544 12232
rect 13495 12192 13544 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 14826 12220 14832 12232
rect 14787 12192 14832 12220
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 16206 12220 16212 12232
rect 15620 12192 16212 12220
rect 15620 12180 15626 12192
rect 16206 12180 16212 12192
rect 16264 12220 16270 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 16264 12192 17417 12220
rect 16264 12180 16270 12192
rect 17405 12189 17417 12192
rect 17451 12220 17463 12223
rect 19426 12220 19432 12232
rect 17451 12192 19432 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20714 12220 20720 12232
rect 20675 12192 20720 12220
rect 20714 12180 20720 12192
rect 20772 12220 20778 12232
rect 21450 12220 21456 12232
rect 20772 12192 21456 12220
rect 20772 12180 20778 12192
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 23216 12229 23244 12260
rect 28184 12232 28212 12260
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12189 24087 12223
rect 24578 12220 24584 12232
rect 24539 12192 24584 12220
rect 24029 12183 24087 12189
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 13035 12124 14381 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 14369 12121 14381 12124
rect 14415 12152 14427 12155
rect 14458 12152 14464 12164
rect 14415 12124 14464 12152
rect 14415 12121 14427 12124
rect 14369 12115 14427 12121
rect 14458 12112 14464 12124
rect 14516 12152 14522 12164
rect 15580 12152 15608 12180
rect 14516 12124 15608 12152
rect 14516 12112 14522 12124
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15810 12155 15868 12161
rect 15810 12152 15822 12155
rect 15712 12124 15822 12152
rect 15712 12112 15718 12124
rect 15810 12121 15822 12124
rect 15856 12121 15868 12155
rect 15810 12115 15868 12121
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 17650 12155 17708 12161
rect 17650 12152 17662 12155
rect 16356 12124 17662 12152
rect 16356 12112 16362 12124
rect 17650 12121 17662 12124
rect 17696 12121 17708 12155
rect 20165 12155 20223 12161
rect 20165 12152 20177 12155
rect 17650 12115 17708 12121
rect 17880 12124 20177 12152
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4212 12056 4445 12084
rect 4212 12044 4218 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 9582 12084 9588 12096
rect 8619 12056 9588 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 14918 12084 14924 12096
rect 12483 12056 14924 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15013 12087 15071 12093
rect 15013 12053 15025 12087
rect 15059 12084 15071 12087
rect 16114 12084 16120 12096
rect 15059 12056 16120 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17880 12084 17908 12124
rect 20165 12121 20177 12124
rect 20211 12152 20223 12155
rect 20962 12155 21020 12161
rect 20962 12152 20974 12155
rect 20211 12124 20974 12152
rect 20211 12121 20223 12124
rect 20165 12115 20223 12121
rect 20962 12121 20974 12124
rect 21008 12121 21020 12155
rect 24044 12152 24072 12183
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 27338 12220 27344 12232
rect 24780 12192 27344 12220
rect 24780 12152 24808 12192
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12189 27491 12223
rect 28166 12220 28172 12232
rect 28079 12192 28172 12220
rect 27433 12183 27491 12189
rect 24854 12161 24860 12164
rect 24044 12124 24808 12152
rect 20962 12115 21020 12121
rect 24848 12115 24860 12161
rect 24912 12152 24918 12164
rect 26602 12152 26608 12164
rect 24912 12124 24948 12152
rect 25056 12124 26096 12152
rect 26563 12124 26608 12152
rect 24854 12112 24860 12115
rect 24912 12112 24918 12124
rect 17276 12056 17908 12084
rect 18785 12087 18843 12093
rect 17276 12044 17282 12056
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 18874 12084 18880 12096
rect 18831 12056 18880 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19300 12056 19625 12084
rect 19300 12044 19306 12056
rect 19613 12053 19625 12056
rect 19659 12084 19671 12087
rect 20714 12084 20720 12096
rect 19659 12056 20720 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 24118 12044 24124 12096
rect 24176 12084 24182 12096
rect 25056 12084 25084 12124
rect 24176 12056 25084 12084
rect 24176 12044 24182 12056
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 25961 12087 26019 12093
rect 25961 12084 25973 12087
rect 25832 12056 25973 12084
rect 25832 12044 25838 12056
rect 25961 12053 25973 12056
rect 26007 12053 26019 12087
rect 26068 12084 26096 12124
rect 26602 12112 26608 12124
rect 26660 12112 26666 12164
rect 26970 12112 26976 12164
rect 27028 12152 27034 12164
rect 27448 12152 27476 12183
rect 28166 12180 28172 12192
rect 28224 12180 28230 12232
rect 28350 12180 28356 12232
rect 28408 12220 28414 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 28408 12192 29745 12220
rect 28408 12180 28414 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29840 12220 29868 12260
rect 32030 12248 32036 12260
rect 32088 12248 32094 12300
rect 32232 12220 32260 12328
rect 38102 12316 38108 12328
rect 38160 12316 38166 12368
rect 38194 12316 38200 12368
rect 38252 12356 38258 12368
rect 40052 12356 40080 12396
rect 38252 12328 40080 12356
rect 41386 12356 41414 12396
rect 41690 12384 41696 12436
rect 41748 12424 41754 12436
rect 44266 12424 44272 12436
rect 41748 12396 44272 12424
rect 41748 12384 41754 12396
rect 44266 12384 44272 12396
rect 44324 12384 44330 12436
rect 44545 12427 44603 12433
rect 44545 12393 44557 12427
rect 44591 12424 44603 12427
rect 45554 12424 45560 12436
rect 44591 12396 45560 12424
rect 44591 12393 44603 12396
rect 44545 12387 44603 12393
rect 45554 12384 45560 12396
rect 45612 12384 45618 12436
rect 47026 12384 47032 12436
rect 47084 12424 47090 12436
rect 48774 12424 48780 12436
rect 47084 12396 48780 12424
rect 47084 12384 47090 12396
rect 48774 12384 48780 12396
rect 48832 12384 48838 12436
rect 49789 12427 49847 12433
rect 49789 12393 49801 12427
rect 49835 12424 49847 12427
rect 52362 12424 52368 12436
rect 49835 12396 51074 12424
rect 49835 12393 49847 12396
rect 49789 12387 49847 12393
rect 42150 12356 42156 12368
rect 41386 12328 42156 12356
rect 38252 12316 38258 12328
rect 42150 12316 42156 12328
rect 42208 12316 42214 12368
rect 42245 12359 42303 12365
rect 42245 12325 42257 12359
rect 42291 12356 42303 12359
rect 43530 12356 43536 12368
rect 42291 12328 43536 12356
rect 42291 12325 42303 12328
rect 42245 12319 42303 12325
rect 43530 12316 43536 12328
rect 43588 12316 43594 12368
rect 43809 12359 43867 12365
rect 43809 12325 43821 12359
rect 43855 12356 43867 12359
rect 43898 12356 43904 12368
rect 43855 12328 43904 12356
rect 43855 12325 43867 12328
rect 43809 12319 43867 12325
rect 43898 12316 43904 12328
rect 43956 12316 43962 12368
rect 50801 12359 50859 12365
rect 50801 12325 50813 12359
rect 50847 12325 50859 12359
rect 51046 12356 51074 12396
rect 52104 12396 52368 12424
rect 51442 12356 51448 12368
rect 51046 12328 51448 12356
rect 50801 12319 50859 12325
rect 34256 12260 40356 12288
rect 34256 12229 34284 12260
rect 29840 12192 32260 12220
rect 32493 12223 32551 12229
rect 29733 12183 29791 12189
rect 32493 12189 32505 12223
rect 32539 12189 32551 12223
rect 32493 12183 32551 12189
rect 34241 12223 34299 12229
rect 34241 12189 34253 12223
rect 34287 12189 34299 12223
rect 35342 12220 35348 12232
rect 35303 12192 35348 12220
rect 34241 12183 34299 12189
rect 27028 12124 27476 12152
rect 27028 12112 27034 12124
rect 28534 12112 28540 12164
rect 28592 12152 28598 12164
rect 31766 12155 31824 12161
rect 31766 12152 31778 12155
rect 28592 12124 31778 12152
rect 28592 12112 28598 12124
rect 31766 12121 31778 12124
rect 31812 12121 31824 12155
rect 31766 12115 31824 12121
rect 28552 12084 28580 12112
rect 29178 12084 29184 12096
rect 26068 12056 28580 12084
rect 29091 12056 29184 12084
rect 25961 12047 26019 12053
rect 29178 12044 29184 12056
rect 29236 12084 29242 12096
rect 30650 12084 30656 12096
rect 29236 12056 30656 12084
rect 29236 12044 29242 12056
rect 30650 12044 30656 12056
rect 30708 12044 30714 12096
rect 30926 12044 30932 12096
rect 30984 12084 30990 12096
rect 32508 12084 32536 12183
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 36170 12220 36176 12232
rect 36131 12192 36176 12220
rect 36170 12180 36176 12192
rect 36228 12180 36234 12232
rect 36354 12180 36360 12232
rect 36412 12220 36418 12232
rect 37553 12223 37611 12229
rect 37553 12220 37565 12223
rect 36412 12192 37565 12220
rect 36412 12180 36418 12192
rect 37553 12189 37565 12192
rect 37599 12220 37611 12223
rect 38194 12220 38200 12232
rect 37599 12192 38200 12220
rect 37599 12189 37611 12192
rect 37553 12183 37611 12189
rect 38194 12180 38200 12192
rect 38252 12180 38258 12232
rect 38378 12220 38384 12232
rect 38339 12192 38384 12220
rect 38378 12180 38384 12192
rect 38436 12180 38442 12232
rect 39206 12220 39212 12232
rect 39167 12192 39212 12220
rect 39206 12180 39212 12192
rect 39264 12180 39270 12232
rect 40218 12220 40224 12232
rect 40179 12192 40224 12220
rect 40218 12180 40224 12192
rect 40276 12180 40282 12232
rect 40328 12220 40356 12260
rect 41230 12248 41236 12300
rect 41288 12288 41294 12300
rect 42705 12291 42763 12297
rect 42705 12288 42717 12291
rect 41288 12260 42717 12288
rect 41288 12248 41294 12260
rect 42705 12257 42717 12260
rect 42751 12257 42763 12291
rect 43990 12288 43996 12300
rect 42705 12251 42763 12257
rect 43548 12260 43996 12288
rect 41414 12220 41420 12232
rect 40328 12192 41420 12220
rect 41414 12180 41420 12192
rect 41472 12180 41478 12232
rect 42058 12220 42064 12232
rect 42019 12192 42064 12220
rect 42058 12180 42064 12192
rect 42116 12180 42122 12232
rect 42889 12223 42947 12229
rect 42889 12189 42901 12223
rect 42935 12220 42947 12223
rect 43548 12220 43576 12260
rect 43990 12248 43996 12260
rect 44048 12248 44054 12300
rect 50816 12288 50844 12319
rect 51442 12316 51448 12328
rect 51500 12316 51506 12368
rect 51074 12288 51080 12300
rect 50816 12260 51080 12288
rect 51074 12248 51080 12260
rect 51132 12248 51138 12300
rect 42935 12192 43576 12220
rect 43625 12223 43683 12229
rect 42935 12189 42947 12192
rect 42889 12183 42947 12189
rect 43625 12189 43637 12223
rect 43671 12189 43683 12223
rect 43625 12183 43683 12189
rect 44361 12223 44419 12229
rect 44361 12189 44373 12223
rect 44407 12220 44419 12223
rect 45002 12220 45008 12232
rect 44407 12192 45008 12220
rect 44407 12189 44419 12192
rect 44361 12183 44419 12189
rect 34330 12112 34336 12164
rect 34388 12152 34394 12164
rect 37642 12152 37648 12164
rect 34388 12124 37648 12152
rect 34388 12112 34394 12124
rect 37642 12112 37648 12124
rect 37700 12112 37706 12164
rect 38102 12112 38108 12164
rect 38160 12152 38166 12164
rect 39850 12152 39856 12164
rect 38160 12124 39856 12152
rect 38160 12112 38166 12124
rect 39850 12112 39856 12124
rect 39908 12112 39914 12164
rect 40310 12112 40316 12164
rect 40368 12152 40374 12164
rect 40466 12155 40524 12161
rect 40466 12152 40478 12155
rect 40368 12124 40478 12152
rect 40368 12112 40374 12124
rect 40466 12121 40478 12124
rect 40512 12121 40524 12155
rect 43640 12152 43668 12183
rect 45002 12180 45008 12192
rect 45060 12180 45066 12232
rect 45462 12220 45468 12232
rect 45423 12192 45468 12220
rect 45462 12180 45468 12192
rect 45520 12180 45526 12232
rect 45922 12220 45928 12232
rect 45883 12192 45928 12220
rect 45922 12180 45928 12192
rect 45980 12220 45986 12232
rect 49145 12223 49203 12229
rect 49145 12220 49157 12223
rect 45980 12192 49157 12220
rect 45980 12180 45986 12192
rect 49145 12189 49157 12192
rect 49191 12220 49203 12223
rect 49694 12220 49700 12232
rect 49191 12192 49700 12220
rect 49191 12189 49203 12192
rect 49145 12183 49203 12189
rect 49694 12180 49700 12192
rect 49752 12180 49758 12232
rect 49786 12180 49792 12232
rect 49844 12220 49850 12232
rect 50246 12220 50252 12232
rect 49844 12192 50252 12220
rect 49844 12180 49850 12192
rect 50246 12180 50252 12192
rect 50304 12220 50310 12232
rect 50617 12223 50675 12229
rect 50617 12220 50629 12223
rect 50304 12192 50629 12220
rect 50304 12180 50310 12192
rect 50617 12189 50629 12192
rect 50663 12189 50675 12223
rect 51626 12220 51632 12232
rect 51587 12192 51632 12220
rect 50617 12183 50675 12189
rect 51626 12180 51632 12192
rect 51684 12180 51690 12232
rect 51718 12180 51724 12232
rect 51776 12220 51782 12232
rect 52104 12229 52132 12396
rect 52362 12384 52368 12396
rect 52420 12424 52426 12436
rect 55582 12424 55588 12436
rect 52420 12396 55588 12424
rect 52420 12384 52426 12396
rect 55582 12384 55588 12396
rect 55640 12384 55646 12436
rect 56134 12384 56140 12436
rect 56192 12424 56198 12436
rect 56413 12427 56471 12433
rect 56413 12424 56425 12427
rect 56192 12396 56425 12424
rect 56192 12384 56198 12396
rect 56413 12393 56425 12396
rect 56459 12393 56471 12427
rect 56413 12387 56471 12393
rect 56778 12384 56784 12436
rect 56836 12424 56842 12436
rect 57882 12424 57888 12436
rect 56836 12396 57888 12424
rect 56836 12384 56842 12396
rect 57882 12384 57888 12396
rect 57940 12424 57946 12436
rect 57940 12396 58204 12424
rect 57940 12384 57946 12396
rect 54021 12359 54079 12365
rect 54021 12325 54033 12359
rect 54067 12325 54079 12359
rect 54021 12319 54079 12325
rect 54036 12288 54064 12319
rect 54294 12316 54300 12368
rect 54352 12356 54358 12368
rect 57238 12356 57244 12368
rect 54352 12328 57244 12356
rect 54352 12316 54358 12328
rect 57238 12316 57244 12328
rect 57296 12316 57302 12368
rect 58176 12356 58204 12396
rect 58250 12384 58256 12436
rect 58308 12424 58314 12436
rect 59265 12427 59323 12433
rect 59265 12424 59277 12427
rect 58308 12396 59277 12424
rect 58308 12384 58314 12396
rect 59265 12393 59277 12396
rect 59311 12393 59323 12427
rect 63218 12424 63224 12436
rect 63179 12396 63224 12424
rect 59265 12387 59323 12393
rect 63218 12384 63224 12396
rect 63276 12384 63282 12436
rect 63770 12384 63776 12436
rect 63828 12424 63834 12436
rect 63957 12427 64015 12433
rect 63957 12424 63969 12427
rect 63828 12396 63969 12424
rect 63828 12384 63834 12396
rect 63957 12393 63969 12396
rect 64003 12393 64015 12427
rect 63957 12387 64015 12393
rect 64782 12384 64788 12436
rect 64840 12424 64846 12436
rect 64969 12427 65027 12433
rect 64969 12424 64981 12427
rect 64840 12396 64981 12424
rect 64840 12384 64846 12396
rect 64969 12393 64981 12396
rect 65015 12393 65027 12427
rect 64969 12387 65027 12393
rect 68646 12384 68652 12436
rect 68704 12424 68710 12436
rect 68833 12427 68891 12433
rect 68833 12424 68845 12427
rect 68704 12396 68845 12424
rect 68704 12384 68710 12396
rect 68833 12393 68845 12396
rect 68879 12393 68891 12427
rect 68833 12387 68891 12393
rect 69750 12384 69756 12436
rect 69808 12424 69814 12436
rect 70029 12427 70087 12433
rect 70029 12424 70041 12427
rect 69808 12396 70041 12424
rect 69808 12384 69814 12396
rect 70029 12393 70041 12396
rect 70075 12393 70087 12427
rect 70029 12387 70087 12393
rect 71774 12384 71780 12436
rect 71832 12424 71838 12436
rect 72421 12427 72479 12433
rect 72421 12424 72433 12427
rect 71832 12396 72433 12424
rect 71832 12384 71838 12396
rect 72421 12393 72433 12396
rect 72467 12424 72479 12427
rect 73062 12424 73068 12436
rect 72467 12396 73068 12424
rect 72467 12393 72479 12396
rect 72421 12387 72479 12393
rect 73062 12384 73068 12396
rect 73120 12384 73126 12436
rect 75362 12424 75368 12436
rect 73172 12396 74948 12424
rect 75323 12396 75368 12424
rect 61010 12356 61016 12368
rect 58176 12328 61016 12356
rect 61010 12316 61016 12328
rect 61068 12316 61074 12368
rect 62393 12359 62451 12365
rect 62393 12325 62405 12359
rect 62439 12356 62451 12359
rect 66162 12356 66168 12368
rect 62439 12328 66168 12356
rect 62439 12325 62451 12328
rect 62393 12319 62451 12325
rect 66162 12316 66168 12328
rect 66220 12316 66226 12368
rect 66625 12359 66683 12365
rect 66625 12325 66637 12359
rect 66671 12356 66683 12359
rect 69106 12356 69112 12368
rect 66671 12328 69112 12356
rect 66671 12325 66683 12328
rect 66625 12319 66683 12325
rect 69106 12316 69112 12328
rect 69164 12356 69170 12368
rect 69934 12356 69940 12368
rect 69164 12328 69940 12356
rect 69164 12316 69170 12328
rect 69934 12316 69940 12328
rect 69992 12356 69998 12368
rect 69992 12328 70394 12356
rect 69992 12316 69998 12328
rect 56686 12288 56692 12300
rect 54036 12260 56692 12288
rect 56686 12248 56692 12260
rect 56744 12248 56750 12300
rect 56781 12291 56839 12297
rect 56781 12257 56793 12291
rect 56827 12288 56839 12291
rect 57146 12288 57152 12300
rect 56827 12260 57152 12288
rect 56827 12257 56839 12260
rect 56781 12251 56839 12257
rect 57146 12248 57152 12260
rect 57204 12248 57210 12300
rect 67910 12248 67916 12300
rect 67968 12288 67974 12300
rect 67968 12260 69888 12288
rect 67968 12248 67974 12260
rect 52089 12223 52147 12229
rect 52089 12220 52101 12223
rect 51776 12192 52101 12220
rect 51776 12180 51782 12192
rect 52089 12189 52101 12192
rect 52135 12189 52147 12223
rect 52089 12183 52147 12189
rect 54205 12223 54263 12229
rect 54205 12189 54217 12223
rect 54251 12220 54263 12223
rect 54294 12220 54300 12232
rect 54251 12192 54300 12220
rect 54251 12189 54263 12192
rect 54205 12183 54263 12189
rect 54294 12180 54300 12192
rect 54352 12180 54358 12232
rect 54846 12220 54852 12232
rect 54404 12192 54852 12220
rect 40466 12115 40524 12121
rect 41386 12124 43668 12152
rect 46192 12155 46250 12161
rect 30984 12056 32536 12084
rect 33505 12087 33563 12093
rect 30984 12044 30990 12056
rect 33505 12053 33517 12087
rect 33551 12084 33563 12087
rect 33686 12084 33692 12096
rect 33551 12056 33692 12084
rect 33551 12053 33563 12056
rect 33505 12047 33563 12053
rect 33686 12044 33692 12056
rect 33744 12084 33750 12096
rect 33962 12084 33968 12096
rect 33744 12056 33968 12084
rect 33744 12044 33750 12056
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 34882 12044 34888 12096
rect 34940 12084 34946 12096
rect 41386 12084 41414 12124
rect 46192 12121 46204 12155
rect 46238 12152 46250 12155
rect 48774 12152 48780 12164
rect 46238 12124 48780 12152
rect 46238 12121 46250 12124
rect 46192 12115 46250 12121
rect 48774 12112 48780 12124
rect 48832 12112 48838 12164
rect 48900 12155 48958 12161
rect 48900 12121 48912 12155
rect 48946 12152 48958 12155
rect 50154 12152 50160 12164
rect 48946 12124 50160 12152
rect 48946 12121 48958 12124
rect 48900 12115 48958 12121
rect 50154 12112 50160 12124
rect 50212 12112 50218 12164
rect 51994 12152 52000 12164
rect 51046 12124 52000 12152
rect 34940 12056 41414 12084
rect 41601 12087 41659 12093
rect 34940 12044 34946 12056
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 42150 12084 42156 12096
rect 41647 12056 42156 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 42150 12044 42156 12056
rect 42208 12044 42214 12096
rect 42702 12044 42708 12096
rect 42760 12084 42766 12096
rect 42886 12084 42892 12096
rect 42760 12056 42892 12084
rect 42760 12044 42766 12056
rect 42886 12044 42892 12056
rect 42944 12044 42950 12096
rect 43073 12087 43131 12093
rect 43073 12053 43085 12087
rect 43119 12084 43131 12087
rect 44082 12084 44088 12096
rect 43119 12056 44088 12084
rect 43119 12053 43131 12056
rect 43073 12047 43131 12053
rect 44082 12044 44088 12056
rect 44140 12044 44146 12096
rect 45281 12087 45339 12093
rect 45281 12053 45293 12087
rect 45327 12084 45339 12087
rect 46658 12084 46664 12096
rect 45327 12056 46664 12084
rect 45327 12053 45339 12056
rect 45281 12047 45339 12053
rect 46658 12044 46664 12056
rect 46716 12044 46722 12096
rect 47302 12084 47308 12096
rect 47263 12056 47308 12084
rect 47302 12044 47308 12056
rect 47360 12044 47366 12096
rect 47762 12084 47768 12096
rect 47675 12056 47768 12084
rect 47762 12044 47768 12056
rect 47820 12084 47826 12096
rect 51046 12084 51074 12124
rect 51994 12112 52000 12124
rect 52052 12112 52058 12164
rect 52356 12155 52414 12161
rect 52356 12121 52368 12155
rect 52402 12152 52414 12155
rect 53006 12152 53012 12164
rect 52402 12124 53012 12152
rect 52402 12121 52414 12124
rect 52356 12115 52414 12121
rect 53006 12112 53012 12124
rect 53064 12112 53070 12164
rect 54404 12152 54432 12192
rect 54846 12180 54852 12192
rect 54904 12180 54910 12232
rect 55674 12220 55680 12232
rect 55635 12192 55680 12220
rect 55674 12180 55680 12192
rect 55732 12180 55738 12232
rect 55861 12223 55919 12229
rect 55861 12189 55873 12223
rect 55907 12220 55919 12223
rect 55950 12220 55956 12232
rect 55907 12192 55956 12220
rect 55907 12189 55919 12192
rect 55861 12183 55919 12189
rect 55950 12180 55956 12192
rect 56008 12180 56014 12232
rect 56042 12180 56048 12232
rect 56100 12220 56106 12232
rect 56318 12220 56324 12232
rect 56100 12192 56324 12220
rect 56100 12180 56106 12192
rect 56318 12180 56324 12192
rect 56376 12180 56382 12232
rect 56597 12223 56655 12229
rect 56597 12189 56609 12223
rect 56643 12220 56655 12223
rect 57054 12220 57060 12232
rect 56643 12192 57060 12220
rect 56643 12189 56655 12192
rect 56597 12183 56655 12189
rect 57054 12180 57060 12192
rect 57112 12180 57118 12232
rect 57238 12220 57244 12232
rect 57199 12192 57244 12220
rect 57238 12180 57244 12192
rect 57296 12180 57302 12232
rect 57330 12180 57336 12232
rect 57388 12220 57394 12232
rect 59449 12223 59507 12229
rect 59449 12220 59461 12223
rect 57388 12192 59461 12220
rect 57388 12180 57394 12192
rect 59449 12189 59461 12192
rect 59495 12189 59507 12223
rect 59449 12183 59507 12189
rect 59538 12180 59544 12232
rect 59596 12220 59602 12232
rect 61010 12220 61016 12232
rect 59596 12192 59641 12220
rect 60971 12192 61016 12220
rect 59596 12180 59602 12192
rect 61010 12180 61016 12192
rect 61068 12180 61074 12232
rect 62390 12220 62396 12232
rect 61212 12192 62396 12220
rect 53116 12124 54432 12152
rect 54757 12155 54815 12161
rect 47820 12056 51074 12084
rect 51445 12087 51503 12093
rect 47820 12044 47826 12056
rect 51445 12053 51457 12087
rect 51491 12084 51503 12087
rect 53116 12084 53144 12124
rect 54757 12121 54769 12155
rect 54803 12152 54815 12155
rect 57508 12155 57566 12161
rect 54803 12124 55812 12152
rect 54803 12121 54815 12124
rect 54757 12115 54815 12121
rect 51491 12056 53144 12084
rect 53469 12087 53527 12093
rect 51491 12053 51503 12056
rect 51445 12047 51503 12053
rect 53469 12053 53481 12087
rect 53515 12084 53527 12087
rect 54570 12084 54576 12096
rect 53515 12056 54576 12084
rect 53515 12053 53527 12056
rect 53469 12047 53527 12053
rect 54570 12044 54576 12056
rect 54628 12044 54634 12096
rect 54849 12087 54907 12093
rect 54849 12053 54861 12087
rect 54895 12084 54907 12087
rect 55306 12084 55312 12096
rect 54895 12056 55312 12084
rect 54895 12053 54907 12056
rect 54849 12047 54907 12053
rect 55306 12044 55312 12056
rect 55364 12044 55370 12096
rect 55490 12084 55496 12096
rect 55451 12056 55496 12084
rect 55490 12044 55496 12056
rect 55548 12044 55554 12096
rect 55784 12084 55812 12124
rect 57508 12121 57520 12155
rect 57554 12152 57566 12155
rect 61212 12152 61240 12192
rect 62390 12180 62396 12192
rect 62448 12180 62454 12232
rect 62482 12180 62488 12232
rect 62540 12220 62546 12232
rect 63037 12223 63095 12229
rect 63037 12220 63049 12223
rect 62540 12192 63049 12220
rect 62540 12180 62546 12192
rect 63037 12189 63049 12192
rect 63083 12189 63095 12223
rect 63037 12183 63095 12189
rect 63773 12223 63831 12229
rect 63773 12189 63785 12223
rect 63819 12189 63831 12223
rect 63773 12183 63831 12189
rect 65153 12223 65211 12229
rect 65153 12189 65165 12223
rect 65199 12220 65211 12223
rect 65794 12220 65800 12232
rect 65199 12192 65800 12220
rect 65199 12189 65211 12192
rect 65153 12183 65211 12189
rect 57554 12124 61240 12152
rect 61280 12155 61338 12161
rect 57554 12121 57566 12124
rect 57508 12115 57566 12121
rect 61280 12121 61292 12155
rect 61326 12152 61338 12155
rect 61654 12152 61660 12164
rect 61326 12124 61660 12152
rect 61326 12121 61338 12124
rect 61280 12115 61338 12121
rect 61654 12112 61660 12124
rect 61712 12112 61718 12164
rect 63788 12152 63816 12183
rect 65794 12180 65800 12192
rect 65852 12180 65858 12232
rect 69860 12229 69888 12260
rect 67729 12223 67787 12229
rect 67729 12189 67741 12223
rect 67775 12220 67787 12223
rect 69017 12223 69075 12229
rect 69017 12220 69029 12223
rect 67775 12192 69029 12220
rect 67775 12189 67787 12192
rect 67729 12183 67787 12189
rect 69017 12189 69029 12192
rect 69063 12189 69075 12223
rect 69017 12183 69075 12189
rect 69845 12223 69903 12229
rect 69845 12189 69857 12223
rect 69891 12189 69903 12223
rect 70366 12220 70394 12328
rect 72326 12316 72332 12368
rect 72384 12356 72390 12368
rect 73172 12356 73200 12396
rect 72384 12328 73200 12356
rect 74920 12356 74948 12396
rect 75362 12384 75368 12396
rect 75420 12384 75426 12436
rect 76190 12384 76196 12436
rect 76248 12424 76254 12436
rect 77478 12424 77484 12436
rect 76248 12396 77484 12424
rect 76248 12384 76254 12396
rect 77478 12384 77484 12396
rect 77536 12384 77542 12436
rect 77754 12424 77760 12436
rect 77715 12396 77760 12424
rect 77754 12384 77760 12396
rect 77812 12384 77818 12436
rect 84746 12424 84752 12436
rect 78232 12396 84752 12424
rect 78232 12356 78260 12396
rect 84746 12384 84752 12396
rect 84804 12384 84810 12436
rect 85206 12384 85212 12436
rect 85264 12424 85270 12436
rect 85393 12427 85451 12433
rect 85393 12424 85405 12427
rect 85264 12396 85405 12424
rect 85264 12384 85270 12396
rect 85393 12393 85405 12396
rect 85439 12393 85451 12427
rect 85393 12387 85451 12393
rect 85758 12384 85764 12436
rect 85816 12424 85822 12436
rect 86589 12427 86647 12433
rect 86589 12424 86601 12427
rect 85816 12396 86601 12424
rect 85816 12384 85822 12396
rect 86589 12393 86601 12396
rect 86635 12393 86647 12427
rect 86589 12387 86647 12393
rect 87322 12384 87328 12436
rect 87380 12424 87386 12436
rect 87785 12427 87843 12433
rect 87785 12424 87797 12427
rect 87380 12396 87797 12424
rect 87380 12384 87386 12396
rect 87785 12393 87797 12396
rect 87831 12393 87843 12427
rect 87785 12387 87843 12393
rect 87874 12384 87880 12436
rect 87932 12424 87938 12436
rect 87932 12396 96200 12424
rect 87932 12384 87938 12396
rect 74920 12328 78260 12356
rect 72384 12316 72390 12328
rect 79686 12316 79692 12368
rect 79744 12356 79750 12368
rect 80514 12356 80520 12368
rect 79744 12328 80520 12356
rect 79744 12316 79750 12328
rect 80514 12316 80520 12328
rect 80572 12316 80578 12368
rect 82170 12316 82176 12368
rect 82228 12356 82234 12368
rect 88150 12356 88156 12368
rect 82228 12328 88156 12356
rect 82228 12316 82234 12328
rect 88150 12316 88156 12328
rect 88208 12316 88214 12368
rect 89162 12316 89168 12368
rect 89220 12356 89226 12368
rect 89809 12359 89867 12365
rect 89809 12356 89821 12359
rect 89220 12328 89821 12356
rect 89220 12316 89226 12328
rect 89809 12325 89821 12328
rect 89855 12325 89867 12359
rect 89809 12319 89867 12325
rect 89898 12316 89904 12368
rect 89956 12356 89962 12368
rect 90545 12359 90603 12365
rect 90545 12356 90557 12359
rect 89956 12328 90557 12356
rect 89956 12316 89962 12328
rect 90545 12325 90557 12328
rect 90591 12325 90603 12359
rect 90545 12319 90603 12325
rect 75914 12248 75920 12300
rect 75972 12288 75978 12300
rect 76653 12291 76711 12297
rect 76653 12288 76665 12291
rect 75972 12260 76665 12288
rect 75972 12248 75978 12260
rect 76653 12257 76665 12260
rect 76699 12288 76711 12291
rect 76742 12288 76748 12300
rect 76699 12260 76748 12288
rect 76699 12257 76711 12260
rect 76653 12251 76711 12257
rect 76742 12248 76748 12260
rect 76800 12248 76806 12300
rect 77386 12248 77392 12300
rect 77444 12288 77450 12300
rect 77754 12288 77760 12300
rect 77444 12260 77760 12288
rect 77444 12248 77450 12260
rect 77754 12248 77760 12260
rect 77812 12248 77818 12300
rect 81253 12291 81311 12297
rect 81253 12257 81265 12291
rect 81299 12288 81311 12291
rect 81299 12260 82032 12288
rect 81299 12257 81311 12260
rect 81253 12251 81311 12257
rect 72881 12223 72939 12229
rect 72881 12220 72893 12223
rect 70366 12192 72893 12220
rect 69845 12183 69903 12189
rect 72881 12189 72893 12192
rect 72927 12220 72939 12223
rect 73154 12220 73160 12232
rect 72927 12192 73160 12220
rect 72927 12189 72939 12192
rect 72881 12183 72939 12189
rect 62224 12124 63816 12152
rect 67177 12155 67235 12161
rect 56778 12084 56784 12096
rect 55784 12056 56784 12084
rect 56778 12044 56784 12056
rect 56836 12044 56842 12096
rect 58621 12087 58679 12093
rect 58621 12053 58633 12087
rect 58667 12084 58679 12087
rect 62224 12084 62252 12124
rect 67177 12121 67189 12155
rect 67223 12152 67235 12155
rect 68830 12152 68836 12164
rect 67223 12124 68836 12152
rect 67223 12121 67235 12124
rect 67177 12115 67235 12121
rect 68830 12112 68836 12124
rect 68888 12112 68894 12164
rect 69032 12152 69060 12183
rect 73154 12180 73160 12192
rect 73212 12220 73218 12232
rect 73985 12223 74043 12229
rect 73985 12220 73997 12223
rect 73212 12192 73997 12220
rect 73212 12180 73218 12192
rect 73985 12189 73997 12192
rect 74031 12189 74043 12223
rect 74252 12223 74310 12229
rect 74252 12220 74264 12223
rect 73985 12183 74043 12189
rect 74184 12192 74264 12220
rect 73525 12155 73583 12161
rect 69032 12124 73476 12152
rect 58667 12056 62252 12084
rect 66073 12087 66131 12093
rect 58667 12053 58679 12056
rect 58621 12047 58679 12053
rect 66073 12053 66085 12087
rect 66119 12084 66131 12087
rect 66162 12084 66168 12096
rect 66119 12056 66168 12084
rect 66119 12053 66131 12056
rect 66073 12047 66131 12053
rect 66162 12044 66168 12056
rect 66220 12084 66226 12096
rect 66806 12084 66812 12096
rect 66220 12056 66812 12084
rect 66220 12044 66226 12056
rect 66806 12044 66812 12056
rect 66864 12044 66870 12096
rect 68281 12087 68339 12093
rect 68281 12053 68293 12087
rect 68327 12084 68339 12087
rect 68738 12084 68744 12096
rect 68327 12056 68744 12084
rect 68327 12053 68339 12056
rect 68281 12047 68339 12053
rect 68738 12044 68744 12056
rect 68796 12044 68802 12096
rect 71041 12087 71099 12093
rect 71041 12053 71053 12087
rect 71087 12084 71099 12087
rect 71130 12084 71136 12096
rect 71087 12056 71136 12084
rect 71087 12053 71099 12056
rect 71041 12047 71099 12053
rect 71130 12044 71136 12056
rect 71188 12044 71194 12096
rect 71682 12084 71688 12096
rect 71643 12056 71688 12084
rect 71682 12044 71688 12056
rect 71740 12044 71746 12096
rect 73448 12084 73476 12124
rect 73525 12121 73537 12155
rect 73571 12152 73583 12155
rect 74184 12152 74212 12192
rect 74252 12189 74264 12192
rect 74298 12220 74310 12223
rect 78582 12220 78588 12232
rect 74298 12192 78588 12220
rect 74298 12189 74310 12192
rect 74252 12183 74310 12189
rect 78582 12180 78588 12192
rect 78640 12180 78646 12232
rect 79137 12223 79195 12229
rect 79137 12189 79149 12223
rect 79183 12220 79195 12223
rect 80514 12220 80520 12232
rect 79183 12192 80520 12220
rect 79183 12189 79195 12192
rect 79137 12183 79195 12189
rect 77294 12152 77300 12164
rect 73571 12124 74212 12152
rect 77255 12124 77300 12152
rect 73571 12121 73583 12124
rect 73525 12115 73583 12121
rect 77294 12112 77300 12124
rect 77352 12112 77358 12164
rect 78870 12155 78928 12161
rect 78870 12152 78882 12155
rect 77404 12124 78882 12152
rect 75270 12084 75276 12096
rect 73448 12056 75276 12084
rect 75270 12044 75276 12056
rect 75328 12044 75334 12096
rect 75546 12044 75552 12096
rect 75604 12084 75610 12096
rect 77404 12084 77432 12124
rect 78870 12121 78882 12124
rect 78916 12121 78928 12155
rect 79152 12152 79180 12183
rect 80514 12180 80520 12192
rect 80572 12180 80578 12232
rect 81437 12223 81495 12229
rect 81437 12189 81449 12223
rect 81483 12220 81495 12223
rect 81710 12220 81716 12232
rect 81483 12192 81716 12220
rect 81483 12189 81495 12192
rect 81437 12183 81495 12189
rect 81710 12180 81716 12192
rect 81768 12180 81774 12232
rect 82004 12220 82032 12260
rect 83090 12248 83096 12300
rect 83148 12288 83154 12300
rect 83737 12291 83795 12297
rect 83737 12288 83749 12291
rect 83148 12260 83749 12288
rect 83148 12248 83154 12260
rect 83737 12257 83749 12260
rect 83783 12288 83795 12291
rect 84102 12288 84108 12300
rect 83783 12260 84108 12288
rect 83783 12257 83795 12260
rect 83737 12251 83795 12257
rect 84102 12248 84108 12260
rect 84160 12248 84166 12300
rect 85390 12248 85396 12300
rect 85448 12288 85454 12300
rect 87141 12291 87199 12297
rect 87141 12288 87153 12291
rect 85448 12260 87153 12288
rect 85448 12248 85454 12260
rect 82078 12220 82084 12232
rect 81991 12192 82084 12220
rect 82078 12180 82084 12192
rect 82136 12180 82142 12232
rect 85592 12229 85620 12260
rect 87141 12257 87153 12260
rect 87187 12257 87199 12291
rect 87141 12251 87199 12257
rect 89530 12248 89536 12300
rect 89588 12288 89594 12300
rect 90082 12288 90088 12300
rect 89588 12260 90088 12288
rect 89588 12248 89594 12260
rect 90082 12248 90088 12260
rect 90140 12248 90146 12300
rect 90174 12248 90180 12300
rect 90232 12288 90238 12300
rect 93026 12288 93032 12300
rect 90232 12260 90496 12288
rect 90232 12248 90238 12260
rect 85577 12223 85635 12229
rect 85577 12189 85589 12223
rect 85623 12189 85635 12223
rect 86402 12220 86408 12232
rect 86363 12192 86408 12220
rect 85577 12183 85635 12189
rect 86402 12180 86408 12192
rect 86460 12180 86466 12232
rect 89162 12220 89168 12232
rect 89123 12192 89168 12220
rect 89162 12180 89168 12192
rect 89220 12220 89226 12232
rect 89438 12220 89444 12232
rect 89220 12192 89444 12220
rect 89220 12180 89226 12192
rect 89438 12180 89444 12192
rect 89496 12180 89502 12232
rect 89625 12223 89683 12229
rect 89625 12189 89637 12223
rect 89671 12189 89683 12223
rect 90358 12220 90364 12232
rect 90319 12192 90364 12220
rect 89625 12183 89683 12189
rect 78870 12115 78928 12121
rect 79060 12124 79180 12152
rect 75604 12056 77432 12084
rect 75604 12044 75610 12056
rect 77478 12044 77484 12096
rect 77536 12084 77542 12096
rect 79060 12084 79088 12124
rect 82446 12112 82452 12164
rect 82504 12152 82510 12164
rect 82504 12124 84608 12152
rect 82504 12112 82510 12124
rect 77536 12056 79088 12084
rect 77536 12044 77542 12056
rect 79134 12044 79140 12096
rect 79192 12084 79198 12096
rect 80698 12084 80704 12096
rect 79192 12056 80704 12084
rect 79192 12044 79198 12056
rect 80698 12044 80704 12056
rect 80756 12044 80762 12096
rect 81618 12084 81624 12096
rect 81579 12056 81624 12084
rect 81618 12044 81624 12056
rect 81676 12044 81682 12096
rect 81710 12044 81716 12096
rect 81768 12084 81774 12096
rect 82630 12084 82636 12096
rect 81768 12056 82636 12084
rect 81768 12044 81774 12056
rect 82630 12044 82636 12056
rect 82688 12044 82694 12096
rect 83274 12084 83280 12096
rect 83235 12056 83280 12084
rect 83274 12044 83280 12056
rect 83332 12044 83338 12096
rect 84286 12044 84292 12096
rect 84344 12084 84350 12096
rect 84381 12087 84439 12093
rect 84381 12084 84393 12087
rect 84344 12056 84393 12084
rect 84344 12044 84350 12056
rect 84381 12053 84393 12056
rect 84427 12084 84439 12087
rect 84470 12084 84476 12096
rect 84427 12056 84476 12084
rect 84427 12053 84439 12056
rect 84381 12047 84439 12053
rect 84470 12044 84476 12056
rect 84528 12044 84534 12096
rect 84580 12084 84608 12124
rect 84746 12112 84752 12164
rect 84804 12152 84810 12164
rect 88058 12152 88064 12164
rect 84804 12124 88064 12152
rect 84804 12112 84810 12124
rect 88058 12112 88064 12124
rect 88116 12112 88122 12164
rect 88886 12152 88892 12164
rect 88944 12161 88950 12164
rect 88856 12124 88892 12152
rect 88886 12112 88892 12124
rect 88944 12115 88956 12161
rect 88944 12112 88950 12115
rect 89640 12084 89668 12183
rect 90358 12180 90364 12192
rect 90416 12180 90422 12232
rect 90468 12220 90496 12260
rect 92860 12260 93032 12288
rect 92860 12220 92888 12260
rect 93026 12248 93032 12260
rect 93084 12248 93090 12300
rect 93302 12248 93308 12300
rect 93360 12288 93366 12300
rect 94133 12291 94191 12297
rect 94133 12288 94145 12291
rect 93360 12260 94145 12288
rect 93360 12248 93366 12260
rect 94133 12257 94145 12260
rect 94179 12257 94191 12291
rect 96172 12288 96200 12396
rect 96246 12384 96252 12436
rect 96304 12424 96310 12436
rect 96801 12427 96859 12433
rect 96801 12424 96813 12427
rect 96304 12396 96813 12424
rect 96304 12384 96310 12396
rect 96801 12393 96813 12396
rect 96847 12393 96859 12427
rect 98730 12424 98736 12436
rect 98691 12396 98736 12424
rect 96801 12387 96859 12393
rect 98730 12384 98736 12396
rect 98788 12384 98794 12436
rect 99377 12427 99435 12433
rect 99377 12393 99389 12427
rect 99423 12424 99435 12427
rect 99926 12424 99932 12436
rect 99423 12396 99932 12424
rect 99423 12393 99435 12396
rect 99377 12387 99435 12393
rect 99926 12384 99932 12396
rect 99984 12384 99990 12436
rect 102042 12384 102048 12436
rect 102100 12424 102106 12436
rect 104618 12424 104624 12436
rect 102100 12396 104624 12424
rect 102100 12384 102106 12396
rect 104618 12384 104624 12396
rect 104676 12384 104682 12436
rect 105078 12384 105084 12436
rect 105136 12424 105142 12436
rect 105357 12427 105415 12433
rect 105357 12424 105369 12427
rect 105136 12396 105369 12424
rect 105136 12384 105142 12396
rect 105357 12393 105369 12396
rect 105403 12393 105415 12427
rect 105357 12387 105415 12393
rect 105630 12384 105636 12436
rect 105688 12424 105694 12436
rect 106001 12427 106059 12433
rect 106001 12424 106013 12427
rect 105688 12396 106013 12424
rect 105688 12384 105694 12396
rect 106001 12393 106013 12396
rect 106047 12393 106059 12427
rect 106001 12387 106059 12393
rect 106734 12384 106740 12436
rect 106792 12424 106798 12436
rect 107105 12427 107163 12433
rect 107105 12424 107117 12427
rect 106792 12396 107117 12424
rect 106792 12384 106798 12396
rect 107105 12393 107117 12396
rect 107151 12393 107163 12427
rect 107105 12387 107163 12393
rect 107286 12384 107292 12436
rect 107344 12424 107350 12436
rect 110230 12424 110236 12436
rect 107344 12396 110092 12424
rect 110191 12396 110236 12424
rect 107344 12384 107350 12396
rect 98178 12316 98184 12368
rect 98236 12356 98242 12368
rect 101398 12356 101404 12368
rect 98236 12328 101404 12356
rect 98236 12316 98242 12328
rect 101398 12316 101404 12328
rect 101456 12316 101462 12368
rect 101508 12328 106504 12356
rect 101508 12288 101536 12328
rect 96172 12260 101536 12288
rect 94133 12251 94191 12257
rect 101582 12248 101588 12300
rect 101640 12288 101646 12300
rect 106366 12288 106372 12300
rect 101640 12260 106372 12288
rect 101640 12248 101646 12260
rect 90468 12192 92888 12220
rect 92937 12223 92995 12229
rect 92937 12189 92949 12223
rect 92983 12220 92995 12223
rect 93670 12220 93676 12232
rect 92983 12192 93256 12220
rect 93631 12192 93676 12220
rect 92983 12189 92995 12192
rect 92937 12183 92995 12189
rect 93228 12164 93256 12192
rect 93670 12180 93676 12192
rect 93728 12180 93734 12232
rect 96154 12220 96160 12232
rect 94976 12192 96160 12220
rect 89898 12112 89904 12164
rect 89956 12152 89962 12164
rect 90818 12152 90824 12164
rect 89956 12124 90824 12152
rect 89956 12112 89962 12124
rect 90818 12112 90824 12124
rect 90876 12112 90882 12164
rect 92692 12155 92750 12161
rect 92692 12121 92704 12155
rect 92738 12152 92750 12155
rect 93118 12152 93124 12164
rect 92738 12124 93124 12152
rect 92738 12121 92750 12124
rect 92692 12115 92750 12121
rect 93118 12112 93124 12124
rect 93176 12112 93182 12164
rect 93210 12112 93216 12164
rect 93268 12152 93274 12164
rect 94976 12152 95004 12192
rect 96154 12180 96160 12192
rect 96212 12180 96218 12232
rect 96982 12220 96988 12232
rect 96943 12192 96988 12220
rect 96982 12180 96988 12192
rect 97040 12180 97046 12232
rect 97721 12223 97779 12229
rect 97721 12189 97733 12223
rect 97767 12220 97779 12223
rect 99282 12220 99288 12232
rect 97767 12192 99288 12220
rect 97767 12189 97779 12192
rect 97721 12183 97779 12189
rect 99282 12180 99288 12192
rect 99340 12180 99346 12232
rect 99929 12223 99987 12229
rect 99929 12189 99941 12223
rect 99975 12220 99987 12223
rect 100294 12220 100300 12232
rect 99975 12192 100300 12220
rect 99975 12189 99987 12192
rect 99929 12183 99987 12189
rect 100294 12180 100300 12192
rect 100352 12180 100358 12232
rect 102962 12220 102968 12232
rect 102923 12192 102968 12220
rect 102962 12180 102968 12192
rect 103020 12180 103026 12232
rect 103054 12180 103060 12232
rect 103112 12220 103118 12232
rect 104342 12220 104348 12232
rect 103112 12192 104348 12220
rect 103112 12180 103118 12192
rect 104342 12180 104348 12192
rect 104400 12180 104406 12232
rect 104544 12229 104572 12260
rect 106366 12248 106372 12260
rect 106424 12248 106430 12300
rect 106476 12288 106504 12328
rect 108666 12316 108672 12368
rect 108724 12316 108730 12368
rect 110064 12356 110092 12396
rect 110230 12384 110236 12396
rect 110288 12384 110294 12436
rect 111702 12384 111708 12436
rect 111760 12424 111766 12436
rect 112257 12427 112315 12433
rect 112257 12424 112269 12427
rect 111760 12396 112269 12424
rect 111760 12384 111766 12396
rect 112257 12393 112269 12396
rect 112303 12393 112315 12427
rect 112257 12387 112315 12393
rect 112346 12384 112352 12436
rect 112404 12424 112410 12436
rect 118510 12424 118516 12436
rect 112404 12396 118516 12424
rect 112404 12384 112410 12396
rect 118510 12384 118516 12396
rect 118568 12384 118574 12436
rect 118666 12396 120304 12424
rect 118666 12356 118694 12396
rect 110064 12328 118694 12356
rect 120276 12356 120304 12396
rect 121638 12384 121644 12436
rect 121696 12424 121702 12436
rect 121733 12427 121791 12433
rect 121733 12424 121745 12427
rect 121696 12396 121745 12424
rect 121696 12384 121702 12396
rect 121733 12393 121745 12396
rect 121779 12393 121791 12427
rect 121733 12387 121791 12393
rect 121822 12384 121828 12436
rect 121880 12424 121886 12436
rect 126054 12424 126060 12436
rect 121880 12396 126060 12424
rect 121880 12384 121886 12396
rect 126054 12384 126060 12396
rect 126112 12384 126118 12436
rect 127158 12384 127164 12436
rect 127216 12424 127222 12436
rect 127805 12427 127863 12433
rect 127805 12424 127817 12427
rect 127216 12396 127817 12424
rect 127216 12384 127222 12396
rect 127805 12393 127817 12396
rect 127851 12393 127863 12427
rect 128446 12424 128452 12436
rect 128407 12396 128452 12424
rect 127805 12387 127863 12393
rect 128446 12384 128452 12396
rect 128504 12384 128510 12436
rect 129001 12427 129059 12433
rect 129001 12393 129013 12427
rect 129047 12424 129059 12427
rect 129090 12424 129096 12436
rect 129047 12396 129096 12424
rect 129047 12393 129059 12396
rect 129001 12387 129059 12393
rect 129090 12384 129096 12396
rect 129148 12384 129154 12436
rect 130470 12384 130476 12436
rect 130528 12424 130534 12436
rect 132865 12427 132923 12433
rect 132865 12424 132877 12427
rect 130528 12396 132877 12424
rect 130528 12384 130534 12396
rect 132865 12393 132877 12396
rect 132911 12424 132923 12427
rect 135070 12424 135076 12436
rect 132911 12396 135076 12424
rect 132911 12393 132923 12396
rect 132865 12387 132923 12393
rect 135070 12384 135076 12396
rect 135128 12384 135134 12436
rect 135530 12424 135536 12436
rect 135491 12396 135536 12424
rect 135530 12384 135536 12396
rect 135588 12384 135594 12436
rect 137186 12384 137192 12436
rect 137244 12424 137250 12436
rect 141326 12424 141332 12436
rect 137244 12396 141188 12424
rect 141287 12396 141332 12424
rect 137244 12384 137250 12396
rect 122469 12359 122527 12365
rect 122469 12356 122481 12359
rect 120276 12328 122481 12356
rect 122469 12325 122481 12328
rect 122515 12325 122527 12359
rect 125594 12356 125600 12368
rect 122469 12319 122527 12325
rect 123864 12328 125600 12356
rect 108684 12288 108712 12316
rect 114278 12288 114284 12300
rect 106476 12260 108712 12288
rect 110432 12260 114284 12288
rect 104529 12223 104587 12229
rect 104529 12189 104541 12223
rect 104575 12189 104587 12223
rect 104529 12183 104587 12189
rect 104618 12180 104624 12232
rect 104676 12220 104682 12232
rect 105173 12223 105231 12229
rect 105173 12220 105185 12223
rect 104676 12192 105185 12220
rect 104676 12180 104682 12192
rect 105173 12189 105185 12192
rect 105219 12189 105231 12223
rect 106182 12220 106188 12232
rect 106143 12192 106188 12220
rect 105173 12183 105231 12189
rect 106182 12180 106188 12192
rect 106240 12180 106246 12232
rect 107286 12220 107292 12232
rect 107247 12192 107292 12220
rect 107286 12180 107292 12192
rect 107344 12180 107350 12232
rect 107562 12180 107568 12232
rect 107620 12220 107626 12232
rect 110432 12229 110460 12260
rect 114278 12248 114284 12260
rect 114336 12248 114342 12300
rect 117869 12291 117927 12297
rect 117869 12288 117881 12291
rect 115400 12260 117881 12288
rect 109681 12223 109739 12229
rect 109681 12220 109693 12223
rect 107620 12192 109693 12220
rect 107620 12180 107626 12192
rect 109681 12189 109693 12192
rect 109727 12189 109739 12223
rect 109681 12183 109739 12189
rect 110417 12223 110475 12229
rect 110417 12189 110429 12223
rect 110463 12189 110475 12223
rect 110874 12220 110880 12232
rect 110835 12192 110880 12220
rect 110417 12183 110475 12189
rect 93268 12124 95004 12152
rect 95912 12155 95970 12161
rect 93268 12112 93274 12124
rect 95912 12121 95924 12155
rect 95958 12152 95970 12155
rect 98178 12152 98184 12164
rect 95958 12124 98184 12152
rect 95958 12121 95970 12124
rect 95912 12115 95970 12121
rect 98178 12112 98184 12124
rect 98236 12112 98242 12164
rect 101030 12112 101036 12164
rect 101088 12152 101094 12164
rect 109402 12152 109408 12164
rect 109460 12161 109466 12164
rect 101088 12124 103744 12152
rect 101088 12112 101094 12124
rect 91554 12084 91560 12096
rect 84580 12056 89668 12084
rect 91515 12056 91560 12084
rect 91554 12044 91560 12056
rect 91612 12044 91618 12096
rect 91830 12044 91836 12096
rect 91888 12084 91894 12096
rect 93489 12087 93547 12093
rect 93489 12084 93501 12087
rect 91888 12056 93501 12084
rect 91888 12044 91894 12056
rect 93489 12053 93501 12056
rect 93535 12053 93547 12087
rect 94774 12084 94780 12096
rect 94735 12056 94780 12084
rect 93489 12047 93547 12053
rect 94774 12044 94780 12056
rect 94832 12044 94838 12096
rect 96522 12044 96528 12096
rect 96580 12084 96586 12096
rect 97537 12087 97595 12093
rect 97537 12084 97549 12087
rect 96580 12056 97549 12084
rect 96580 12044 96586 12056
rect 97537 12053 97549 12056
rect 97583 12053 97595 12087
rect 100386 12084 100392 12096
rect 100347 12056 100392 12084
rect 97537 12047 97595 12053
rect 100386 12044 100392 12056
rect 100444 12044 100450 12096
rect 101306 12084 101312 12096
rect 101219 12056 101312 12084
rect 101306 12044 101312 12056
rect 101364 12084 101370 12096
rect 101490 12084 101496 12096
rect 101364 12056 101496 12084
rect 101364 12044 101370 12056
rect 101490 12044 101496 12056
rect 101548 12044 101554 12096
rect 101950 12084 101956 12096
rect 101911 12056 101956 12084
rect 101950 12044 101956 12056
rect 102008 12044 102014 12096
rect 102318 12044 102324 12096
rect 102376 12084 102382 12096
rect 102781 12087 102839 12093
rect 102781 12084 102793 12087
rect 102376 12056 102793 12084
rect 102376 12044 102382 12056
rect 102781 12053 102793 12056
rect 102827 12053 102839 12087
rect 102781 12047 102839 12053
rect 103517 12087 103575 12093
rect 103517 12053 103529 12087
rect 103563 12084 103575 12087
rect 103606 12084 103612 12096
rect 103563 12056 103612 12084
rect 103563 12053 103575 12056
rect 103517 12047 103575 12053
rect 103606 12044 103612 12056
rect 103664 12044 103670 12096
rect 103716 12084 103744 12124
rect 104544 12124 109034 12152
rect 109372 12124 109408 12152
rect 104544 12084 104572 12124
rect 103716 12056 104572 12084
rect 104713 12087 104771 12093
rect 104713 12053 104725 12087
rect 104759 12084 104771 12087
rect 105630 12084 105636 12096
rect 104759 12056 105636 12084
rect 104759 12053 104771 12056
rect 104713 12047 104771 12053
rect 105630 12044 105636 12056
rect 105688 12044 105694 12096
rect 105814 12044 105820 12096
rect 105872 12084 105878 12096
rect 107841 12087 107899 12093
rect 107841 12084 107853 12087
rect 105872 12056 107853 12084
rect 105872 12044 105878 12056
rect 107841 12053 107853 12056
rect 107887 12084 107899 12087
rect 107930 12084 107936 12096
rect 107887 12056 107936 12084
rect 107887 12053 107899 12056
rect 107841 12047 107899 12053
rect 107930 12044 107936 12056
rect 107988 12044 107994 12096
rect 108022 12044 108028 12096
rect 108080 12084 108086 12096
rect 108301 12087 108359 12093
rect 108301 12084 108313 12087
rect 108080 12056 108313 12084
rect 108080 12044 108086 12056
rect 108301 12053 108313 12056
rect 108347 12053 108359 12087
rect 109006 12084 109034 12124
rect 109402 12112 109408 12124
rect 109460 12115 109472 12161
rect 109696 12152 109724 12183
rect 110874 12180 110880 12192
rect 110932 12180 110938 12232
rect 111061 12223 111119 12229
rect 111061 12189 111073 12223
rect 111107 12220 111119 12223
rect 111242 12220 111248 12232
rect 111107 12192 111248 12220
rect 111107 12189 111119 12192
rect 111061 12183 111119 12189
rect 111242 12180 111248 12192
rect 111300 12180 111306 12232
rect 112441 12223 112499 12229
rect 112441 12189 112453 12223
rect 112487 12220 112499 12223
rect 114830 12220 114836 12232
rect 112487 12192 114836 12220
rect 112487 12189 112499 12192
rect 112441 12183 112499 12189
rect 114830 12180 114836 12192
rect 114888 12180 114894 12232
rect 115400 12229 115428 12260
rect 117869 12257 117881 12260
rect 117915 12288 117927 12291
rect 117958 12288 117964 12300
rect 117915 12260 117964 12288
rect 117915 12257 117927 12260
rect 117869 12251 117927 12257
rect 117958 12248 117964 12260
rect 118016 12248 118022 12300
rect 120261 12291 120319 12297
rect 120261 12257 120273 12291
rect 120307 12288 120319 12291
rect 122742 12288 122748 12300
rect 120307 12260 122748 12288
rect 120307 12257 120319 12260
rect 120261 12251 120319 12257
rect 115385 12223 115443 12229
rect 115385 12189 115397 12223
rect 115431 12189 115443 12223
rect 116486 12220 116492 12232
rect 116447 12192 116492 12220
rect 115385 12183 115443 12189
rect 116486 12180 116492 12192
rect 116544 12180 116550 12232
rect 117222 12180 117228 12232
rect 117280 12220 117286 12232
rect 118510 12220 118516 12232
rect 117280 12192 118516 12220
rect 117280 12180 117286 12192
rect 118510 12180 118516 12192
rect 118568 12180 118574 12232
rect 120276 12220 120304 12251
rect 122742 12248 122748 12260
rect 122800 12248 122806 12300
rect 123864 12288 123892 12328
rect 125594 12316 125600 12328
rect 125652 12316 125658 12368
rect 126790 12316 126796 12368
rect 126848 12356 126854 12368
rect 127986 12356 127992 12368
rect 126848 12328 127992 12356
rect 126848 12316 126854 12328
rect 127986 12316 127992 12328
rect 128044 12316 128050 12368
rect 133874 12356 133880 12368
rect 129568 12328 133880 12356
rect 128446 12288 128452 12300
rect 123772 12260 123892 12288
rect 124600 12260 128452 12288
rect 118666 12192 120304 12220
rect 112530 12152 112536 12164
rect 109696 12124 112536 12152
rect 109460 12112 109466 12115
rect 112530 12112 112536 12124
rect 112588 12152 112594 12164
rect 112993 12155 113051 12161
rect 112993 12152 113005 12155
rect 112588 12124 113005 12152
rect 112588 12112 112594 12124
rect 112993 12121 113005 12124
rect 113039 12152 113051 12155
rect 115290 12152 115296 12164
rect 113039 12124 115296 12152
rect 113039 12121 113051 12124
rect 112993 12115 113051 12121
rect 115290 12112 115296 12124
rect 115348 12152 115354 12164
rect 118666 12152 118694 12192
rect 120442 12180 120448 12232
rect 120500 12220 120506 12232
rect 121822 12220 121828 12232
rect 120500 12192 121828 12220
rect 120500 12180 120506 12192
rect 121822 12180 121828 12192
rect 121880 12180 121886 12232
rect 121917 12223 121975 12229
rect 121917 12189 121929 12223
rect 121963 12220 121975 12223
rect 123772 12220 123800 12260
rect 121963 12192 123800 12220
rect 121963 12189 121975 12192
rect 121917 12183 121975 12189
rect 123846 12180 123852 12232
rect 123904 12220 123910 12232
rect 124600 12229 124628 12260
rect 128446 12248 128452 12260
rect 128504 12248 128510 12300
rect 128538 12248 128544 12300
rect 128596 12288 128602 12300
rect 129568 12288 129596 12328
rect 133874 12316 133880 12328
rect 133932 12316 133938 12368
rect 131758 12288 131764 12300
rect 128596 12260 129596 12288
rect 129844 12260 131764 12288
rect 128596 12248 128602 12260
rect 124585 12223 124643 12229
rect 123904 12192 123949 12220
rect 123904 12180 123910 12192
rect 124585 12189 124597 12223
rect 124631 12189 124643 12223
rect 124585 12183 124643 12189
rect 125502 12180 125508 12232
rect 125560 12220 125566 12232
rect 125689 12223 125747 12229
rect 125689 12220 125701 12223
rect 125560 12192 125701 12220
rect 125560 12180 125566 12192
rect 125689 12189 125701 12192
rect 125735 12220 125747 12223
rect 126514 12220 126520 12232
rect 125735 12192 126520 12220
rect 125735 12189 125747 12192
rect 125689 12183 125747 12189
rect 126514 12180 126520 12192
rect 126572 12180 126578 12232
rect 127434 12180 127440 12232
rect 127492 12220 127498 12232
rect 127621 12223 127679 12229
rect 127621 12220 127633 12223
rect 127492 12192 127633 12220
rect 127492 12180 127498 12192
rect 127621 12189 127633 12192
rect 127667 12189 127679 12223
rect 127621 12183 127679 12189
rect 127894 12180 127900 12232
rect 127952 12220 127958 12232
rect 129844 12220 129872 12260
rect 131758 12248 131764 12260
rect 131816 12248 131822 12300
rect 137005 12291 137063 12297
rect 137005 12288 137017 12291
rect 136008 12260 137017 12288
rect 130010 12220 130016 12232
rect 127952 12192 129872 12220
rect 129971 12192 130016 12220
rect 127952 12180 127958 12192
rect 130010 12180 130016 12192
rect 130068 12180 130074 12232
rect 130102 12180 130108 12232
rect 130160 12220 130166 12232
rect 132126 12220 132132 12232
rect 130160 12192 132132 12220
rect 130160 12180 130166 12192
rect 132126 12180 132132 12192
rect 132184 12180 132190 12232
rect 133138 12180 133144 12232
rect 133196 12220 133202 12232
rect 134153 12223 134211 12229
rect 134153 12220 134165 12223
rect 133196 12192 134165 12220
rect 133196 12180 133202 12192
rect 134153 12189 134165 12192
rect 134199 12189 134211 12223
rect 134153 12183 134211 12189
rect 134420 12223 134478 12229
rect 134420 12189 134432 12223
rect 134466 12220 134478 12223
rect 135898 12220 135904 12232
rect 134466 12192 135904 12220
rect 134466 12189 134478 12192
rect 134420 12183 134478 12189
rect 135898 12180 135904 12192
rect 135956 12220 135962 12232
rect 136008 12220 136036 12260
rect 137005 12257 137017 12260
rect 137051 12257 137063 12291
rect 141160 12288 141188 12396
rect 141326 12384 141332 12396
rect 141384 12384 141390 12436
rect 143166 12384 143172 12436
rect 143224 12424 143230 12436
rect 146941 12427 146999 12433
rect 146941 12424 146953 12427
rect 143224 12396 146953 12424
rect 143224 12384 143230 12396
rect 146941 12393 146953 12396
rect 146987 12393 146999 12427
rect 146941 12387 146999 12393
rect 147140 12396 148088 12424
rect 141878 12356 141884 12368
rect 141839 12328 141884 12356
rect 141878 12316 141884 12328
rect 141936 12316 141942 12368
rect 143258 12288 143264 12300
rect 141160 12260 143264 12288
rect 137005 12251 137063 12257
rect 143258 12248 143264 12260
rect 143316 12248 143322 12300
rect 135956 12192 136036 12220
rect 136545 12223 136603 12229
rect 135956 12180 135962 12192
rect 136545 12189 136557 12223
rect 136591 12220 136603 12223
rect 138014 12220 138020 12232
rect 136591 12192 138020 12220
rect 136591 12189 136603 12192
rect 136545 12183 136603 12189
rect 138014 12180 138020 12192
rect 138072 12220 138078 12232
rect 140498 12220 140504 12232
rect 138072 12192 138165 12220
rect 140459 12192 140504 12220
rect 138072 12180 138078 12192
rect 140498 12180 140504 12192
rect 140556 12180 140562 12232
rect 140590 12180 140596 12232
rect 140648 12220 140654 12232
rect 141145 12223 141203 12229
rect 141145 12220 141157 12223
rect 140648 12192 141157 12220
rect 140648 12180 140654 12192
rect 141145 12189 141157 12192
rect 141191 12189 141203 12223
rect 141145 12183 141203 12189
rect 141234 12180 141240 12232
rect 141292 12220 141298 12232
rect 144549 12223 144607 12229
rect 141292 12192 144408 12220
rect 141292 12180 141298 12192
rect 115348 12124 118694 12152
rect 120005 12155 120063 12161
rect 115348 12112 115354 12124
rect 120005 12121 120017 12155
rect 120051 12152 120063 12155
rect 123604 12155 123662 12161
rect 120051 12124 123524 12152
rect 120051 12121 120063 12124
rect 120005 12115 120063 12121
rect 111058 12084 111064 12096
rect 109006 12056 111064 12084
rect 108301 12047 108359 12053
rect 111058 12044 111064 12056
rect 111116 12044 111122 12096
rect 111245 12087 111303 12093
rect 111245 12053 111257 12087
rect 111291 12084 111303 12087
rect 111610 12084 111616 12096
rect 111291 12056 111616 12084
rect 111291 12053 111303 12056
rect 111245 12047 111303 12053
rect 111610 12044 111616 12056
rect 111668 12044 111674 12096
rect 113542 12084 113548 12096
rect 113503 12056 113548 12084
rect 113542 12044 113548 12056
rect 113600 12044 113606 12096
rect 114097 12087 114155 12093
rect 114097 12053 114109 12087
rect 114143 12084 114155 12087
rect 114278 12084 114284 12096
rect 114143 12056 114284 12084
rect 114143 12053 114155 12056
rect 114097 12047 114155 12053
rect 114278 12044 114284 12056
rect 114336 12044 114342 12096
rect 114554 12084 114560 12096
rect 114515 12056 114560 12084
rect 114554 12044 114560 12056
rect 114612 12044 114618 12096
rect 115198 12084 115204 12096
rect 115159 12056 115204 12084
rect 115198 12044 115204 12056
rect 115256 12044 115262 12096
rect 116302 12084 116308 12096
rect 116263 12056 116308 12084
rect 116302 12044 116308 12056
rect 116360 12044 116366 12096
rect 116394 12044 116400 12096
rect 116452 12084 116458 12096
rect 117317 12087 117375 12093
rect 117317 12084 117329 12087
rect 116452 12056 117329 12084
rect 116452 12044 116458 12056
rect 117317 12053 117329 12056
rect 117363 12053 117375 12087
rect 118878 12084 118884 12096
rect 118791 12056 118884 12084
rect 117317 12047 117375 12053
rect 118878 12044 118884 12056
rect 118936 12084 118942 12096
rect 119890 12084 119896 12096
rect 118936 12056 119896 12084
rect 118936 12044 118942 12056
rect 119890 12044 119896 12056
rect 119948 12044 119954 12096
rect 120810 12084 120816 12096
rect 120771 12056 120816 12084
rect 120810 12044 120816 12056
rect 120868 12044 120874 12096
rect 123496 12084 123524 12124
rect 123604 12121 123616 12155
rect 123650 12152 123662 12155
rect 123754 12152 123760 12164
rect 123650 12124 123760 12152
rect 123650 12121 123662 12124
rect 123604 12115 123662 12121
rect 123754 12112 123760 12124
rect 123812 12112 123818 12164
rect 124140 12124 133460 12152
rect 124140 12084 124168 12124
rect 123496 12056 124168 12084
rect 124306 12044 124312 12096
rect 124364 12084 124370 12096
rect 124401 12087 124459 12093
rect 124401 12084 124413 12087
rect 124364 12056 124413 12084
rect 124364 12044 124370 12056
rect 124401 12053 124413 12056
rect 124447 12053 124459 12087
rect 124401 12047 124459 12053
rect 124858 12044 124864 12096
rect 124916 12084 124922 12096
rect 125045 12087 125103 12093
rect 125045 12084 125057 12087
rect 124916 12056 125057 12084
rect 124916 12044 124922 12056
rect 125045 12053 125057 12056
rect 125091 12053 125103 12087
rect 125045 12047 125103 12053
rect 126241 12087 126299 12093
rect 126241 12053 126253 12087
rect 126287 12084 126299 12087
rect 126330 12084 126336 12096
rect 126287 12056 126336 12084
rect 126287 12053 126299 12056
rect 126241 12047 126299 12053
rect 126330 12044 126336 12056
rect 126388 12044 126394 12096
rect 126698 12044 126704 12096
rect 126756 12084 126762 12096
rect 126793 12087 126851 12093
rect 126793 12084 126805 12087
rect 126756 12056 126805 12084
rect 126756 12044 126762 12056
rect 126793 12053 126805 12056
rect 126839 12084 126851 12087
rect 126882 12084 126888 12096
rect 126839 12056 126888 12084
rect 126839 12053 126851 12056
rect 126793 12047 126851 12053
rect 126882 12044 126888 12056
rect 126940 12044 126946 12096
rect 126974 12044 126980 12096
rect 127032 12084 127038 12096
rect 129461 12087 129519 12093
rect 129461 12084 129473 12087
rect 127032 12056 129473 12084
rect 127032 12044 127038 12056
rect 129461 12053 129473 12056
rect 129507 12053 129519 12087
rect 130654 12084 130660 12096
rect 130615 12056 130660 12084
rect 129461 12047 129519 12053
rect 130654 12044 130660 12056
rect 130712 12044 130718 12096
rect 131206 12084 131212 12096
rect 131167 12056 131212 12084
rect 131206 12044 131212 12056
rect 131264 12044 131270 12096
rect 131758 12084 131764 12096
rect 131719 12056 131764 12084
rect 131758 12044 131764 12056
rect 131816 12044 131822 12096
rect 132402 12044 132408 12096
rect 132460 12084 132466 12096
rect 133322 12084 133328 12096
rect 132460 12056 133328 12084
rect 132460 12044 132466 12056
rect 133322 12044 133328 12056
rect 133380 12044 133386 12096
rect 133432 12084 133460 12124
rect 135346 12112 135352 12164
rect 135404 12152 135410 12164
rect 140256 12155 140314 12161
rect 135404 12124 139164 12152
rect 135404 12112 135410 12124
rect 139136 12096 139164 12124
rect 140256 12121 140268 12155
rect 140302 12152 140314 12155
rect 141418 12152 141424 12164
rect 140302 12124 141424 12152
rect 140302 12121 140314 12124
rect 140256 12115 140314 12121
rect 141418 12112 141424 12124
rect 141476 12112 141482 12164
rect 141878 12112 141884 12164
rect 141936 12152 141942 12164
rect 142065 12155 142123 12161
rect 142065 12152 142077 12155
rect 141936 12124 142077 12152
rect 141936 12112 141942 12124
rect 142065 12121 142077 12124
rect 142111 12121 142123 12155
rect 144270 12152 144276 12164
rect 144328 12161 144334 12164
rect 144240 12124 144276 12152
rect 142065 12115 142123 12121
rect 144270 12112 144276 12124
rect 144328 12115 144340 12161
rect 144380 12152 144408 12192
rect 144549 12189 144561 12223
rect 144595 12220 144607 12223
rect 144730 12220 144736 12232
rect 144595 12192 144736 12220
rect 144595 12189 144607 12192
rect 144549 12183 144607 12189
rect 144730 12180 144736 12192
rect 144788 12180 144794 12232
rect 144822 12180 144828 12232
rect 144880 12220 144886 12232
rect 146386 12220 146392 12232
rect 144880 12192 146248 12220
rect 146347 12192 146392 12220
rect 144880 12180 144886 12192
rect 146110 12152 146116 12164
rect 146168 12161 146174 12164
rect 144380 12124 145972 12152
rect 146080 12124 146116 12152
rect 144328 12112 144334 12115
rect 136361 12087 136419 12093
rect 136361 12084 136373 12087
rect 133432 12056 136373 12084
rect 136361 12053 136373 12056
rect 136407 12053 136419 12087
rect 136361 12047 136419 12053
rect 138106 12044 138112 12096
rect 138164 12084 138170 12096
rect 138477 12087 138535 12093
rect 138477 12084 138489 12087
rect 138164 12056 138489 12084
rect 138164 12044 138170 12056
rect 138477 12053 138489 12056
rect 138523 12053 138535 12087
rect 139118 12084 139124 12096
rect 139079 12056 139124 12084
rect 138477 12047 138535 12053
rect 139118 12044 139124 12056
rect 139176 12044 139182 12096
rect 140038 12044 140044 12096
rect 140096 12084 140102 12096
rect 142338 12084 142344 12096
rect 140096 12056 142344 12084
rect 140096 12044 140102 12056
rect 142338 12044 142344 12056
rect 142396 12044 142402 12096
rect 143166 12084 143172 12096
rect 143127 12056 143172 12084
rect 143166 12044 143172 12056
rect 143224 12044 143230 12096
rect 145006 12084 145012 12096
rect 144967 12056 145012 12084
rect 145006 12044 145012 12056
rect 145064 12044 145070 12096
rect 145944 12084 145972 12124
rect 146110 12112 146116 12124
rect 146168 12115 146180 12161
rect 146220 12152 146248 12192
rect 146386 12180 146392 12192
rect 146444 12180 146450 12232
rect 147140 12229 147168 12396
rect 148060 12356 148088 12396
rect 148134 12384 148140 12436
rect 148192 12424 148198 12436
rect 149977 12427 150035 12433
rect 149977 12424 149989 12427
rect 148192 12396 149989 12424
rect 148192 12384 148198 12396
rect 149977 12393 149989 12396
rect 150023 12393 150035 12427
rect 149977 12387 150035 12393
rect 150452 12396 151400 12424
rect 150452 12356 150480 12396
rect 148060 12328 150480 12356
rect 151372 12356 151400 12396
rect 153102 12384 153108 12436
rect 153160 12424 153166 12436
rect 153160 12396 156828 12424
rect 153160 12384 153166 12396
rect 153381 12359 153439 12365
rect 153381 12356 153393 12359
rect 151372 12328 153393 12356
rect 153381 12325 153393 12328
rect 153427 12325 153439 12359
rect 153381 12319 153439 12325
rect 154758 12316 154764 12368
rect 154816 12356 154822 12368
rect 156233 12359 156291 12365
rect 156233 12356 156245 12359
rect 154816 12328 156245 12356
rect 154816 12316 154822 12328
rect 156233 12325 156245 12328
rect 156279 12325 156291 12359
rect 156233 12319 156291 12325
rect 148410 12288 148416 12300
rect 147232 12260 148416 12288
rect 147125 12223 147183 12229
rect 147125 12189 147137 12223
rect 147171 12189 147183 12223
rect 147125 12183 147183 12189
rect 147232 12152 147260 12260
rect 148410 12248 148416 12260
rect 148468 12248 148474 12300
rect 155589 12291 155647 12297
rect 151280 12260 153700 12288
rect 148042 12220 148048 12232
rect 146220 12124 147260 12152
rect 147324 12192 148048 12220
rect 146168 12112 146174 12115
rect 147324 12084 147352 12192
rect 148042 12180 148048 12192
rect 148100 12180 148106 12232
rect 148226 12180 148232 12232
rect 148284 12220 148290 12232
rect 148505 12223 148563 12229
rect 148505 12220 148517 12223
rect 148284 12192 148517 12220
rect 148284 12180 148290 12192
rect 148505 12189 148517 12192
rect 148551 12189 148563 12223
rect 148505 12183 148563 12189
rect 148594 12180 148600 12232
rect 148652 12220 148658 12232
rect 148965 12223 149023 12229
rect 148965 12220 148977 12223
rect 148652 12192 148977 12220
rect 148652 12180 148658 12192
rect 148965 12189 148977 12192
rect 149011 12189 149023 12223
rect 148965 12183 149023 12189
rect 150250 12180 150256 12232
rect 150308 12220 150314 12232
rect 151280 12220 151308 12260
rect 150308 12192 151308 12220
rect 150308 12180 150314 12192
rect 151354 12180 151360 12232
rect 151412 12220 151418 12232
rect 152001 12223 152059 12229
rect 151412 12192 151457 12220
rect 151412 12180 151418 12192
rect 152001 12189 152013 12223
rect 152047 12189 152059 12223
rect 152642 12220 152648 12232
rect 152603 12192 152648 12220
rect 152001 12183 152059 12189
rect 147674 12112 147680 12164
rect 147732 12152 147738 12164
rect 150526 12152 150532 12164
rect 147732 12124 150532 12152
rect 147732 12112 147738 12124
rect 150526 12112 150532 12124
rect 150584 12112 150590 12164
rect 151078 12112 151084 12164
rect 151136 12161 151142 12164
rect 151136 12152 151148 12161
rect 152016 12152 152044 12183
rect 152642 12180 152648 12192
rect 152700 12180 152706 12232
rect 152829 12223 152887 12229
rect 152829 12189 152841 12223
rect 152875 12220 152887 12223
rect 153010 12220 153016 12232
rect 152875 12192 153016 12220
rect 152875 12189 152887 12192
rect 152829 12183 152887 12189
rect 153010 12180 153016 12192
rect 153068 12180 153074 12232
rect 153672 12220 153700 12260
rect 155589 12257 155601 12291
rect 155635 12288 155647 12291
rect 155862 12288 155868 12300
rect 155635 12260 155868 12288
rect 155635 12257 155647 12260
rect 155589 12251 155647 12257
rect 155862 12248 155868 12260
rect 155920 12248 155926 12300
rect 153672 12192 154620 12220
rect 151136 12124 151181 12152
rect 152016 12124 153516 12152
rect 151136 12115 151148 12124
rect 151136 12112 151142 12115
rect 147582 12084 147588 12096
rect 145944 12056 147352 12084
rect 147543 12056 147588 12084
rect 147582 12044 147588 12056
rect 147640 12044 147646 12096
rect 148318 12084 148324 12096
rect 148279 12056 148324 12084
rect 148318 12044 148324 12056
rect 148376 12044 148382 12096
rect 148410 12044 148416 12096
rect 148468 12084 148474 12096
rect 149149 12087 149207 12093
rect 149149 12084 149161 12087
rect 148468 12056 149161 12084
rect 148468 12044 148474 12056
rect 149149 12053 149161 12056
rect 149195 12053 149207 12087
rect 149149 12047 149207 12053
rect 149238 12044 149244 12096
rect 149296 12084 149302 12096
rect 151817 12087 151875 12093
rect 151817 12084 151829 12087
rect 149296 12056 151829 12084
rect 149296 12044 149302 12056
rect 151817 12053 151829 12056
rect 151863 12053 151875 12087
rect 151817 12047 151875 12053
rect 151906 12044 151912 12096
rect 151964 12084 151970 12096
rect 152461 12087 152519 12093
rect 152461 12084 152473 12087
rect 151964 12056 152473 12084
rect 151964 12044 151970 12056
rect 152461 12053 152473 12056
rect 152507 12053 152519 12087
rect 153488 12084 153516 12124
rect 153746 12112 153752 12164
rect 153804 12152 153810 12164
rect 154494 12155 154552 12161
rect 154494 12152 154506 12155
rect 153804 12124 154506 12152
rect 153804 12112 153810 12124
rect 154494 12121 154506 12124
rect 154540 12121 154552 12155
rect 154592 12152 154620 12192
rect 154666 12180 154672 12232
rect 154724 12220 154730 12232
rect 154761 12223 154819 12229
rect 154761 12220 154773 12223
rect 154724 12192 154773 12220
rect 154724 12180 154730 12192
rect 154761 12189 154773 12192
rect 154807 12189 154819 12223
rect 154761 12183 154819 12189
rect 155218 12180 155224 12232
rect 155276 12220 155282 12232
rect 155405 12223 155463 12229
rect 155405 12220 155417 12223
rect 155276 12192 155417 12220
rect 155276 12180 155282 12192
rect 155405 12189 155417 12192
rect 155451 12189 155463 12223
rect 155405 12183 155463 12189
rect 155494 12180 155500 12232
rect 155552 12220 155558 12232
rect 156800 12229 156828 12396
rect 156049 12223 156107 12229
rect 156049 12220 156061 12223
rect 155552 12192 156061 12220
rect 155552 12180 155558 12192
rect 156049 12189 156061 12192
rect 156095 12189 156107 12223
rect 156049 12183 156107 12189
rect 156785 12223 156843 12229
rect 156785 12189 156797 12223
rect 156831 12189 156843 12223
rect 156785 12183 156843 12189
rect 157705 12223 157763 12229
rect 157705 12189 157717 12223
rect 157751 12220 157763 12223
rect 159174 12220 159180 12232
rect 157751 12192 159180 12220
rect 157751 12189 157763 12192
rect 157705 12183 157763 12189
rect 159174 12180 159180 12192
rect 159232 12180 159238 12232
rect 154592 12124 157012 12152
rect 154494 12115 154552 12121
rect 156984 12093 157012 12124
rect 155221 12087 155279 12093
rect 155221 12084 155233 12087
rect 153488 12056 155233 12084
rect 152461 12047 152519 12053
rect 155221 12053 155233 12056
rect 155267 12053 155279 12087
rect 155221 12047 155279 12053
rect 156969 12087 157027 12093
rect 156969 12053 156981 12087
rect 157015 12053 157027 12087
rect 156969 12047 157027 12053
rect 157058 12044 157064 12096
rect 157116 12084 157122 12096
rect 157521 12087 157579 12093
rect 157521 12084 157533 12087
rect 157116 12056 157533 12084
rect 157116 12044 157122 12056
rect 157521 12053 157533 12056
rect 157567 12053 157579 12087
rect 157521 12047 157579 12053
rect 1104 11994 159043 12016
rect 1104 11942 40394 11994
rect 40446 11942 40458 11994
rect 40510 11942 40522 11994
rect 40574 11942 40586 11994
rect 40638 11942 40650 11994
rect 40702 11942 79839 11994
rect 79891 11942 79903 11994
rect 79955 11942 79967 11994
rect 80019 11942 80031 11994
rect 80083 11942 80095 11994
rect 80147 11942 119284 11994
rect 119336 11942 119348 11994
rect 119400 11942 119412 11994
rect 119464 11942 119476 11994
rect 119528 11942 119540 11994
rect 119592 11942 158729 11994
rect 158781 11942 158793 11994
rect 158845 11942 158857 11994
rect 158909 11942 158921 11994
rect 158973 11942 158985 11994
rect 159037 11942 159043 11994
rect 1104 11920 159043 11942
rect 10505 11883 10563 11889
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 13170 11880 13176 11892
rect 10551 11852 13176 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 14274 11880 14280 11892
rect 13464 11852 14280 11880
rect 13265 11815 13323 11821
rect 13265 11812 13277 11815
rect 10980 11784 13277 11812
rect 4062 11753 4068 11756
rect 4056 11707 4068 11753
rect 4120 11744 4126 11756
rect 8386 11744 8392 11756
rect 4120 11716 4156 11744
rect 8347 11716 8392 11744
rect 4062 11704 4068 11707
rect 4120 11704 4126 11716
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 10980 11753 11008 11784
rect 13265 11781 13277 11784
rect 13311 11781 13323 11815
rect 13265 11775 13323 11781
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11882 11744 11888 11756
rect 11296 11716 11888 11744
rect 11296 11704 11302 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12526 11744 12532 11756
rect 12268 11716 12532 11744
rect 3786 11676 3792 11688
rect 3747 11648 3792 11676
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 12268 11676 12296 11716
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 13354 11744 13360 11756
rect 12851 11716 13360 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13464 11753 13492 11852
rect 14274 11840 14280 11852
rect 14332 11880 14338 11892
rect 18509 11883 18567 11889
rect 14332 11852 17540 11880
rect 14332 11840 14338 11852
rect 14918 11772 14924 11824
rect 14976 11812 14982 11824
rect 15562 11812 15568 11824
rect 14976 11784 15568 11812
rect 14976 11772 14982 11784
rect 15562 11772 15568 11784
rect 15620 11812 15626 11824
rect 17374 11815 17432 11821
rect 17374 11812 17386 11815
rect 15620 11784 17386 11812
rect 15620 11772 15626 11784
rect 17374 11781 17386 11784
rect 17420 11781 17432 11815
rect 17374 11775 17432 11781
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 13449 11707 13507 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14717 11747 14775 11753
rect 14717 11744 14729 11747
rect 14608 11716 14729 11744
rect 14608 11704 14614 11716
rect 14717 11713 14729 11716
rect 14763 11713 14775 11747
rect 14717 11707 14775 11713
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15470 11744 15476 11756
rect 15252 11716 15476 11744
rect 15252 11704 15258 11716
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 17218 11744 17224 11756
rect 16172 11716 17224 11744
rect 16172 11704 16178 11716
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17512 11744 17540 11852
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 20162 11880 20168 11892
rect 18555 11852 20168 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20588 11852 20821 11880
rect 20588 11840 20594 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 23937 11883 23995 11889
rect 23937 11880 23949 11883
rect 21692 11852 23949 11880
rect 21692 11840 21698 11852
rect 23937 11849 23949 11852
rect 23983 11849 23995 11883
rect 23937 11843 23995 11849
rect 26237 11883 26295 11889
rect 26237 11849 26249 11883
rect 26283 11880 26295 11883
rect 27614 11880 27620 11892
rect 26283 11852 27620 11880
rect 26283 11849 26295 11852
rect 26237 11843 26295 11849
rect 27614 11840 27620 11852
rect 27672 11840 27678 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 31021 11883 31079 11889
rect 31021 11880 31033 11883
rect 28040 11852 31033 11880
rect 28040 11840 28046 11852
rect 31021 11849 31033 11852
rect 31067 11849 31079 11883
rect 31021 11843 31079 11849
rect 31110 11840 31116 11892
rect 31168 11880 31174 11892
rect 31665 11883 31723 11889
rect 31665 11880 31677 11883
rect 31168 11852 31677 11880
rect 31168 11840 31174 11852
rect 31665 11849 31677 11852
rect 31711 11849 31723 11883
rect 31665 11843 31723 11849
rect 32306 11840 32312 11892
rect 32364 11880 32370 11892
rect 32858 11880 32864 11892
rect 32364 11852 32864 11880
rect 32364 11840 32370 11852
rect 32858 11840 32864 11852
rect 32916 11840 32922 11892
rect 36354 11880 36360 11892
rect 36315 11852 36360 11880
rect 36354 11840 36360 11852
rect 36412 11840 36418 11892
rect 37642 11840 37648 11892
rect 37700 11880 37706 11892
rect 39298 11880 39304 11892
rect 37700 11852 39304 11880
rect 37700 11840 37706 11852
rect 39298 11840 39304 11852
rect 39356 11840 39362 11892
rect 39482 11840 39488 11892
rect 39540 11880 39546 11892
rect 39669 11883 39727 11889
rect 39669 11880 39681 11883
rect 39540 11852 39681 11880
rect 39540 11840 39546 11852
rect 39669 11849 39681 11852
rect 39715 11849 39727 11883
rect 39669 11843 39727 11849
rect 40218 11840 40224 11892
rect 40276 11880 40282 11892
rect 41690 11880 41696 11892
rect 40276 11852 41696 11880
rect 40276 11840 40282 11852
rect 41690 11840 41696 11852
rect 41748 11840 41754 11892
rect 41877 11883 41935 11889
rect 41877 11849 41889 11883
rect 41923 11880 41935 11883
rect 43254 11880 43260 11892
rect 41923 11852 43260 11880
rect 41923 11849 41935 11852
rect 41877 11843 41935 11849
rect 43254 11840 43260 11852
rect 43312 11840 43318 11892
rect 44361 11883 44419 11889
rect 44361 11849 44373 11883
rect 44407 11849 44419 11883
rect 44361 11843 44419 11849
rect 45097 11883 45155 11889
rect 45097 11849 45109 11883
rect 45143 11880 45155 11883
rect 45143 11852 46704 11880
rect 45143 11849 45155 11852
rect 45097 11843 45155 11849
rect 19153 11815 19211 11821
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 19794 11812 19800 11824
rect 19199 11784 19800 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 21910 11812 21916 11824
rect 19904 11784 21916 11812
rect 19904 11744 19932 11784
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 25102 11815 25160 11821
rect 25102 11812 25114 11815
rect 22066 11784 25114 11812
rect 17512 11716 19932 11744
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 12618 11676 12624 11688
rect 8573 11639 8631 11645
rect 11164 11648 12296 11676
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 6144 11580 8217 11608
rect 6144 11568 6150 11580
rect 8205 11577 8217 11580
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5534 11540 5540 11552
rect 5215 11512 5540 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 7742 11540 7748 11552
rect 7703 11512 7748 11540
rect 7742 11500 7748 11512
rect 7800 11540 7806 11552
rect 8588 11540 8616 11639
rect 9401 11611 9459 11617
rect 9401 11577 9413 11611
rect 9447 11608 9459 11611
rect 10318 11608 10324 11620
rect 9447 11580 10324 11608
rect 9447 11577 9459 11580
rect 9401 11571 9459 11577
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 11164 11617 11192 11648
rect 12605 11636 12624 11676
rect 12676 11636 12682 11688
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 12952 11648 13645 11676
rect 12952 11636 12958 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 17092 11648 17141 11676
rect 17092 11636 17098 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 19242 11676 19248 11688
rect 18196 11648 19248 11676
rect 18196 11636 18202 11648
rect 19242 11636 19248 11648
rect 19300 11676 19306 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19300 11648 19625 11676
rect 19300 11636 19306 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 21008 11676 21036 11707
rect 21082 11704 21088 11756
rect 21140 11744 21146 11756
rect 22066 11744 22094 11784
rect 25102 11781 25114 11784
rect 25148 11781 25160 11815
rect 25102 11775 25160 11781
rect 28068 11815 28126 11821
rect 28068 11781 28080 11815
rect 28114 11812 28126 11815
rect 29178 11812 29184 11824
rect 28114 11784 29184 11812
rect 28114 11781 28126 11784
rect 28068 11775 28126 11781
rect 29178 11772 29184 11784
rect 29236 11772 29242 11824
rect 29546 11772 29552 11824
rect 29604 11812 29610 11824
rect 30466 11812 30472 11824
rect 29604 11784 30472 11812
rect 29604 11772 29610 11784
rect 30466 11772 30472 11784
rect 30524 11772 30530 11824
rect 35894 11772 35900 11824
rect 35952 11812 35958 11824
rect 40034 11812 40040 11824
rect 35952 11784 40040 11812
rect 35952 11772 35958 11784
rect 40034 11772 40040 11784
rect 40092 11812 40098 11824
rect 43622 11812 43628 11824
rect 40092 11784 40724 11812
rect 40092 11772 40098 11784
rect 21140 11716 22094 11744
rect 21140 11704 21146 11716
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22244 11716 22937 11744
rect 22244 11704 22250 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 24118 11744 24124 11756
rect 22925 11707 22983 11713
rect 23032 11716 23704 11744
rect 24079 11716 24124 11744
rect 23032 11676 23060 11716
rect 21008 11648 23060 11676
rect 23109 11679 23167 11685
rect 19613 11639 19671 11645
rect 23109 11645 23121 11679
rect 23155 11645 23167 11679
rect 23109 11639 23167 11645
rect 11149 11611 11207 11617
rect 11149 11577 11161 11611
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 7800 11512 8616 11540
rect 9953 11543 10011 11549
rect 7800 11500 7806 11512
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10042 11540 10048 11552
rect 9999 11512 10048 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 12066 11540 12072 11552
rect 12027 11512 12072 11540
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12605 11549 12633 11636
rect 18598 11568 18604 11620
rect 18656 11608 18662 11620
rect 22741 11611 22799 11617
rect 22741 11608 22753 11611
rect 18656 11580 22753 11608
rect 18656 11568 18662 11580
rect 22741 11577 22753 11580
rect 22787 11577 22799 11611
rect 23124 11608 23152 11639
rect 22741 11571 22799 11577
rect 22940 11580 23152 11608
rect 12605 11543 12679 11549
rect 12605 11512 12633 11543
rect 12621 11509 12633 11512
rect 12667 11509 12679 11543
rect 15838 11540 15844 11552
rect 15799 11512 15844 11540
rect 12621 11503 12679 11509
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 19334 11540 19340 11552
rect 15988 11512 19340 11540
rect 15988 11500 15994 11512
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 20162 11540 20168 11552
rect 20123 11512 20168 11540
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 22094 11540 22100 11552
rect 20312 11512 22100 11540
rect 20312 11500 20318 11512
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22940 11540 22968 11580
rect 22336 11512 22968 11540
rect 23676 11540 23704 11716
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11744 24915 11747
rect 24946 11744 24952 11756
rect 24903 11716 24952 11744
rect 24903 11713 24915 11716
rect 24857 11707 24915 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 27706 11744 27712 11756
rect 27387 11716 27712 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 27706 11704 27712 11716
rect 27764 11744 27770 11756
rect 28810 11744 28816 11756
rect 27764 11716 28816 11744
rect 27764 11704 27770 11716
rect 28810 11704 28816 11716
rect 28868 11704 28874 11756
rect 29897 11747 29955 11753
rect 29897 11744 29909 11747
rect 28920 11716 29909 11744
rect 23750 11636 23756 11688
rect 23808 11676 23814 11688
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 23808 11648 24317 11676
rect 23808 11636 23814 11648
rect 24305 11645 24317 11648
rect 24351 11645 24363 11679
rect 24305 11639 24363 11645
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 26602 11676 26608 11688
rect 26292 11648 26608 11676
rect 26292 11636 26298 11648
rect 26602 11636 26608 11648
rect 26660 11676 26666 11688
rect 27801 11679 27859 11685
rect 27801 11676 27813 11679
rect 26660 11648 27813 11676
rect 26660 11636 26666 11648
rect 27801 11645 27813 11648
rect 27847 11645 27859 11679
rect 27801 11639 27859 11645
rect 25958 11568 25964 11620
rect 26016 11608 26022 11620
rect 26016 11580 27200 11608
rect 26016 11568 26022 11580
rect 27062 11540 27068 11552
rect 23676 11512 27068 11540
rect 22336 11500 22342 11512
rect 27062 11500 27068 11512
rect 27120 11500 27126 11552
rect 27172 11540 27200 11580
rect 28920 11540 28948 11716
rect 29897 11713 29909 11716
rect 29943 11713 29955 11747
rect 29897 11707 29955 11713
rect 30190 11704 30196 11756
rect 30248 11744 30254 11756
rect 31481 11747 31539 11753
rect 31481 11744 31493 11747
rect 30248 11716 31493 11744
rect 30248 11704 30254 11716
rect 31481 11713 31493 11716
rect 31527 11713 31539 11747
rect 31481 11707 31539 11713
rect 31662 11704 31668 11756
rect 31720 11744 31726 11756
rect 32030 11744 32036 11756
rect 31720 11716 32036 11744
rect 31720 11704 31726 11716
rect 32030 11704 32036 11716
rect 32088 11744 32094 11756
rect 34054 11744 34060 11756
rect 32088 11716 34060 11744
rect 32088 11704 32094 11716
rect 34054 11704 34060 11716
rect 34112 11704 34118 11756
rect 38545 11747 38603 11753
rect 38545 11744 38557 11747
rect 35176 11716 38557 11744
rect 28994 11636 29000 11688
rect 29052 11676 29058 11688
rect 29638 11676 29644 11688
rect 29052 11648 29644 11676
rect 29052 11636 29058 11648
rect 29638 11636 29644 11648
rect 29696 11636 29702 11688
rect 30834 11636 30840 11688
rect 30892 11676 30898 11688
rect 35176 11676 35204 11716
rect 38545 11713 38557 11716
rect 38591 11713 38603 11747
rect 38545 11707 38603 11713
rect 39114 11704 39120 11756
rect 39172 11744 39178 11756
rect 40696 11753 40724 11784
rect 42076 11784 43628 11812
rect 40497 11747 40555 11753
rect 40497 11744 40509 11747
rect 39172 11716 40509 11744
rect 39172 11704 39178 11716
rect 40497 11713 40509 11716
rect 40543 11713 40555 11747
rect 40497 11707 40555 11713
rect 40681 11747 40739 11753
rect 40681 11713 40693 11747
rect 40727 11713 40739 11747
rect 40681 11707 40739 11713
rect 41506 11704 41512 11756
rect 41564 11744 41570 11756
rect 41966 11744 41972 11756
rect 41564 11716 41972 11744
rect 41564 11704 41570 11716
rect 41966 11704 41972 11716
rect 42024 11704 42030 11756
rect 42076 11753 42104 11784
rect 43622 11772 43628 11784
rect 43680 11772 43686 11824
rect 43898 11772 43904 11824
rect 43956 11812 43962 11824
rect 44376 11812 44404 11843
rect 45916 11815 45974 11821
rect 43956 11784 44312 11812
rect 44376 11784 45876 11812
rect 43956 11772 43962 11784
rect 42061 11747 42119 11753
rect 42061 11713 42073 11747
rect 42107 11713 42119 11747
rect 42061 11707 42119 11713
rect 42150 11704 42156 11756
rect 42208 11744 42214 11756
rect 42705 11747 42763 11753
rect 42705 11744 42717 11747
rect 42208 11716 42717 11744
rect 42208 11704 42214 11716
rect 42705 11713 42717 11716
rect 42751 11713 42763 11747
rect 42705 11707 42763 11713
rect 42794 11704 42800 11756
rect 42852 11744 42858 11756
rect 43441 11747 43499 11753
rect 43441 11744 43453 11747
rect 42852 11716 43453 11744
rect 42852 11704 42858 11716
rect 43441 11713 43453 11716
rect 43487 11713 43499 11747
rect 44174 11744 44180 11756
rect 44135 11716 44180 11744
rect 43441 11707 43499 11713
rect 44174 11704 44180 11716
rect 44232 11704 44238 11756
rect 44284 11744 44312 11784
rect 44913 11747 44971 11753
rect 44913 11744 44925 11747
rect 44284 11716 44925 11744
rect 44913 11713 44925 11716
rect 44959 11713 44971 11747
rect 45646 11744 45652 11756
rect 45607 11716 45652 11744
rect 44913 11707 44971 11713
rect 45646 11704 45652 11716
rect 45704 11704 45710 11756
rect 45848 11744 45876 11784
rect 45916 11781 45928 11815
rect 45962 11812 45974 11815
rect 46382 11812 46388 11824
rect 45962 11784 46388 11812
rect 45962 11781 45974 11784
rect 45916 11775 45974 11781
rect 46382 11772 46388 11784
rect 46440 11772 46446 11824
rect 46676 11812 46704 11852
rect 46934 11840 46940 11892
rect 46992 11880 46998 11892
rect 47029 11883 47087 11889
rect 47029 11880 47041 11883
rect 46992 11852 47041 11880
rect 46992 11840 46998 11852
rect 47029 11849 47041 11852
rect 47075 11880 47087 11883
rect 48130 11880 48136 11892
rect 47075 11852 48136 11880
rect 47075 11849 47087 11852
rect 47029 11843 47087 11849
rect 48130 11840 48136 11852
rect 48188 11840 48194 11892
rect 48409 11883 48467 11889
rect 48409 11849 48421 11883
rect 48455 11880 48467 11883
rect 50982 11880 50988 11892
rect 48455 11852 50988 11880
rect 48455 11849 48467 11852
rect 48409 11843 48467 11849
rect 50982 11840 50988 11852
rect 51040 11840 51046 11892
rect 52089 11883 52147 11889
rect 51828 11852 52040 11880
rect 48222 11812 48228 11824
rect 46676 11784 48228 11812
rect 48222 11772 48228 11784
rect 48280 11772 48286 11824
rect 49510 11772 49516 11824
rect 49568 11812 49574 11824
rect 51828 11812 51856 11852
rect 49568 11784 51856 11812
rect 52012 11812 52040 11852
rect 52089 11849 52101 11883
rect 52135 11880 52147 11883
rect 52362 11880 52368 11892
rect 52135 11852 52368 11880
rect 52135 11849 52147 11852
rect 52089 11843 52147 11849
rect 52362 11840 52368 11852
rect 52420 11840 52426 11892
rect 52822 11840 52828 11892
rect 52880 11880 52886 11892
rect 52917 11883 52975 11889
rect 52917 11880 52929 11883
rect 52880 11852 52929 11880
rect 52880 11840 52886 11852
rect 52917 11849 52929 11852
rect 52963 11849 52975 11883
rect 52917 11843 52975 11849
rect 53745 11883 53803 11889
rect 53745 11849 53757 11883
rect 53791 11849 53803 11883
rect 54294 11880 54300 11892
rect 54255 11852 54300 11880
rect 53745 11843 53803 11849
rect 53760 11812 53788 11843
rect 54294 11840 54300 11852
rect 54352 11840 54358 11892
rect 54386 11840 54392 11892
rect 54444 11880 54450 11892
rect 56042 11880 56048 11892
rect 54444 11852 56048 11880
rect 54444 11840 54450 11852
rect 56042 11840 56048 11852
rect 56100 11840 56106 11892
rect 57238 11880 57244 11892
rect 56336 11852 57244 11880
rect 55214 11812 55220 11824
rect 52012 11784 53696 11812
rect 53760 11784 55220 11812
rect 49568 11772 49574 11784
rect 47670 11744 47676 11756
rect 45848 11716 47676 11744
rect 47670 11704 47676 11716
rect 47728 11704 47734 11756
rect 48593 11747 48651 11753
rect 48593 11713 48605 11747
rect 48639 11744 48651 11747
rect 49142 11744 49148 11756
rect 48639 11716 49148 11744
rect 48639 11713 48651 11716
rect 48593 11707 48651 11713
rect 49142 11704 49148 11716
rect 49200 11704 49206 11756
rect 49326 11744 49332 11756
rect 49287 11716 49332 11744
rect 49326 11704 49332 11716
rect 49384 11704 49390 11756
rect 50062 11753 50068 11756
rect 50056 11707 50068 11753
rect 50120 11744 50126 11756
rect 51902 11744 51908 11756
rect 50120 11716 50156 11744
rect 51863 11716 51908 11744
rect 50062 11704 50068 11707
rect 50120 11704 50126 11716
rect 51902 11704 51908 11716
rect 51960 11704 51966 11756
rect 52454 11704 52460 11756
rect 52512 11744 52518 11756
rect 53101 11747 53159 11753
rect 53101 11744 53113 11747
rect 52512 11716 53113 11744
rect 52512 11704 52518 11716
rect 53101 11713 53113 11716
rect 53147 11713 53159 11747
rect 53558 11744 53564 11756
rect 53519 11716 53564 11744
rect 53101 11707 53159 11713
rect 53558 11704 53564 11716
rect 53616 11704 53622 11756
rect 53668 11744 53696 11784
rect 55214 11772 55220 11784
rect 55272 11772 55278 11824
rect 55306 11772 55312 11824
rect 55364 11812 55370 11824
rect 56336 11812 56364 11852
rect 57238 11840 57244 11852
rect 57296 11880 57302 11892
rect 58618 11880 58624 11892
rect 57296 11852 58624 11880
rect 57296 11840 57302 11852
rect 58618 11840 58624 11852
rect 58676 11880 58682 11892
rect 59078 11880 59084 11892
rect 58676 11852 59084 11880
rect 58676 11840 58682 11852
rect 59078 11840 59084 11852
rect 59136 11840 59142 11892
rect 59446 11880 59452 11892
rect 59407 11852 59452 11880
rect 59446 11840 59452 11852
rect 59504 11840 59510 11892
rect 59740 11852 59952 11880
rect 56410 11821 56416 11824
rect 55364 11784 56364 11812
rect 56393 11815 56416 11821
rect 55364 11772 55370 11784
rect 56393 11781 56405 11815
rect 56393 11775 56416 11781
rect 56410 11772 56416 11775
rect 56468 11772 56474 11824
rect 59740 11812 59768 11852
rect 58176 11784 59768 11812
rect 55410 11747 55468 11753
rect 55410 11744 55422 11747
rect 53668 11716 55422 11744
rect 55410 11713 55422 11716
rect 55456 11744 55468 11747
rect 57330 11744 57336 11756
rect 55456 11716 57336 11744
rect 55456 11713 55468 11716
rect 55410 11707 55468 11713
rect 57330 11704 57336 11716
rect 57388 11704 57394 11756
rect 57882 11704 57888 11756
rect 57940 11744 57946 11756
rect 58069 11747 58127 11753
rect 58069 11744 58081 11747
rect 57940 11716 58081 11744
rect 57940 11704 57946 11716
rect 58069 11713 58081 11716
rect 58115 11713 58127 11747
rect 58069 11707 58127 11713
rect 30892 11648 35204 11676
rect 30892 11636 30898 11648
rect 37182 11636 37188 11688
rect 37240 11676 37246 11688
rect 38289 11679 38347 11685
rect 38289 11676 38301 11679
rect 37240 11648 38301 11676
rect 37240 11636 37246 11648
rect 38289 11645 38301 11648
rect 38335 11645 38347 11679
rect 38289 11639 38347 11645
rect 40865 11679 40923 11685
rect 40865 11645 40877 11679
rect 40911 11676 40923 11679
rect 42610 11676 42616 11688
rect 40911 11648 42616 11676
rect 40911 11645 40923 11648
rect 40865 11639 40923 11645
rect 42610 11636 42616 11648
rect 42668 11636 42674 11688
rect 44358 11676 44364 11688
rect 42996 11648 44364 11676
rect 30650 11568 30656 11620
rect 30708 11608 30714 11620
rect 34790 11608 34796 11620
rect 30708 11580 34652 11608
rect 34751 11580 34796 11608
rect 30708 11568 30714 11580
rect 27172 11512 28948 11540
rect 29181 11543 29239 11549
rect 29181 11509 29193 11543
rect 29227 11540 29239 11543
rect 30742 11540 30748 11552
rect 29227 11512 30748 11540
rect 29227 11509 29239 11512
rect 29181 11503 29239 11509
rect 30742 11500 30748 11512
rect 30800 11500 30806 11552
rect 31754 11500 31760 11552
rect 31812 11540 31818 11552
rect 32309 11543 32367 11549
rect 32309 11540 32321 11543
rect 31812 11512 32321 11540
rect 31812 11500 31818 11512
rect 32309 11509 32321 11512
rect 32355 11509 32367 11543
rect 32309 11503 32367 11509
rect 33597 11543 33655 11549
rect 33597 11509 33609 11543
rect 33643 11540 33655 11543
rect 33870 11540 33876 11552
rect 33643 11512 33876 11540
rect 33643 11509 33655 11512
rect 33597 11503 33655 11509
rect 33870 11500 33876 11512
rect 33928 11500 33934 11552
rect 34238 11540 34244 11552
rect 34199 11512 34244 11540
rect 34238 11500 34244 11512
rect 34296 11500 34302 11552
rect 34624 11540 34652 11580
rect 34790 11568 34796 11580
rect 34848 11568 34854 11620
rect 36909 11611 36967 11617
rect 36909 11577 36921 11611
rect 36955 11608 36967 11611
rect 36955 11580 38332 11608
rect 36955 11577 36967 11580
rect 36909 11571 36967 11577
rect 36538 11540 36544 11552
rect 34624 11512 36544 11540
rect 36538 11500 36544 11512
rect 36596 11500 36602 11552
rect 37826 11540 37832 11552
rect 37787 11512 37832 11540
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 38304 11540 38332 11580
rect 39298 11568 39304 11620
rect 39356 11608 39362 11620
rect 41322 11608 41328 11620
rect 39356 11580 41328 11608
rect 39356 11568 39362 11580
rect 41322 11568 41328 11580
rect 41380 11568 41386 11620
rect 39206 11540 39212 11552
rect 38304 11512 39212 11540
rect 39206 11500 39212 11512
rect 39264 11540 39270 11552
rect 42426 11540 42432 11552
rect 39264 11512 42432 11540
rect 39264 11500 39270 11512
rect 42426 11500 42432 11512
rect 42484 11500 42490 11552
rect 42889 11543 42947 11549
rect 42889 11509 42901 11543
rect 42935 11540 42947 11543
rect 42996 11540 43024 11648
rect 44358 11636 44364 11648
rect 44416 11636 44422 11688
rect 46658 11636 46664 11688
rect 46716 11676 46722 11688
rect 49234 11676 49240 11688
rect 46716 11648 49240 11676
rect 46716 11636 46722 11648
rect 49234 11636 49240 11648
rect 49292 11636 49298 11688
rect 49786 11676 49792 11688
rect 49747 11648 49792 11676
rect 49786 11636 49792 11648
rect 49844 11636 49850 11688
rect 51074 11636 51080 11688
rect 51132 11676 51138 11688
rect 51534 11676 51540 11688
rect 51132 11648 51540 11676
rect 51132 11636 51138 11648
rect 51534 11636 51540 11648
rect 51592 11676 51598 11688
rect 51721 11679 51779 11685
rect 51721 11676 51733 11679
rect 51592 11648 51733 11676
rect 51592 11636 51598 11648
rect 51721 11645 51733 11648
rect 51767 11645 51779 11679
rect 51721 11639 51779 11645
rect 52086 11636 52092 11688
rect 52144 11636 52150 11688
rect 53006 11636 53012 11688
rect 53064 11676 53070 11688
rect 54018 11676 54024 11688
rect 53064 11648 54024 11676
rect 53064 11636 53070 11648
rect 54018 11636 54024 11648
rect 54076 11636 54082 11688
rect 55677 11679 55735 11685
rect 55677 11645 55689 11679
rect 55723 11676 55735 11679
rect 55766 11676 55772 11688
rect 55723 11648 55772 11676
rect 55723 11645 55735 11648
rect 55677 11639 55735 11645
rect 55766 11636 55772 11648
rect 55824 11636 55830 11688
rect 56134 11676 56140 11688
rect 56095 11648 56140 11676
rect 56134 11636 56140 11648
rect 56192 11636 56198 11688
rect 58176 11676 58204 11784
rect 58336 11747 58394 11753
rect 58336 11713 58348 11747
rect 58382 11744 58394 11747
rect 59538 11744 59544 11756
rect 58382 11716 59544 11744
rect 58382 11713 58394 11716
rect 58336 11707 58394 11713
rect 59538 11704 59544 11716
rect 59596 11704 59602 11756
rect 59924 11744 59952 11852
rect 59998 11840 60004 11892
rect 60056 11880 60062 11892
rect 60918 11880 60924 11892
rect 60056 11852 60924 11880
rect 60056 11840 60062 11852
rect 60918 11840 60924 11852
rect 60976 11840 60982 11892
rect 61010 11840 61016 11892
rect 61068 11880 61074 11892
rect 61286 11880 61292 11892
rect 61068 11852 61292 11880
rect 61068 11840 61074 11852
rect 61286 11840 61292 11852
rect 61344 11880 61350 11892
rect 62298 11880 62304 11892
rect 61344 11852 62304 11880
rect 61344 11840 61350 11852
rect 62298 11840 62304 11852
rect 62356 11840 62362 11892
rect 62574 11840 62580 11892
rect 62632 11880 62638 11892
rect 63405 11883 63463 11889
rect 63405 11880 63417 11883
rect 62632 11852 63417 11880
rect 62632 11840 62638 11852
rect 63405 11849 63417 11852
rect 63451 11849 63463 11883
rect 70946 11880 70952 11892
rect 63405 11843 63463 11849
rect 68296 11852 70952 11880
rect 60090 11772 60096 11824
rect 60148 11812 60154 11824
rect 67174 11812 67180 11824
rect 60148 11784 64000 11812
rect 60148 11772 60154 11784
rect 60642 11744 60648 11756
rect 59924 11716 60648 11744
rect 60642 11704 60648 11716
rect 60700 11704 60706 11756
rect 61562 11753 61568 11756
rect 61556 11744 61568 11753
rect 60752 11716 61568 11744
rect 57532 11648 58204 11676
rect 60001 11679 60059 11685
rect 43625 11611 43683 11617
rect 43625 11577 43637 11611
rect 43671 11608 43683 11611
rect 43671 11580 45232 11608
rect 43671 11577 43683 11580
rect 43625 11571 43683 11577
rect 42935 11512 43024 11540
rect 45204 11540 45232 11580
rect 46750 11568 46756 11620
rect 46808 11608 46814 11620
rect 46808 11580 48360 11608
rect 46808 11568 46814 11580
rect 46014 11540 46020 11552
rect 45204 11512 46020 11540
rect 42935 11509 42947 11512
rect 42889 11503 42947 11509
rect 46014 11500 46020 11512
rect 46072 11500 46078 11552
rect 46382 11500 46388 11552
rect 46440 11540 46446 11552
rect 47578 11540 47584 11552
rect 46440 11512 47584 11540
rect 46440 11500 46446 11512
rect 47578 11500 47584 11512
rect 47636 11500 47642 11552
rect 47670 11500 47676 11552
rect 47728 11540 47734 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 47728 11512 47777 11540
rect 47728 11500 47734 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 48332 11540 48360 11580
rect 48774 11568 48780 11620
rect 48832 11608 48838 11620
rect 49804 11608 49832 11636
rect 52104 11608 52132 11636
rect 57532 11617 57560 11648
rect 60001 11645 60013 11679
rect 60047 11676 60059 11679
rect 60752 11676 60780 11716
rect 61556 11707 61568 11716
rect 61562 11704 61568 11707
rect 61620 11704 61626 11756
rect 61930 11704 61936 11756
rect 61988 11744 61994 11756
rect 63972 11753 64000 11784
rect 65628 11784 67180 11812
rect 65628 11753 65656 11784
rect 67174 11772 67180 11784
rect 67232 11772 67238 11824
rect 63221 11747 63279 11753
rect 63221 11744 63233 11747
rect 61988 11716 63233 11744
rect 61988 11704 61994 11716
rect 63221 11713 63233 11716
rect 63267 11713 63279 11747
rect 63221 11707 63279 11713
rect 63957 11747 64015 11753
rect 63957 11713 63969 11747
rect 64003 11713 64015 11747
rect 63957 11707 64015 11713
rect 65613 11747 65671 11753
rect 65613 11713 65625 11747
rect 65659 11713 65671 11747
rect 65613 11707 65671 11713
rect 60047 11648 60780 11676
rect 60829 11679 60887 11685
rect 60047 11645 60059 11648
rect 60001 11639 60059 11645
rect 60829 11645 60841 11679
rect 60875 11676 60887 11679
rect 61010 11676 61016 11688
rect 60875 11648 61016 11676
rect 60875 11645 60887 11648
rect 60829 11639 60887 11645
rect 61010 11636 61016 11648
rect 61068 11636 61074 11688
rect 61286 11676 61292 11688
rect 61247 11648 61292 11676
rect 61286 11636 61292 11648
rect 61344 11636 61350 11688
rect 62298 11636 62304 11688
rect 62356 11676 62362 11688
rect 65628 11676 65656 11707
rect 65702 11704 65708 11756
rect 65760 11744 65766 11756
rect 65869 11747 65927 11753
rect 65869 11744 65881 11747
rect 65760 11716 65881 11744
rect 65760 11704 65766 11716
rect 65869 11713 65881 11716
rect 65915 11713 65927 11747
rect 65869 11707 65927 11713
rect 67821 11747 67879 11753
rect 67821 11713 67833 11747
rect 67867 11744 67879 11747
rect 68296 11744 68324 11852
rect 70946 11840 70952 11852
rect 71004 11840 71010 11892
rect 71133 11883 71191 11889
rect 71133 11849 71145 11883
rect 71179 11880 71191 11883
rect 71179 11852 78904 11880
rect 71179 11849 71191 11852
rect 71133 11843 71191 11849
rect 69468 11815 69526 11821
rect 67867 11716 68324 11744
rect 68388 11784 68692 11812
rect 67867 11713 67879 11716
rect 67821 11707 67879 11713
rect 62356 11648 65656 11676
rect 62356 11636 62362 11648
rect 57517 11611 57575 11617
rect 48832 11580 49832 11608
rect 51046 11580 52132 11608
rect 52472 11580 54800 11608
rect 48832 11568 48838 11580
rect 49050 11540 49056 11552
rect 48332 11512 49056 11540
rect 47765 11503 47823 11509
rect 49050 11500 49056 11512
rect 49108 11500 49114 11552
rect 49145 11543 49203 11549
rect 49145 11509 49157 11543
rect 49191 11540 49203 11543
rect 51046 11540 51074 11580
rect 49191 11512 51074 11540
rect 51169 11543 51227 11549
rect 49191 11509 49203 11512
rect 49145 11503 49203 11509
rect 51169 11509 51181 11543
rect 51215 11540 51227 11543
rect 52472 11540 52500 11580
rect 51215 11512 52500 11540
rect 51215 11509 51227 11512
rect 51169 11503 51227 11509
rect 52546 11500 52552 11552
rect 52604 11540 52610 11552
rect 54386 11540 54392 11552
rect 52604 11512 54392 11540
rect 52604 11500 52610 11512
rect 54386 11500 54392 11512
rect 54444 11500 54450 11552
rect 54772 11540 54800 11580
rect 57517 11577 57529 11611
rect 57563 11577 57575 11611
rect 57517 11571 57575 11577
rect 60366 11568 60372 11620
rect 60424 11608 60430 11620
rect 64141 11611 64199 11617
rect 64141 11608 64153 11611
rect 60424 11580 60734 11608
rect 60424 11568 60430 11580
rect 60090 11540 60096 11552
rect 54772 11512 60096 11540
rect 60090 11500 60096 11512
rect 60148 11500 60154 11552
rect 60461 11543 60519 11549
rect 60461 11509 60473 11543
rect 60507 11540 60519 11543
rect 60550 11540 60556 11552
rect 60507 11512 60556 11540
rect 60507 11509 60519 11512
rect 60461 11503 60519 11509
rect 60550 11500 60556 11512
rect 60608 11500 60614 11552
rect 60706 11540 60734 11580
rect 62224 11580 64153 11608
rect 62224 11540 62252 11580
rect 64141 11577 64153 11580
rect 64187 11577 64199 11611
rect 64141 11571 64199 11577
rect 66993 11611 67051 11617
rect 66993 11577 67005 11611
rect 67039 11608 67051 11611
rect 68388 11608 68416 11784
rect 68554 11744 68560 11756
rect 68515 11716 68560 11744
rect 68554 11704 68560 11716
rect 68612 11704 68618 11756
rect 68664 11744 68692 11784
rect 69468 11781 69480 11815
rect 69514 11812 69526 11815
rect 71148 11812 71176 11843
rect 72326 11812 72332 11824
rect 69514 11784 71176 11812
rect 72287 11784 72332 11812
rect 69514 11781 69526 11784
rect 69468 11775 69526 11781
rect 72326 11772 72332 11784
rect 72384 11772 72390 11824
rect 72602 11772 72608 11824
rect 72660 11812 72666 11824
rect 74353 11815 74411 11821
rect 74353 11812 74365 11815
rect 72660 11784 74365 11812
rect 72660 11772 72666 11784
rect 74353 11781 74365 11784
rect 74399 11812 74411 11815
rect 74718 11812 74724 11824
rect 74399 11784 74724 11812
rect 74399 11781 74411 11784
rect 74353 11775 74411 11781
rect 74718 11772 74724 11784
rect 74776 11772 74782 11824
rect 78766 11812 78772 11824
rect 74828 11784 78772 11812
rect 74828 11744 74856 11784
rect 78766 11772 78772 11784
rect 78824 11772 78830 11824
rect 78876 11812 78904 11852
rect 78950 11840 78956 11892
rect 79008 11880 79014 11892
rect 79137 11883 79195 11889
rect 79137 11880 79149 11883
rect 79008 11852 79149 11880
rect 79008 11840 79014 11852
rect 79137 11849 79149 11852
rect 79183 11849 79195 11883
rect 81342 11880 81348 11892
rect 79137 11843 79195 11849
rect 79244 11852 81348 11880
rect 79244 11812 79272 11852
rect 81342 11840 81348 11852
rect 81400 11840 81406 11892
rect 82630 11840 82636 11892
rect 82688 11880 82694 11892
rect 84194 11880 84200 11892
rect 82688 11852 84200 11880
rect 82688 11840 82694 11852
rect 84194 11840 84200 11852
rect 84252 11840 84258 11892
rect 85393 11883 85451 11889
rect 85393 11849 85405 11883
rect 85439 11880 85451 11883
rect 86402 11880 86408 11892
rect 85439 11852 86408 11880
rect 85439 11849 85451 11852
rect 85393 11843 85451 11849
rect 86402 11840 86408 11852
rect 86460 11840 86466 11892
rect 86862 11840 86868 11892
rect 86920 11880 86926 11892
rect 87417 11883 87475 11889
rect 87417 11880 87429 11883
rect 86920 11852 87429 11880
rect 86920 11840 86926 11852
rect 87417 11849 87429 11852
rect 87463 11849 87475 11883
rect 88978 11880 88984 11892
rect 88939 11852 88984 11880
rect 87417 11843 87475 11849
rect 88978 11840 88984 11852
rect 89036 11840 89042 11892
rect 89088 11852 93808 11880
rect 78876 11784 79272 11812
rect 81434 11772 81440 11824
rect 81492 11812 81498 11824
rect 81492 11784 87368 11812
rect 81492 11772 81498 11784
rect 68664 11716 74856 11744
rect 74905 11747 74963 11753
rect 74905 11713 74917 11747
rect 74951 11744 74963 11747
rect 75914 11744 75920 11756
rect 74951 11716 75920 11744
rect 74951 11713 74963 11716
rect 74905 11707 74963 11713
rect 68741 11679 68799 11685
rect 68741 11645 68753 11679
rect 68787 11676 68799 11679
rect 68922 11676 68928 11688
rect 68787 11648 68928 11676
rect 68787 11645 68799 11648
rect 68741 11639 68799 11645
rect 68922 11636 68928 11648
rect 68980 11636 68986 11688
rect 69201 11679 69259 11685
rect 69201 11645 69213 11679
rect 69247 11645 69259 11679
rect 69201 11639 69259 11645
rect 69216 11608 69244 11639
rect 70946 11636 70952 11688
rect 71004 11676 71010 11688
rect 72694 11676 72700 11688
rect 71004 11648 72700 11676
rect 71004 11636 71010 11648
rect 72694 11636 72700 11648
rect 72752 11636 72758 11688
rect 73893 11679 73951 11685
rect 73893 11676 73905 11679
rect 72804 11648 73905 11676
rect 67039 11580 68416 11608
rect 68756 11580 69244 11608
rect 67039 11577 67051 11580
rect 66993 11571 67051 11577
rect 68756 11552 68784 11580
rect 60706 11512 62252 11540
rect 62669 11543 62727 11549
rect 62669 11509 62681 11543
rect 62715 11540 62727 11543
rect 63586 11540 63592 11552
rect 62715 11512 63592 11540
rect 62715 11509 62727 11512
rect 62669 11503 62727 11509
rect 63586 11500 63592 11512
rect 63644 11500 63650 11552
rect 65058 11540 65064 11552
rect 65019 11512 65064 11540
rect 65058 11500 65064 11512
rect 65116 11540 65122 11552
rect 65610 11540 65616 11552
rect 65116 11512 65616 11540
rect 65116 11500 65122 11512
rect 65610 11500 65616 11512
rect 65668 11500 65674 11552
rect 65886 11500 65892 11552
rect 65944 11540 65950 11552
rect 67637 11543 67695 11549
rect 67637 11540 67649 11543
rect 65944 11512 67649 11540
rect 65944 11500 65950 11512
rect 67637 11509 67649 11512
rect 67683 11509 67695 11543
rect 68370 11540 68376 11552
rect 68331 11512 68376 11540
rect 67637 11503 67695 11509
rect 68370 11500 68376 11512
rect 68428 11500 68434 11552
rect 68738 11500 68744 11552
rect 68796 11500 68802 11552
rect 69216 11540 69244 11580
rect 70210 11568 70216 11620
rect 70268 11608 70274 11620
rect 72602 11608 72608 11620
rect 70268 11580 72608 11608
rect 70268 11568 70274 11580
rect 72602 11568 72608 11580
rect 72660 11568 72666 11620
rect 70302 11540 70308 11552
rect 69216 11512 70308 11540
rect 70302 11500 70308 11512
rect 70360 11500 70366 11552
rect 70578 11540 70584 11552
rect 70539 11512 70584 11540
rect 70578 11500 70584 11512
rect 70636 11500 70642 11552
rect 71866 11500 71872 11552
rect 71924 11540 71930 11552
rect 72804 11540 72832 11648
rect 73893 11645 73905 11648
rect 73939 11676 73951 11679
rect 74920 11676 74948 11707
rect 75914 11704 75920 11716
rect 75972 11704 75978 11756
rect 76190 11744 76196 11756
rect 76024 11716 76196 11744
rect 76024 11676 76052 11716
rect 76190 11704 76196 11716
rect 76248 11704 76254 11756
rect 76368 11747 76426 11753
rect 76368 11713 76380 11747
rect 76414 11744 76426 11747
rect 77294 11744 77300 11756
rect 76414 11716 77300 11744
rect 76414 11713 76426 11716
rect 76368 11707 76426 11713
rect 77294 11704 77300 11716
rect 77352 11704 77358 11756
rect 80261 11747 80319 11753
rect 80261 11713 80273 11747
rect 80307 11744 80319 11747
rect 80307 11716 80468 11744
rect 80307 11713 80319 11716
rect 80261 11707 80319 11713
rect 73939 11648 74948 11676
rect 75012 11648 76052 11676
rect 76101 11679 76159 11685
rect 73939 11645 73951 11648
rect 73893 11639 73951 11645
rect 75012 11608 75040 11648
rect 76101 11645 76113 11679
rect 76147 11645 76159 11679
rect 78674 11676 78680 11688
rect 76101 11639 76159 11645
rect 77128 11648 78680 11676
rect 75089 11611 75147 11617
rect 75089 11608 75101 11611
rect 75012 11580 75101 11608
rect 75089 11577 75101 11580
rect 75135 11577 75147 11611
rect 75914 11608 75920 11620
rect 75089 11571 75147 11577
rect 75196 11580 75920 11608
rect 72970 11540 72976 11552
rect 71924 11512 72832 11540
rect 72931 11512 72976 11540
rect 71924 11500 71930 11512
rect 72970 11500 72976 11512
rect 73028 11500 73034 11552
rect 74718 11500 74724 11552
rect 74776 11540 74782 11552
rect 75196 11540 75224 11580
rect 75914 11568 75920 11580
rect 75972 11608 75978 11620
rect 76116 11608 76144 11639
rect 75972 11580 76144 11608
rect 75972 11568 75978 11580
rect 74776 11512 75224 11540
rect 74776 11500 74782 11512
rect 75270 11500 75276 11552
rect 75328 11540 75334 11552
rect 77128 11540 77156 11648
rect 78674 11636 78680 11648
rect 78732 11636 78738 11688
rect 80440 11676 80468 11716
rect 80514 11704 80520 11756
rect 80572 11744 80578 11756
rect 80572 11716 80665 11744
rect 80572 11704 80578 11716
rect 80624 11676 80652 11716
rect 81618 11704 81624 11756
rect 81676 11744 81682 11756
rect 83001 11747 83059 11753
rect 83001 11744 83013 11747
rect 81676 11716 83013 11744
rect 81676 11704 81682 11716
rect 83001 11713 83013 11716
rect 83047 11713 83059 11747
rect 83001 11707 83059 11713
rect 84013 11747 84071 11753
rect 84013 11713 84025 11747
rect 84059 11744 84071 11747
rect 86218 11744 86224 11756
rect 84059 11716 86224 11744
rect 84059 11713 84071 11716
rect 84013 11707 84071 11713
rect 86218 11704 86224 11716
rect 86276 11704 86282 11756
rect 86517 11747 86575 11753
rect 86517 11713 86529 11747
rect 86563 11744 86575 11747
rect 86773 11747 86831 11753
rect 86563 11716 86724 11744
rect 86563 11713 86575 11716
rect 86517 11707 86575 11713
rect 83918 11676 83924 11688
rect 80440 11648 80560 11676
rect 80624 11648 83924 11676
rect 77481 11611 77539 11617
rect 77481 11577 77493 11611
rect 77527 11608 77539 11611
rect 79134 11608 79140 11620
rect 77527 11580 79140 11608
rect 77527 11577 77539 11580
rect 77481 11571 77539 11577
rect 79134 11568 79140 11580
rect 79192 11568 79198 11620
rect 80532 11608 80560 11648
rect 83918 11636 83924 11648
rect 83976 11636 83982 11688
rect 84102 11636 84108 11688
rect 84160 11676 84166 11688
rect 84197 11679 84255 11685
rect 84197 11676 84209 11679
rect 84160 11648 84209 11676
rect 84160 11636 84166 11648
rect 84197 11645 84209 11648
rect 84243 11645 84255 11679
rect 86696 11676 86724 11716
rect 86773 11713 86785 11747
rect 86819 11744 86831 11747
rect 86862 11744 86868 11756
rect 86819 11716 86868 11744
rect 86819 11713 86831 11716
rect 86773 11707 86831 11713
rect 86862 11704 86868 11716
rect 86920 11704 86926 11756
rect 86954 11704 86960 11756
rect 87012 11744 87018 11756
rect 87233 11747 87291 11753
rect 87233 11744 87245 11747
rect 87012 11716 87245 11744
rect 87012 11704 87018 11716
rect 87233 11713 87245 11716
rect 87279 11713 87291 11747
rect 87340 11744 87368 11784
rect 87506 11772 87512 11824
rect 87564 11812 87570 11824
rect 89088 11812 89116 11852
rect 87564 11784 89116 11812
rect 87564 11772 87570 11784
rect 89254 11772 89260 11824
rect 89312 11812 89318 11824
rect 89898 11812 89904 11824
rect 89312 11784 89904 11812
rect 89312 11772 89318 11784
rect 89898 11772 89904 11784
rect 89956 11812 89962 11824
rect 90094 11815 90152 11821
rect 90094 11812 90106 11815
rect 89956 11784 90106 11812
rect 89956 11772 89962 11784
rect 90094 11781 90106 11784
rect 90140 11781 90152 11815
rect 93670 11812 93676 11824
rect 90094 11775 90152 11781
rect 90284 11784 93676 11812
rect 90284 11744 90312 11784
rect 93670 11772 93676 11784
rect 93728 11772 93734 11824
rect 93780 11812 93808 11852
rect 94590 11840 94596 11892
rect 94648 11880 94654 11892
rect 94961 11883 95019 11889
rect 94961 11880 94973 11883
rect 94648 11852 94973 11880
rect 94648 11840 94654 11852
rect 94961 11849 94973 11852
rect 95007 11849 95019 11883
rect 94961 11843 95019 11849
rect 96154 11840 96160 11892
rect 96212 11880 96218 11892
rect 97813 11883 97871 11889
rect 97813 11880 97825 11883
rect 96212 11852 97825 11880
rect 96212 11840 96218 11852
rect 97813 11849 97825 11852
rect 97859 11880 97871 11883
rect 98178 11880 98184 11892
rect 97859 11852 98184 11880
rect 97859 11849 97871 11852
rect 97813 11843 97871 11849
rect 98178 11840 98184 11852
rect 98236 11840 98242 11892
rect 98454 11880 98460 11892
rect 98415 11852 98460 11880
rect 98454 11840 98460 11852
rect 98512 11840 98518 11892
rect 99926 11880 99932 11892
rect 99839 11852 99932 11880
rect 99926 11840 99932 11852
rect 99984 11880 99990 11892
rect 100202 11880 100208 11892
rect 99984 11852 100208 11880
rect 99984 11840 99990 11852
rect 100202 11840 100208 11852
rect 100260 11880 100266 11892
rect 103054 11880 103060 11892
rect 100260 11852 103060 11880
rect 100260 11840 100266 11852
rect 103054 11840 103060 11852
rect 103112 11840 103118 11892
rect 103514 11880 103520 11892
rect 103427 11852 103520 11880
rect 103514 11840 103520 11852
rect 103572 11880 103578 11892
rect 104250 11880 104256 11892
rect 103572 11852 104256 11880
rect 103572 11840 103578 11852
rect 104250 11840 104256 11852
rect 104308 11840 104314 11892
rect 104529 11883 104587 11889
rect 104529 11849 104541 11883
rect 104575 11880 104587 11883
rect 104710 11880 104716 11892
rect 104575 11852 104716 11880
rect 104575 11849 104587 11852
rect 104529 11843 104587 11849
rect 104710 11840 104716 11852
rect 104768 11840 104774 11892
rect 106182 11840 106188 11892
rect 106240 11880 106246 11892
rect 108577 11883 108635 11889
rect 108577 11880 108589 11883
rect 106240 11852 108589 11880
rect 106240 11840 106246 11852
rect 108577 11849 108589 11852
rect 108623 11880 108635 11883
rect 108666 11880 108672 11892
rect 108623 11852 108672 11880
rect 108623 11849 108635 11852
rect 108577 11843 108635 11849
rect 108666 11840 108672 11852
rect 108724 11840 108730 11892
rect 109678 11880 109684 11892
rect 108776 11852 109034 11880
rect 109591 11852 109684 11880
rect 101582 11812 101588 11824
rect 93780 11784 101588 11812
rect 101582 11772 101588 11784
rect 101640 11772 101646 11824
rect 108776 11812 108804 11852
rect 101692 11784 108804 11812
rect 109006 11812 109034 11852
rect 109678 11840 109684 11852
rect 109736 11880 109742 11892
rect 112346 11880 112352 11892
rect 109736 11852 112352 11880
rect 109736 11840 109742 11852
rect 112346 11840 112352 11852
rect 112404 11840 112410 11892
rect 113266 11880 113272 11892
rect 113227 11852 113272 11880
rect 113266 11840 113272 11852
rect 113324 11840 113330 11892
rect 114830 11880 114836 11892
rect 114743 11852 114836 11880
rect 114830 11840 114836 11852
rect 114888 11880 114894 11892
rect 118694 11880 118700 11892
rect 114888 11852 118700 11880
rect 114888 11840 114894 11852
rect 118694 11840 118700 11852
rect 118752 11840 118758 11892
rect 119062 11880 119068 11892
rect 119023 11852 119068 11880
rect 119062 11840 119068 11852
rect 119120 11840 119126 11892
rect 119430 11840 119436 11892
rect 119488 11880 119494 11892
rect 125134 11880 125140 11892
rect 119488 11852 125140 11880
rect 119488 11840 119494 11852
rect 125134 11840 125140 11852
rect 125192 11840 125198 11892
rect 125594 11880 125600 11892
rect 125244 11852 125447 11880
rect 125555 11852 125600 11880
rect 125244 11812 125272 11852
rect 109006 11784 125272 11812
rect 125419 11812 125447 11852
rect 125594 11840 125600 11852
rect 125652 11840 125658 11892
rect 129277 11883 129335 11889
rect 129277 11880 129289 11883
rect 126348 11852 129289 11880
rect 126348 11812 126376 11852
rect 129277 11849 129289 11852
rect 129323 11849 129335 11883
rect 130194 11880 130200 11892
rect 130155 11852 130200 11880
rect 129277 11843 129335 11849
rect 130194 11840 130200 11852
rect 130252 11840 130258 11892
rect 132310 11840 132316 11892
rect 132368 11880 132374 11892
rect 134978 11880 134984 11892
rect 132368 11852 134984 11880
rect 132368 11840 132374 11852
rect 134978 11840 134984 11852
rect 135036 11840 135042 11892
rect 135254 11840 135260 11892
rect 135312 11880 135318 11892
rect 135349 11883 135407 11889
rect 135349 11880 135361 11883
rect 135312 11852 135361 11880
rect 135312 11840 135318 11852
rect 135349 11849 135361 11852
rect 135395 11849 135407 11883
rect 135349 11843 135407 11849
rect 135456 11852 138014 11880
rect 125419 11784 126376 11812
rect 87340 11716 88104 11744
rect 87233 11707 87291 11713
rect 87966 11676 87972 11688
rect 86696 11648 87972 11676
rect 84197 11639 84255 11645
rect 87966 11636 87972 11648
rect 88024 11636 88030 11688
rect 88076 11676 88104 11716
rect 89364 11716 90312 11744
rect 91456 11747 91514 11753
rect 89364 11676 89392 11716
rect 91456 11713 91468 11747
rect 91502 11744 91514 11747
rect 92750 11744 92756 11756
rect 91502 11716 92756 11744
rect 91502 11713 91514 11716
rect 91456 11707 91514 11713
rect 92750 11704 92756 11716
rect 92808 11704 92814 11756
rect 92842 11704 92848 11756
rect 92900 11744 92906 11756
rect 93121 11747 93179 11753
rect 93121 11744 93133 11747
rect 92900 11716 93133 11744
rect 92900 11704 92906 11716
rect 93121 11713 93133 11716
rect 93167 11744 93179 11747
rect 93394 11744 93400 11756
rect 93167 11716 93400 11744
rect 93167 11713 93179 11716
rect 93121 11707 93179 11713
rect 93394 11704 93400 11716
rect 93452 11704 93458 11756
rect 93688 11744 93716 11772
rect 94314 11744 94320 11756
rect 93688 11716 94320 11744
rect 94314 11704 94320 11716
rect 94372 11704 94378 11756
rect 94409 11747 94467 11753
rect 94409 11713 94421 11747
rect 94455 11744 94467 11747
rect 95050 11744 95056 11756
rect 94455 11716 95056 11744
rect 94455 11713 94467 11716
rect 94409 11707 94467 11713
rect 95050 11704 95056 11716
rect 95108 11704 95114 11756
rect 95145 11747 95203 11753
rect 95145 11713 95157 11747
rect 95191 11713 95203 11747
rect 95145 11707 95203 11713
rect 88076 11648 89392 11676
rect 90361 11679 90419 11685
rect 90361 11645 90373 11679
rect 90407 11676 90419 11679
rect 90450 11676 90456 11688
rect 90407 11648 90456 11676
rect 90407 11645 90419 11648
rect 90361 11639 90419 11645
rect 90450 11636 90456 11648
rect 90508 11676 90514 11688
rect 90634 11676 90640 11688
rect 90508 11648 90640 11676
rect 90508 11636 90514 11648
rect 90634 11636 90640 11648
rect 90692 11676 90698 11688
rect 91189 11679 91247 11685
rect 91189 11676 91201 11679
rect 90692 11648 91201 11676
rect 90692 11636 90698 11648
rect 91189 11645 91201 11648
rect 91235 11645 91247 11679
rect 94682 11676 94688 11688
rect 91189 11639 91247 11645
rect 92584 11648 94688 11676
rect 81069 11611 81127 11617
rect 81069 11608 81081 11611
rect 80532 11580 81081 11608
rect 81069 11577 81081 11580
rect 81115 11608 81127 11611
rect 81115 11580 84976 11608
rect 81115 11577 81127 11580
rect 81069 11571 81127 11577
rect 75328 11512 77156 11540
rect 75328 11500 75334 11512
rect 77938 11500 77944 11552
rect 77996 11540 78002 11552
rect 78033 11543 78091 11549
rect 78033 11540 78045 11543
rect 77996 11512 78045 11540
rect 77996 11500 78002 11512
rect 78033 11509 78045 11512
rect 78079 11509 78091 11543
rect 82814 11540 82820 11552
rect 82775 11512 82820 11540
rect 78033 11503 78091 11509
rect 82814 11500 82820 11512
rect 82872 11500 82878 11552
rect 83826 11540 83832 11552
rect 83787 11512 83832 11540
rect 83826 11500 83832 11512
rect 83884 11500 83890 11552
rect 84838 11540 84844 11552
rect 84799 11512 84844 11540
rect 84838 11500 84844 11512
rect 84896 11500 84902 11552
rect 84948 11540 84976 11580
rect 86862 11568 86868 11620
rect 86920 11608 86926 11620
rect 89254 11608 89260 11620
rect 86920 11580 89260 11608
rect 86920 11568 86926 11580
rect 89254 11568 89260 11580
rect 89312 11568 89318 11620
rect 92584 11617 92612 11648
rect 94682 11636 94688 11648
rect 94740 11636 94746 11688
rect 95160 11676 95188 11707
rect 95234 11704 95240 11756
rect 95292 11744 95298 11756
rect 96157 11747 96215 11753
rect 96157 11744 96169 11747
rect 95292 11716 96169 11744
rect 95292 11704 95298 11716
rect 96157 11713 96169 11716
rect 96203 11713 96215 11747
rect 96157 11707 96215 11713
rect 96614 11704 96620 11756
rect 96672 11744 96678 11756
rect 97261 11747 97319 11753
rect 97261 11744 97273 11747
rect 96672 11716 97273 11744
rect 96672 11704 96678 11716
rect 97261 11713 97273 11716
rect 97307 11713 97319 11747
rect 97261 11707 97319 11713
rect 99006 11704 99012 11756
rect 99064 11744 99070 11756
rect 101692 11744 101720 11784
rect 99064 11716 101720 11744
rect 99064 11704 99070 11716
rect 101766 11704 101772 11756
rect 101824 11753 101830 11756
rect 101824 11744 101836 11753
rect 101824 11716 101869 11744
rect 101824 11707 101836 11716
rect 101824 11704 101830 11707
rect 101950 11704 101956 11756
rect 102008 11744 102014 11756
rect 105653 11747 105711 11753
rect 102008 11716 104664 11744
rect 102008 11704 102014 11716
rect 96430 11676 96436 11688
rect 95160 11648 96436 11676
rect 96430 11636 96436 11648
rect 96488 11636 96494 11688
rect 96706 11636 96712 11688
rect 96764 11676 96770 11688
rect 96801 11679 96859 11685
rect 96801 11676 96813 11679
rect 96764 11648 96813 11676
rect 96764 11636 96770 11648
rect 96801 11645 96813 11648
rect 96847 11676 96859 11679
rect 99024 11676 99052 11704
rect 96847 11648 99052 11676
rect 96847 11645 96859 11648
rect 96801 11639 96859 11645
rect 99374 11636 99380 11688
rect 99432 11676 99438 11688
rect 102045 11679 102103 11685
rect 99432 11648 99477 11676
rect 99432 11636 99438 11648
rect 102045 11645 102057 11679
rect 102091 11676 102103 11679
rect 102091 11648 102640 11676
rect 102091 11645 102103 11648
rect 102045 11639 102103 11645
rect 92569 11611 92627 11617
rect 92569 11577 92581 11611
rect 92615 11577 92627 11611
rect 92569 11571 92627 11577
rect 92676 11580 93164 11608
rect 87782 11540 87788 11552
rect 84948 11512 87788 11540
rect 87782 11500 87788 11512
rect 87840 11500 87846 11552
rect 88058 11500 88064 11552
rect 88116 11540 88122 11552
rect 89990 11540 89996 11552
rect 88116 11512 89996 11540
rect 88116 11500 88122 11512
rect 89990 11500 89996 11512
rect 90048 11500 90054 11552
rect 90082 11500 90088 11552
rect 90140 11540 90146 11552
rect 92676 11540 92704 11580
rect 90140 11512 92704 11540
rect 93136 11540 93164 11580
rect 93486 11568 93492 11620
rect 93544 11608 93550 11620
rect 94225 11611 94283 11617
rect 94225 11608 94237 11611
rect 93544 11580 94237 11608
rect 93544 11568 93550 11580
rect 94225 11577 94237 11580
rect 94271 11577 94283 11611
rect 101030 11608 101036 11620
rect 94225 11571 94283 11577
rect 94332 11580 101036 11608
rect 94332 11540 94360 11580
rect 101030 11568 101036 11580
rect 101088 11568 101094 11620
rect 93136 11512 94360 11540
rect 90140 11500 90146 11512
rect 94406 11500 94412 11552
rect 94464 11540 94470 11552
rect 95605 11543 95663 11549
rect 95605 11540 95617 11543
rect 94464 11512 95617 11540
rect 94464 11500 94470 11512
rect 95605 11509 95617 11512
rect 95651 11509 95663 11543
rect 100662 11540 100668 11552
rect 100623 11512 100668 11540
rect 95605 11503 95663 11509
rect 100662 11500 100668 11512
rect 100720 11500 100726 11552
rect 102612 11549 102640 11648
rect 102597 11543 102655 11549
rect 102597 11509 102609 11543
rect 102643 11540 102655 11543
rect 103422 11540 103428 11552
rect 102643 11512 103428 11540
rect 102643 11509 102655 11512
rect 102597 11503 102655 11509
rect 103422 11500 103428 11512
rect 103480 11500 103486 11552
rect 104636 11540 104664 11716
rect 105653 11713 105665 11747
rect 105699 11744 105711 11747
rect 107470 11744 107476 11756
rect 105699 11716 107476 11744
rect 105699 11713 105711 11716
rect 105653 11707 105711 11713
rect 107470 11704 107476 11716
rect 107528 11704 107534 11756
rect 108117 11747 108175 11753
rect 108117 11713 108129 11747
rect 108163 11744 108175 11747
rect 108758 11744 108764 11756
rect 108163 11716 108764 11744
rect 108163 11713 108175 11716
rect 108117 11707 108175 11713
rect 108758 11704 108764 11716
rect 108816 11704 108822 11756
rect 108850 11704 108856 11756
rect 108908 11744 108914 11756
rect 112070 11744 112076 11756
rect 108908 11716 112076 11744
rect 108908 11704 108914 11716
rect 112070 11704 112076 11716
rect 112128 11704 112134 11756
rect 112162 11704 112168 11756
rect 112220 11744 112226 11756
rect 112533 11747 112591 11753
rect 112533 11744 112545 11747
rect 112220 11716 112545 11744
rect 112220 11704 112226 11716
rect 112533 11713 112545 11716
rect 112579 11713 112591 11747
rect 112533 11707 112591 11713
rect 113453 11747 113511 11753
rect 113453 11713 113465 11747
rect 113499 11744 113511 11747
rect 113634 11744 113640 11756
rect 113499 11716 113640 11744
rect 113499 11713 113511 11716
rect 113453 11707 113511 11713
rect 113634 11704 113640 11716
rect 113692 11704 113698 11756
rect 113836 11716 115612 11744
rect 105909 11679 105967 11685
rect 105909 11645 105921 11679
rect 105955 11676 105967 11679
rect 107562 11676 107568 11688
rect 105955 11648 107568 11676
rect 105955 11645 105967 11648
rect 105909 11639 105967 11645
rect 107562 11636 107568 11648
rect 107620 11636 107626 11688
rect 108666 11636 108672 11688
rect 108724 11676 108730 11688
rect 113836 11676 113864 11716
rect 115474 11676 115480 11688
rect 108724 11648 113864 11676
rect 115435 11648 115480 11676
rect 108724 11636 108730 11648
rect 115474 11636 115480 11648
rect 115532 11636 115538 11688
rect 115584 11676 115612 11716
rect 115658 11704 115664 11756
rect 115716 11744 115722 11756
rect 116394 11744 116400 11756
rect 115716 11716 116400 11744
rect 115716 11704 115722 11716
rect 116394 11704 116400 11716
rect 116452 11704 116458 11756
rect 117429 11747 117487 11753
rect 117429 11713 117441 11747
rect 117475 11744 117487 11747
rect 117475 11716 118096 11744
rect 117475 11713 117487 11716
rect 117429 11707 117487 11713
rect 117685 11679 117743 11685
rect 115584 11648 116440 11676
rect 106366 11608 106372 11620
rect 106327 11580 106372 11608
rect 106366 11568 106372 11580
rect 106424 11568 106430 11620
rect 107194 11608 107200 11620
rect 106476 11580 107200 11608
rect 106476 11540 106504 11580
rect 107194 11568 107200 11580
rect 107252 11568 107258 11620
rect 107286 11568 107292 11620
rect 107344 11608 107350 11620
rect 111245 11611 111303 11617
rect 107344 11580 111196 11608
rect 107344 11568 107350 11580
rect 107010 11540 107016 11552
rect 104636 11512 106504 11540
rect 106971 11512 107016 11540
rect 107010 11500 107016 11512
rect 107068 11500 107074 11552
rect 107378 11500 107384 11552
rect 107436 11540 107442 11552
rect 107933 11543 107991 11549
rect 107933 11540 107945 11543
rect 107436 11512 107945 11540
rect 107436 11500 107442 11512
rect 107933 11509 107945 11512
rect 107979 11509 107991 11543
rect 107933 11503 107991 11509
rect 109034 11500 109040 11552
rect 109092 11540 109098 11552
rect 109678 11540 109684 11552
rect 109092 11512 109684 11540
rect 109092 11500 109098 11512
rect 109678 11500 109684 11512
rect 109736 11500 109742 11552
rect 110233 11543 110291 11549
rect 110233 11509 110245 11543
rect 110279 11540 110291 11543
rect 110414 11540 110420 11552
rect 110279 11512 110420 11540
rect 110279 11509 110291 11512
rect 110233 11503 110291 11509
rect 110414 11500 110420 11512
rect 110472 11500 110478 11552
rect 111168 11540 111196 11580
rect 111245 11577 111257 11611
rect 111291 11608 111303 11611
rect 112530 11608 112536 11620
rect 111291 11580 112536 11608
rect 111291 11577 111303 11580
rect 111245 11571 111303 11577
rect 112530 11568 112536 11580
rect 112588 11568 112594 11620
rect 116305 11611 116363 11617
rect 116305 11608 116317 11611
rect 112640 11580 116317 11608
rect 112640 11540 112668 11580
rect 116305 11577 116317 11580
rect 116351 11577 116363 11611
rect 116305 11571 116363 11577
rect 111168 11512 112668 11540
rect 112714 11500 112720 11552
rect 112772 11540 112778 11552
rect 113913 11543 113971 11549
rect 113913 11540 113925 11543
rect 112772 11512 113925 11540
rect 112772 11500 112778 11512
rect 113913 11509 113925 11512
rect 113959 11509 113971 11543
rect 115842 11540 115848 11552
rect 115803 11512 115848 11540
rect 113913 11503 113971 11509
rect 115842 11500 115848 11512
rect 115900 11500 115906 11552
rect 116412 11540 116440 11648
rect 117685 11645 117697 11679
rect 117731 11645 117743 11679
rect 117685 11639 117743 11645
rect 117314 11540 117320 11552
rect 116412 11512 117320 11540
rect 117314 11500 117320 11512
rect 117372 11500 117378 11552
rect 117406 11500 117412 11552
rect 117464 11540 117470 11552
rect 117700 11540 117728 11639
rect 118068 11608 118096 11716
rect 118234 11704 118240 11756
rect 118292 11744 118298 11756
rect 118329 11747 118387 11753
rect 118329 11744 118341 11747
rect 118292 11716 118341 11744
rect 118292 11704 118298 11716
rect 118329 11713 118341 11716
rect 118375 11744 118387 11747
rect 120445 11747 120503 11753
rect 120445 11744 120457 11747
rect 118375 11716 120457 11744
rect 118375 11713 118387 11716
rect 118329 11707 118387 11713
rect 120445 11713 120457 11716
rect 120491 11713 120503 11747
rect 121178 11744 121184 11756
rect 121139 11716 121184 11744
rect 120445 11707 120503 11713
rect 121178 11704 121184 11716
rect 121236 11704 121242 11756
rect 122101 11747 122159 11753
rect 122101 11744 122113 11747
rect 121288 11716 122113 11744
rect 118510 11676 118516 11688
rect 118471 11648 118516 11676
rect 118510 11636 118516 11648
rect 118568 11636 118574 11688
rect 118694 11636 118700 11688
rect 118752 11676 118758 11688
rect 118752 11648 119016 11676
rect 118752 11636 118758 11648
rect 118878 11608 118884 11620
rect 118068 11580 118884 11608
rect 118878 11568 118884 11580
rect 118936 11568 118942 11620
rect 118988 11608 119016 11648
rect 119154 11636 119160 11688
rect 119212 11676 119218 11688
rect 119985 11679 120043 11685
rect 119985 11676 119997 11679
rect 119212 11648 119997 11676
rect 119212 11636 119218 11648
rect 119985 11645 119997 11648
rect 120031 11676 120043 11679
rect 121288 11676 121316 11716
rect 122101 11713 122113 11716
rect 122147 11744 122159 11747
rect 125042 11744 125048 11756
rect 122147 11716 125048 11744
rect 122147 11713 122159 11716
rect 122101 11707 122159 11713
rect 125042 11704 125048 11716
rect 125100 11704 125106 11756
rect 125962 11744 125968 11756
rect 125566 11716 125968 11744
rect 120031 11648 121316 11676
rect 120031 11645 120043 11648
rect 119985 11639 120043 11645
rect 121362 11636 121368 11688
rect 121420 11676 121426 11688
rect 121420 11648 121465 11676
rect 121420 11636 121426 11648
rect 122006 11636 122012 11688
rect 122064 11676 122070 11688
rect 123846 11676 123852 11688
rect 122064 11648 123852 11676
rect 122064 11636 122070 11648
rect 123846 11636 123852 11648
rect 123904 11636 123910 11688
rect 125134 11636 125140 11688
rect 125192 11676 125198 11688
rect 125566 11676 125594 11716
rect 125962 11704 125968 11716
rect 126020 11704 126026 11756
rect 126348 11753 126376 11784
rect 126517 11815 126575 11821
rect 126517 11781 126529 11815
rect 126563 11812 126575 11815
rect 126563 11784 128032 11812
rect 126563 11781 126575 11784
rect 126517 11775 126575 11781
rect 126333 11747 126391 11753
rect 126072 11716 126284 11744
rect 125192 11648 125594 11676
rect 125192 11636 125198 11648
rect 118988 11580 119752 11608
rect 118142 11540 118148 11552
rect 117464 11512 117728 11540
rect 118103 11512 118148 11540
rect 117464 11500 117470 11512
rect 118142 11500 118148 11512
rect 118200 11500 118206 11552
rect 118510 11500 118516 11552
rect 118568 11540 118574 11552
rect 119614 11540 119620 11552
rect 118568 11512 119620 11540
rect 118568 11500 118574 11512
rect 119614 11500 119620 11512
rect 119672 11500 119678 11552
rect 119724 11540 119752 11580
rect 124950 11568 124956 11620
rect 125008 11608 125014 11620
rect 126072 11608 126100 11716
rect 126149 11679 126207 11685
rect 126149 11645 126161 11679
rect 126195 11645 126207 11679
rect 126256 11676 126284 11716
rect 126333 11713 126345 11747
rect 126379 11713 126391 11747
rect 126974 11744 126980 11756
rect 126935 11716 126980 11744
rect 126333 11707 126391 11713
rect 126974 11704 126980 11716
rect 127032 11704 127038 11756
rect 127158 11744 127164 11756
rect 127119 11716 127164 11744
rect 127158 11704 127164 11716
rect 127216 11704 127222 11756
rect 127342 11744 127348 11756
rect 127303 11716 127348 11744
rect 127342 11704 127348 11716
rect 127400 11704 127406 11756
rect 128004 11753 128032 11784
rect 129366 11772 129372 11824
rect 129424 11812 129430 11824
rect 135456 11812 135484 11852
rect 137186 11812 137192 11824
rect 129424 11784 135484 11812
rect 135548 11784 137192 11812
rect 129424 11772 129430 11784
rect 127989 11747 128047 11753
rect 127989 11713 128001 11747
rect 128035 11713 128047 11747
rect 128630 11744 128636 11756
rect 128591 11716 128636 11744
rect 127989 11707 128047 11713
rect 128630 11704 128636 11716
rect 128688 11744 128694 11756
rect 130749 11747 130807 11753
rect 130749 11744 130761 11747
rect 128688 11716 130761 11744
rect 128688 11704 128694 11716
rect 130749 11713 130761 11716
rect 130795 11713 130807 11747
rect 134173 11747 134231 11753
rect 130749 11707 130807 11713
rect 130856 11716 132540 11744
rect 126992 11676 127020 11704
rect 127250 11676 127256 11688
rect 126256 11648 127256 11676
rect 126149 11639 126207 11645
rect 125008 11580 126100 11608
rect 126164 11608 126192 11639
rect 127250 11636 127256 11648
rect 127308 11636 127314 11688
rect 128354 11676 128360 11688
rect 127360 11648 128360 11676
rect 127360 11608 127388 11648
rect 128354 11636 128360 11648
rect 128412 11676 128418 11688
rect 128817 11679 128875 11685
rect 128817 11676 128829 11679
rect 128412 11648 128829 11676
rect 128412 11636 128418 11648
rect 128817 11645 128829 11648
rect 128863 11676 128875 11679
rect 130856 11676 130884 11716
rect 132512 11688 132540 11716
rect 134173 11713 134185 11747
rect 134219 11744 134231 11747
rect 134219 11716 134932 11744
rect 134219 11713 134231 11716
rect 134173 11707 134231 11713
rect 132494 11676 132500 11688
rect 128863 11648 130884 11676
rect 132407 11648 132500 11676
rect 128863 11645 128875 11648
rect 128817 11639 128875 11645
rect 132494 11636 132500 11648
rect 132552 11676 132558 11688
rect 133414 11676 133420 11688
rect 132552 11648 133420 11676
rect 132552 11636 132558 11648
rect 133414 11636 133420 11648
rect 133472 11636 133478 11688
rect 134426 11676 134432 11688
rect 134387 11648 134432 11676
rect 134426 11636 134432 11648
rect 134484 11636 134490 11688
rect 133230 11608 133236 11620
rect 126164 11580 127388 11608
rect 127728 11580 133236 11608
rect 125008 11568 125014 11580
rect 120442 11540 120448 11552
rect 119724 11512 120448 11540
rect 120442 11500 120448 11512
rect 120500 11500 120506 11552
rect 120534 11500 120540 11552
rect 120592 11540 120598 11552
rect 120997 11543 121055 11549
rect 120997 11540 121009 11543
rect 120592 11512 121009 11540
rect 120592 11500 120598 11512
rect 120997 11509 121009 11512
rect 121043 11509 121055 11543
rect 121914 11540 121920 11552
rect 121875 11512 121920 11540
rect 120997 11503 121055 11509
rect 121914 11500 121920 11512
rect 121972 11500 121978 11552
rect 122653 11543 122711 11549
rect 122653 11509 122665 11543
rect 122699 11540 122711 11543
rect 122742 11540 122748 11552
rect 122699 11512 122748 11540
rect 122699 11509 122711 11512
rect 122653 11503 122711 11509
rect 122742 11500 122748 11512
rect 122800 11500 122806 11552
rect 123202 11540 123208 11552
rect 123163 11512 123208 11540
rect 123202 11500 123208 11512
rect 123260 11500 123266 11552
rect 123662 11540 123668 11552
rect 123623 11512 123668 11540
rect 123662 11500 123668 11512
rect 123720 11500 123726 11552
rect 124214 11540 124220 11552
rect 124175 11512 124220 11540
rect 124214 11500 124220 11512
rect 124272 11500 124278 11552
rect 125502 11500 125508 11552
rect 125560 11540 125566 11552
rect 127728 11540 127756 11580
rect 133230 11568 133236 11580
rect 133288 11568 133294 11620
rect 134904 11608 134932 11716
rect 134978 11636 134984 11688
rect 135036 11676 135042 11688
rect 135548 11676 135576 11784
rect 137186 11772 137192 11784
rect 137244 11772 137250 11824
rect 137986 11812 138014 11852
rect 138474 11840 138480 11892
rect 138532 11880 138538 11892
rect 138658 11880 138664 11892
rect 138532 11852 138664 11880
rect 138532 11840 138538 11852
rect 138658 11840 138664 11852
rect 138716 11880 138722 11892
rect 143810 11880 143816 11892
rect 138716 11852 138879 11880
rect 138716 11840 138722 11852
rect 138851 11821 138879 11852
rect 142816 11852 143816 11880
rect 138836 11815 138894 11821
rect 137986 11784 138796 11812
rect 136450 11704 136456 11756
rect 136508 11753 136514 11756
rect 136508 11744 136520 11753
rect 136508 11716 136956 11744
rect 136508 11707 136520 11716
rect 136508 11704 136514 11707
rect 136726 11676 136732 11688
rect 135036 11648 135576 11676
rect 136687 11648 136732 11676
rect 135036 11636 135042 11648
rect 136726 11636 136732 11648
rect 136784 11636 136790 11688
rect 136928 11676 136956 11716
rect 137002 11704 137008 11756
rect 137060 11744 137066 11756
rect 138658 11744 138664 11756
rect 137060 11716 138664 11744
rect 137060 11704 137066 11716
rect 138658 11704 138664 11716
rect 138716 11704 138722 11756
rect 138768 11744 138796 11784
rect 138836 11781 138848 11815
rect 138882 11781 138894 11815
rect 142648 11815 142706 11821
rect 138836 11775 138894 11781
rect 138952 11784 141648 11812
rect 138952 11744 138980 11784
rect 138768 11716 138980 11744
rect 139118 11704 139124 11756
rect 139176 11744 139182 11756
rect 140685 11747 140743 11753
rect 140685 11744 140697 11747
rect 139176 11716 140697 11744
rect 139176 11704 139182 11716
rect 140685 11713 140697 11716
rect 140731 11713 140743 11747
rect 140685 11707 140743 11713
rect 137189 11679 137247 11685
rect 137189 11676 137201 11679
rect 136928 11648 137201 11676
rect 137189 11645 137201 11648
rect 137235 11645 137247 11679
rect 137189 11639 137247 11645
rect 135714 11608 135720 11620
rect 134904 11580 135720 11608
rect 135714 11568 135720 11580
rect 135772 11568 135778 11620
rect 137204 11608 137232 11639
rect 138198 11636 138204 11688
rect 138256 11676 138262 11688
rect 138569 11679 138627 11685
rect 138569 11676 138581 11679
rect 138256 11648 138581 11676
rect 138256 11636 138262 11648
rect 138569 11645 138581 11648
rect 138615 11645 138627 11679
rect 138569 11639 138627 11645
rect 140222 11636 140228 11688
rect 140280 11676 140286 11688
rect 140501 11679 140559 11685
rect 140501 11676 140513 11679
rect 140280 11648 140513 11676
rect 140280 11636 140286 11648
rect 140501 11645 140513 11648
rect 140547 11645 140559 11679
rect 141510 11676 141516 11688
rect 140501 11639 140559 11645
rect 140792 11648 141516 11676
rect 139946 11608 139952 11620
rect 137204 11580 138612 11608
rect 139907 11580 139952 11608
rect 125560 11512 127756 11540
rect 127805 11543 127863 11549
rect 125560 11500 125566 11512
rect 127805 11509 127817 11543
rect 127851 11540 127863 11543
rect 127894 11540 127900 11552
rect 127851 11512 127900 11540
rect 127851 11509 127863 11512
rect 127805 11503 127863 11509
rect 127894 11500 127900 11512
rect 127952 11500 127958 11552
rect 128446 11540 128452 11552
rect 128407 11512 128452 11540
rect 128446 11500 128452 11512
rect 128504 11500 128510 11552
rect 128722 11500 128728 11552
rect 128780 11540 128786 11552
rect 131393 11543 131451 11549
rect 131393 11540 131405 11543
rect 128780 11512 131405 11540
rect 128780 11500 128786 11512
rect 131393 11509 131405 11512
rect 131439 11540 131451 11543
rect 131850 11540 131856 11552
rect 131439 11512 131856 11540
rect 131439 11509 131451 11512
rect 131393 11503 131451 11509
rect 131850 11500 131856 11512
rect 131908 11500 131914 11552
rect 131945 11543 132003 11549
rect 131945 11509 131957 11543
rect 131991 11540 132003 11543
rect 132126 11540 132132 11552
rect 131991 11512 132132 11540
rect 131991 11509 132003 11512
rect 131945 11503 132003 11509
rect 132126 11500 132132 11512
rect 132184 11540 132190 11552
rect 132402 11540 132408 11552
rect 132184 11512 132408 11540
rect 132184 11500 132190 11512
rect 132402 11500 132408 11512
rect 132460 11500 132466 11552
rect 133046 11540 133052 11552
rect 133007 11512 133052 11540
rect 133046 11500 133052 11512
rect 133104 11500 133110 11552
rect 138109 11543 138167 11549
rect 138109 11509 138121 11543
rect 138155 11540 138167 11543
rect 138198 11540 138204 11552
rect 138155 11512 138204 11540
rect 138155 11509 138167 11512
rect 138109 11503 138167 11509
rect 138198 11500 138204 11512
rect 138256 11500 138262 11552
rect 138584 11540 138612 11580
rect 139946 11568 139952 11580
rect 140004 11568 140010 11620
rect 140792 11540 140820 11648
rect 141510 11636 141516 11648
rect 141568 11636 141574 11688
rect 138584 11512 140820 11540
rect 140869 11543 140927 11549
rect 140869 11509 140881 11543
rect 140915 11540 140927 11543
rect 141142 11540 141148 11552
rect 140915 11512 141148 11540
rect 140915 11509 140927 11512
rect 140869 11503 140927 11509
rect 141142 11500 141148 11512
rect 141200 11500 141206 11552
rect 141510 11540 141516 11552
rect 141471 11512 141516 11540
rect 141510 11500 141516 11512
rect 141568 11500 141574 11552
rect 141620 11540 141648 11784
rect 142648 11781 142660 11815
rect 142694 11812 142706 11815
rect 142816 11812 142844 11852
rect 143810 11840 143816 11852
rect 143868 11840 143874 11892
rect 143902 11840 143908 11892
rect 143960 11880 143966 11892
rect 148318 11880 148324 11892
rect 143960 11852 148324 11880
rect 143960 11840 143966 11852
rect 148318 11840 148324 11852
rect 148376 11840 148382 11892
rect 148686 11840 148692 11892
rect 148744 11880 148750 11892
rect 148744 11852 152504 11880
rect 148744 11840 148750 11852
rect 146386 11812 146392 11824
rect 142694 11784 142844 11812
rect 142908 11784 146392 11812
rect 142694 11781 142706 11784
rect 142648 11775 142706 11781
rect 142908 11688 142936 11784
rect 142982 11704 142988 11756
rect 143040 11744 143046 11756
rect 144178 11744 144184 11756
rect 143040 11716 144184 11744
rect 143040 11704 143046 11716
rect 144178 11704 144184 11716
rect 144236 11704 144242 11756
rect 144454 11704 144460 11756
rect 144512 11753 144518 11756
rect 144748 11753 144776 11784
rect 146386 11772 146392 11784
rect 146444 11812 146450 11824
rect 147582 11812 147588 11824
rect 146444 11784 147588 11812
rect 146444 11772 146450 11784
rect 144512 11744 144524 11753
rect 144733 11747 144791 11753
rect 144512 11716 144557 11744
rect 144512 11707 144524 11716
rect 144733 11713 144745 11747
rect 144779 11744 144791 11747
rect 144822 11744 144828 11756
rect 144779 11716 144828 11744
rect 144779 11713 144791 11716
rect 144733 11707 144791 11713
rect 144512 11704 144518 11707
rect 144822 11704 144828 11716
rect 144880 11704 144886 11756
rect 146777 11747 146835 11753
rect 146777 11713 146789 11747
rect 146823 11744 146835 11747
rect 146938 11744 146944 11756
rect 146823 11716 146944 11744
rect 146823 11713 146835 11716
rect 146777 11707 146835 11713
rect 146938 11704 146944 11716
rect 146996 11704 147002 11756
rect 147048 11753 147076 11784
rect 147582 11772 147588 11784
rect 147640 11812 147646 11824
rect 147640 11784 148916 11812
rect 147640 11772 147646 11784
rect 147033 11747 147091 11753
rect 147033 11713 147045 11747
rect 147079 11713 147091 11747
rect 148318 11744 148324 11756
rect 147033 11707 147091 11713
rect 147646 11716 148324 11744
rect 142890 11676 142896 11688
rect 142851 11648 142896 11676
rect 142890 11636 142896 11648
rect 142948 11636 142954 11688
rect 147122 11636 147128 11688
rect 147180 11676 147186 11688
rect 147490 11676 147496 11688
rect 147180 11648 147496 11676
rect 147180 11636 147186 11648
rect 147490 11636 147496 11648
rect 147548 11636 147554 11688
rect 147646 11608 147674 11716
rect 148318 11704 148324 11716
rect 148376 11704 148382 11756
rect 148888 11753 148916 11784
rect 150434 11772 150440 11824
rect 150492 11812 150498 11824
rect 151050 11815 151108 11821
rect 151050 11812 151062 11815
rect 150492 11784 151062 11812
rect 150492 11772 150498 11784
rect 151050 11781 151062 11784
rect 151096 11781 151108 11815
rect 152476 11812 152504 11852
rect 152550 11840 152556 11892
rect 152608 11880 152614 11892
rect 152645 11883 152703 11889
rect 152645 11880 152657 11883
rect 152608 11852 152657 11880
rect 152608 11840 152614 11852
rect 152645 11849 152657 11852
rect 152691 11849 152703 11883
rect 152645 11843 152703 11849
rect 153286 11840 153292 11892
rect 153344 11880 153350 11892
rect 156785 11883 156843 11889
rect 156785 11880 156797 11883
rect 153344 11852 156797 11880
rect 153344 11840 153350 11852
rect 156785 11849 156797 11852
rect 156831 11849 156843 11883
rect 157610 11880 157616 11892
rect 157571 11852 157616 11880
rect 156785 11843 156843 11849
rect 157610 11840 157616 11852
rect 157668 11840 157674 11892
rect 152476 11784 153424 11812
rect 151050 11775 151108 11781
rect 148617 11747 148675 11753
rect 148617 11713 148629 11747
rect 148663 11744 148675 11747
rect 148873 11747 148931 11753
rect 148663 11716 148824 11744
rect 148663 11713 148675 11716
rect 148617 11707 148675 11713
rect 148796 11676 148824 11716
rect 148873 11713 148885 11747
rect 148919 11713 148931 11747
rect 148873 11707 148931 11713
rect 149425 11747 149483 11753
rect 149425 11713 149437 11747
rect 149471 11744 149483 11747
rect 150158 11744 150164 11756
rect 149471 11716 150164 11744
rect 149471 11713 149483 11716
rect 149425 11707 149483 11713
rect 150158 11704 150164 11716
rect 150216 11704 150222 11756
rect 150253 11747 150311 11753
rect 150253 11713 150265 11747
rect 150299 11744 150311 11747
rect 153286 11744 153292 11756
rect 150299 11716 153292 11744
rect 150299 11713 150311 11716
rect 150253 11707 150311 11713
rect 153286 11704 153292 11716
rect 153344 11704 153350 11756
rect 153396 11744 153424 11784
rect 153672 11784 154068 11812
rect 153672 11744 153700 11784
rect 153396 11716 153700 11744
rect 153769 11747 153827 11753
rect 153769 11713 153781 11747
rect 153815 11744 153827 11747
rect 153930 11744 153936 11756
rect 153815 11716 153936 11744
rect 153815 11713 153827 11716
rect 153769 11707 153827 11713
rect 153930 11704 153936 11716
rect 153988 11704 153994 11756
rect 154040 11744 154068 11784
rect 154206 11772 154212 11824
rect 154264 11812 154270 11824
rect 155310 11812 155316 11824
rect 154264 11784 155316 11812
rect 154264 11772 154270 11784
rect 155310 11772 155316 11784
rect 155368 11772 155374 11824
rect 155678 11772 155684 11824
rect 155736 11812 155742 11824
rect 155736 11784 157840 11812
rect 155736 11772 155742 11784
rect 154574 11744 154580 11756
rect 154040 11716 154580 11744
rect 154574 11704 154580 11716
rect 154632 11704 154638 11756
rect 154666 11704 154672 11756
rect 154724 11744 154730 11756
rect 154724 11716 154769 11744
rect 154724 11704 154730 11716
rect 156138 11704 156144 11756
rect 156196 11742 156202 11756
rect 157812 11753 157840 11784
rect 156969 11747 157027 11753
rect 156196 11714 156239 11742
rect 156196 11704 156202 11714
rect 156969 11713 156981 11747
rect 157015 11713 157027 11747
rect 156969 11707 157027 11713
rect 157797 11747 157855 11753
rect 157797 11713 157809 11747
rect 157843 11713 157855 11747
rect 157797 11707 157855 11713
rect 150342 11676 150348 11688
rect 148796 11648 150348 11676
rect 150342 11636 150348 11648
rect 150400 11636 150406 11688
rect 150802 11676 150808 11688
rect 150763 11648 150808 11676
rect 150802 11636 150808 11648
rect 150860 11636 150866 11688
rect 154025 11679 154083 11685
rect 154025 11645 154037 11679
rect 154071 11676 154083 11679
rect 154298 11676 154304 11688
rect 154071 11648 154304 11676
rect 154071 11645 154083 11648
rect 154025 11639 154083 11645
rect 154298 11636 154304 11648
rect 154356 11636 154362 11688
rect 154390 11636 154396 11688
rect 154448 11676 154454 11688
rect 154485 11679 154543 11685
rect 154485 11676 154497 11679
rect 154448 11648 154497 11676
rect 154448 11636 154454 11648
rect 154485 11645 154497 11648
rect 154531 11645 154543 11679
rect 154485 11639 154543 11645
rect 154853 11679 154911 11685
rect 154853 11645 154865 11679
rect 154899 11676 154911 11679
rect 155678 11676 155684 11688
rect 154899 11648 155684 11676
rect 154899 11645 154911 11648
rect 154853 11639 154911 11645
rect 155678 11636 155684 11648
rect 155736 11636 155742 11688
rect 155957 11679 156015 11685
rect 155957 11676 155969 11679
rect 155788 11648 155969 11676
rect 150069 11611 150127 11617
rect 150069 11608 150081 11611
rect 142908 11580 143488 11608
rect 142908 11540 142936 11580
rect 141620 11512 142936 11540
rect 143258 11500 143264 11552
rect 143316 11540 143322 11552
rect 143353 11543 143411 11549
rect 143353 11540 143365 11543
rect 143316 11512 143365 11540
rect 143316 11500 143322 11512
rect 143353 11509 143365 11512
rect 143399 11509 143411 11543
rect 143460 11540 143488 11580
rect 144748 11580 145788 11608
rect 144748 11540 144776 11580
rect 143460 11512 144776 11540
rect 143353 11503 143411 11509
rect 144914 11500 144920 11552
rect 144972 11540 144978 11552
rect 145650 11540 145656 11552
rect 144972 11512 145656 11540
rect 144972 11500 144978 11512
rect 145650 11500 145656 11512
rect 145708 11500 145714 11552
rect 145760 11540 145788 11580
rect 147048 11580 147674 11608
rect 148888 11580 150081 11608
rect 147048 11540 147076 11580
rect 147490 11540 147496 11552
rect 145760 11512 147076 11540
rect 147451 11512 147496 11540
rect 147490 11500 147496 11512
rect 147548 11500 147554 11552
rect 147582 11500 147588 11552
rect 147640 11540 147646 11552
rect 148134 11540 148140 11552
rect 147640 11512 148140 11540
rect 147640 11500 147646 11512
rect 148134 11500 148140 11512
rect 148192 11500 148198 11552
rect 148502 11500 148508 11552
rect 148560 11540 148566 11552
rect 148888 11540 148916 11580
rect 150069 11577 150081 11580
rect 150115 11577 150127 11611
rect 150069 11571 150127 11577
rect 150158 11568 150164 11620
rect 150216 11608 150222 11620
rect 150820 11608 150848 11636
rect 152366 11608 152372 11620
rect 150216 11580 150848 11608
rect 151740 11580 152372 11608
rect 150216 11568 150222 11580
rect 148560 11512 148916 11540
rect 149517 11543 149575 11549
rect 148560 11500 148566 11512
rect 149517 11509 149529 11543
rect 149563 11540 149575 11543
rect 149606 11540 149612 11552
rect 149563 11512 149612 11540
rect 149563 11509 149575 11512
rect 149517 11503 149575 11509
rect 149606 11500 149612 11512
rect 149664 11500 149670 11552
rect 149974 11500 149980 11552
rect 150032 11540 150038 11552
rect 151740 11540 151768 11580
rect 152366 11568 152372 11580
rect 152424 11568 152430 11620
rect 155494 11608 155500 11620
rect 154132 11580 154712 11608
rect 150032 11512 151768 11540
rect 152185 11543 152243 11549
rect 150032 11500 150038 11512
rect 152185 11509 152197 11543
rect 152231 11540 152243 11543
rect 154132 11540 154160 11580
rect 152231 11512 154160 11540
rect 154684 11540 154712 11580
rect 154868 11580 155500 11608
rect 154868 11540 154896 11580
rect 155494 11568 155500 11580
rect 155552 11568 155558 11620
rect 155310 11540 155316 11552
rect 154684 11512 154896 11540
rect 155271 11512 155316 11540
rect 152231 11509 152243 11512
rect 152185 11503 152243 11509
rect 155310 11500 155316 11512
rect 155368 11500 155374 11552
rect 155402 11500 155408 11552
rect 155460 11540 155466 11552
rect 155678 11540 155684 11552
rect 155460 11512 155684 11540
rect 155460 11500 155466 11512
rect 155678 11500 155684 11512
rect 155736 11540 155742 11552
rect 155788 11540 155816 11648
rect 155957 11645 155969 11648
rect 156003 11645 156015 11679
rect 156984 11676 157012 11707
rect 155957 11639 156015 11645
rect 156156 11648 157012 11676
rect 157153 11679 157211 11685
rect 156156 11620 156184 11648
rect 157153 11645 157165 11679
rect 157199 11645 157211 11679
rect 157153 11639 157211 11645
rect 156138 11568 156144 11620
rect 156196 11568 156202 11620
rect 157168 11608 157196 11639
rect 156248 11580 157196 11608
rect 155736 11512 155816 11540
rect 155736 11500 155742 11512
rect 155862 11500 155868 11552
rect 155920 11540 155926 11552
rect 156248 11540 156276 11580
rect 155920 11512 156276 11540
rect 156325 11543 156383 11549
rect 155920 11500 155926 11512
rect 156325 11509 156337 11543
rect 156371 11540 156383 11543
rect 156506 11540 156512 11552
rect 156371 11512 156512 11540
rect 156371 11509 156383 11512
rect 156325 11503 156383 11509
rect 156506 11500 156512 11512
rect 156564 11500 156570 11552
rect 158254 11540 158260 11552
rect 158215 11512 158260 11540
rect 158254 11500 158260 11512
rect 158312 11500 158318 11552
rect 1104 11450 158884 11472
rect 1104 11398 20672 11450
rect 20724 11398 20736 11450
rect 20788 11398 20800 11450
rect 20852 11398 20864 11450
rect 20916 11398 20928 11450
rect 20980 11398 60117 11450
rect 60169 11398 60181 11450
rect 60233 11398 60245 11450
rect 60297 11398 60309 11450
rect 60361 11398 60373 11450
rect 60425 11398 99562 11450
rect 99614 11398 99626 11450
rect 99678 11398 99690 11450
rect 99742 11398 99754 11450
rect 99806 11398 99818 11450
rect 99870 11398 139007 11450
rect 139059 11398 139071 11450
rect 139123 11398 139135 11450
rect 139187 11398 139199 11450
rect 139251 11398 139263 11450
rect 139315 11398 158884 11450
rect 1104 11376 158884 11398
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 11238 11336 11244 11348
rect 10183 11308 11244 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 13630 11336 13636 11348
rect 11808 11308 13636 11336
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 8444 11240 9229 11268
rect 8444 11228 8450 11240
rect 9217 11237 9229 11240
rect 9263 11268 9275 11271
rect 11808 11268 11836 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 25590 11336 25596 11348
rect 13771 11308 25596 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 26145 11339 26203 11345
rect 26145 11305 26157 11339
rect 26191 11336 26203 11339
rect 28166 11336 28172 11348
rect 26191 11308 28172 11336
rect 26191 11305 26203 11308
rect 26145 11299 26203 11305
rect 28166 11296 28172 11308
rect 28224 11296 28230 11348
rect 30926 11336 30932 11348
rect 28276 11308 30932 11336
rect 9263 11240 11836 11268
rect 11885 11271 11943 11277
rect 9263 11237 9275 11240
rect 9217 11231 9275 11237
rect 11885 11237 11897 11271
rect 11931 11237 11943 11271
rect 17586 11268 17592 11280
rect 17547 11240 17592 11268
rect 11885 11231 11943 11237
rect 4890 11200 4896 11212
rect 4632 11172 4896 11200
rect 4632 11141 4660 11172
rect 4890 11160 4896 11172
rect 4948 11200 4954 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4948 11172 5365 11200
rect 4948 11160 4954 11172
rect 5353 11169 5365 11172
rect 5399 11200 5411 11203
rect 10502 11200 10508 11212
rect 5399 11172 10508 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 10686 11200 10692 11212
rect 10647 11172 10692 11200
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11900 11200 11928 11231
rect 17586 11228 17592 11240
rect 17644 11228 17650 11280
rect 23017 11271 23075 11277
rect 23017 11237 23029 11271
rect 23063 11268 23075 11271
rect 28276 11268 28304 11308
rect 30926 11296 30932 11308
rect 30984 11296 30990 11348
rect 31113 11339 31171 11345
rect 31113 11305 31125 11339
rect 31159 11336 31171 11339
rect 31386 11336 31392 11348
rect 31159 11308 31392 11336
rect 31159 11305 31171 11308
rect 31113 11299 31171 11305
rect 31386 11296 31392 11308
rect 31444 11296 31450 11348
rect 33045 11339 33103 11345
rect 31496 11308 32996 11336
rect 23063 11240 28304 11268
rect 23063 11237 23075 11240
rect 23017 11231 23075 11237
rect 30742 11228 30748 11280
rect 30800 11268 30806 11280
rect 31496 11268 31524 11308
rect 30800 11240 31524 11268
rect 32968 11268 32996 11308
rect 33045 11305 33057 11339
rect 33091 11336 33103 11339
rect 36170 11336 36176 11348
rect 33091 11308 36176 11336
rect 33091 11305 33103 11308
rect 33045 11299 33103 11305
rect 36170 11296 36176 11308
rect 36228 11296 36234 11348
rect 36265 11339 36323 11345
rect 36265 11305 36277 11339
rect 36311 11336 36323 11339
rect 36722 11336 36728 11348
rect 36311 11308 36728 11336
rect 36311 11305 36323 11308
rect 36265 11299 36323 11305
rect 36722 11296 36728 11308
rect 36780 11296 36786 11348
rect 37826 11296 37832 11348
rect 37884 11336 37890 11348
rect 38749 11339 38807 11345
rect 38749 11336 38761 11339
rect 37884 11308 38761 11336
rect 37884 11296 37890 11308
rect 38749 11305 38761 11308
rect 38795 11336 38807 11339
rect 40034 11336 40040 11348
rect 38795 11308 40040 11336
rect 38795 11305 38807 11308
rect 38749 11299 38807 11305
rect 40034 11296 40040 11308
rect 40092 11296 40098 11348
rect 40681 11339 40739 11345
rect 40681 11305 40693 11339
rect 40727 11336 40739 11339
rect 40770 11336 40776 11348
rect 40727 11308 40776 11336
rect 40727 11305 40739 11308
rect 40681 11299 40739 11305
rect 40770 11296 40776 11308
rect 40828 11296 40834 11348
rect 41969 11339 42027 11345
rect 41969 11305 41981 11339
rect 42015 11336 42027 11339
rect 42613 11339 42671 11345
rect 42015 11308 42564 11336
rect 42015 11305 42027 11308
rect 41969 11299 42027 11305
rect 34882 11268 34888 11280
rect 32968 11240 34888 11268
rect 30800 11228 30806 11240
rect 34882 11228 34888 11240
rect 34940 11228 34946 11280
rect 38289 11271 38347 11277
rect 38289 11237 38301 11271
rect 38335 11268 38347 11271
rect 38562 11268 38568 11280
rect 38335 11240 38568 11268
rect 38335 11237 38347 11240
rect 38289 11231 38347 11237
rect 38562 11228 38568 11240
rect 38620 11268 38626 11280
rect 39485 11271 39543 11277
rect 38620 11240 39436 11268
rect 38620 11228 38626 11240
rect 16206 11200 16212 11212
rect 11900 11172 12480 11200
rect 16167 11172 16212 11200
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 4847 11104 5917 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5905 11101 5917 11104
rect 5951 11132 5963 11135
rect 7742 11132 7748 11144
rect 5951 11104 7748 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 7742 11092 7748 11104
rect 7800 11132 7806 11144
rect 8202 11132 8208 11144
rect 7800 11104 8208 11132
rect 7800 11092 7806 11104
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10870 11132 10876 11144
rect 9640 11104 10876 11132
rect 9640 11092 9646 11104
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11132 11759 11135
rect 11882 11132 11888 11144
rect 11747 11104 11888 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12250 11132 12256 11144
rect 11992 11104 12256 11132
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11064 7987 11067
rect 11054 11064 11060 11076
rect 7975 11036 11060 11064
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11241 11067 11299 11073
rect 11241 11064 11253 11067
rect 11204 11036 11253 11064
rect 11204 11024 11210 11036
rect 11241 11033 11253 11036
rect 11287 11064 11299 11067
rect 11992 11064 12020 11104
rect 12250 11092 12256 11104
rect 12308 11132 12314 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12308 11104 12357 11132
rect 12308 11092 12314 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12452 11132 12480 11172
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 19426 11200 19432 11212
rect 17368 11172 18736 11200
rect 19387 11172 19432 11200
rect 17368 11160 17374 11172
rect 14369 11135 14427 11141
rect 12452 11104 12756 11132
rect 12345 11095 12403 11101
rect 12590 11067 12648 11073
rect 12590 11064 12602 11067
rect 11287 11036 12020 11064
rect 12084 11036 12602 11064
rect 11287 11033 11299 11036
rect 11241 11027 11299 11033
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 12084 10996 12112 11036
rect 12590 11033 12602 11036
rect 12636 11033 12648 11067
rect 12728 11064 12756 11104
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 15194 11132 15200 11144
rect 14415 11104 15200 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 15194 11092 15200 11104
rect 15252 11132 15258 11144
rect 16224 11132 16252 11160
rect 15252 11104 16252 11132
rect 16476 11135 16534 11141
rect 15252 11092 15258 11104
rect 16476 11101 16488 11135
rect 16522 11132 16534 11135
rect 18414 11132 18420 11144
rect 16522 11104 18420 11132
rect 16522 11101 16534 11104
rect 16476 11095 16534 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18598 11132 18604 11144
rect 18559 11104 18604 11132
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 18708 11132 18736 11172
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 20588 11172 21772 11200
rect 20588 11160 20594 11172
rect 21082 11132 21088 11144
rect 18708 11104 21088 11132
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11101 21695 11135
rect 21744 11132 21772 11172
rect 24394 11160 24400 11212
rect 24452 11200 24458 11212
rect 28537 11203 28595 11209
rect 28537 11200 28549 11203
rect 24452 11172 28549 11200
rect 24452 11160 24458 11172
rect 28537 11169 28549 11172
rect 28583 11200 28595 11203
rect 29546 11200 29552 11212
rect 28583 11172 29552 11200
rect 28583 11169 28595 11172
rect 28537 11163 28595 11169
rect 29546 11160 29552 11172
rect 29604 11160 29610 11212
rect 30852 11172 31800 11200
rect 23937 11135 23995 11141
rect 23937 11132 23949 11135
rect 21744 11104 23949 11132
rect 21637 11095 21695 11101
rect 23937 11101 23949 11104
rect 23983 11132 23995 11135
rect 24578 11132 24584 11144
rect 23983 11104 24584 11132
rect 23983 11101 23995 11104
rect 23937 11095 23995 11101
rect 14614 11067 14672 11073
rect 14614 11064 14626 11067
rect 12728 11036 14626 11064
rect 12590 11027 12648 11033
rect 14614 11033 14626 11036
rect 14660 11033 14672 11067
rect 18322 11064 18328 11076
rect 14614 11027 14672 11033
rect 15764 11036 18328 11064
rect 11480 10968 12112 10996
rect 11480 10956 11486 10968
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 15764 11005 15792 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 20254 11064 20260 11076
rect 18564 11036 20260 11064
rect 18564 11024 18570 11036
rect 20254 11024 20260 11036
rect 20312 11024 20318 11076
rect 21177 11067 21235 11073
rect 21177 11033 21189 11067
rect 21223 11064 21235 11067
rect 21358 11064 21364 11076
rect 21223 11036 21364 11064
rect 21223 11033 21235 11036
rect 21177 11027 21235 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 15749 10999 15807 11005
rect 15749 10996 15761 10999
rect 13688 10968 15761 10996
rect 13688 10956 13694 10968
rect 15749 10965 15761 10968
rect 15795 10965 15807 10999
rect 18414 10996 18420 11008
rect 18375 10968 18420 10996
rect 15749 10959 15807 10965
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 21652 10996 21680 11095
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 26602 11132 26608 11144
rect 24688 11104 26372 11132
rect 26563 11104 26608 11132
rect 21910 11073 21916 11076
rect 21904 11027 21916 11073
rect 21968 11064 21974 11076
rect 21968 11036 22004 11064
rect 21910 11024 21916 11027
rect 21968 11024 21974 11036
rect 22094 11024 22100 11076
rect 22152 11064 22158 11076
rect 24688 11064 24716 11104
rect 25130 11064 25136 11076
rect 22152 11036 24716 11064
rect 25091 11036 25136 11064
rect 22152 11024 22158 11036
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25317 11067 25375 11073
rect 25317 11033 25329 11067
rect 25363 11064 25375 11067
rect 26234 11064 26240 11076
rect 25363 11036 26240 11064
rect 25363 11033 25375 11036
rect 25317 11027 25375 11033
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 26344 11064 26372 11104
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 26789 11135 26847 11141
rect 26789 11101 26801 11135
rect 26835 11132 26847 11135
rect 27706 11132 27712 11144
rect 26835 11104 27712 11132
rect 26835 11101 26847 11104
rect 26789 11095 26847 11101
rect 27706 11092 27712 11104
rect 27764 11092 27770 11144
rect 29638 11092 29644 11144
rect 29696 11132 29702 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29696 11104 29745 11132
rect 29696 11092 29702 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 30000 11135 30058 11141
rect 30000 11101 30012 11135
rect 30046 11132 30058 11135
rect 30852 11132 30880 11172
rect 31772 11144 31800 11172
rect 33594 11160 33600 11212
rect 33652 11200 33658 11212
rect 34241 11203 34299 11209
rect 34241 11200 34253 11203
rect 33652 11172 34253 11200
rect 33652 11160 33658 11172
rect 34241 11169 34253 11172
rect 34287 11200 34299 11203
rect 34330 11200 34336 11212
rect 34287 11172 34336 11200
rect 34287 11169 34299 11172
rect 34241 11163 34299 11169
rect 34330 11160 34336 11172
rect 34388 11160 34394 11212
rect 39408 11200 39436 11240
rect 39485 11237 39497 11271
rect 39531 11268 39543 11271
rect 42242 11268 42248 11280
rect 39531 11240 42248 11268
rect 39531 11237 39543 11240
rect 39485 11231 39543 11237
rect 42242 11228 42248 11240
rect 42300 11228 42306 11280
rect 42536 11268 42564 11308
rect 42613 11305 42625 11339
rect 42659 11336 42671 11339
rect 43254 11336 43260 11348
rect 42659 11308 43260 11336
rect 42659 11305 42671 11308
rect 42613 11299 42671 11305
rect 43254 11296 43260 11308
rect 43312 11296 43318 11348
rect 44637 11339 44695 11345
rect 44637 11305 44649 11339
rect 44683 11336 44695 11339
rect 51626 11336 51632 11348
rect 44683 11308 51632 11336
rect 44683 11305 44695 11308
rect 44637 11299 44695 11305
rect 51626 11296 51632 11308
rect 51684 11296 51690 11348
rect 53466 11296 53472 11348
rect 53524 11336 53530 11348
rect 53561 11339 53619 11345
rect 53561 11336 53573 11339
rect 53524 11308 53573 11336
rect 53524 11296 53530 11308
rect 53561 11305 53573 11308
rect 53607 11305 53619 11339
rect 57885 11339 57943 11345
rect 53561 11299 53619 11305
rect 54036 11308 57836 11336
rect 42702 11268 42708 11280
rect 42536 11240 42708 11268
rect 42702 11228 42708 11240
rect 42760 11228 42766 11280
rect 45370 11268 45376 11280
rect 45331 11240 45376 11268
rect 45370 11228 45376 11240
rect 45428 11228 45434 11280
rect 45646 11228 45652 11280
rect 45704 11268 45710 11280
rect 47581 11271 47639 11277
rect 45704 11240 46244 11268
rect 45704 11228 45710 11240
rect 41230 11200 41236 11212
rect 36924 11172 39252 11200
rect 39408 11172 41236 11200
rect 31662 11132 31668 11144
rect 30046 11104 30880 11132
rect 31623 11104 31668 11132
rect 30046 11101 30058 11104
rect 30000 11095 30058 11101
rect 26878 11064 26884 11076
rect 26344 11036 26884 11064
rect 26878 11024 26884 11036
rect 26936 11024 26942 11076
rect 26973 11067 27031 11073
rect 26973 11033 26985 11067
rect 27019 11064 27031 11067
rect 27154 11064 27160 11076
rect 27019 11036 27160 11064
rect 27019 11033 27031 11036
rect 26973 11027 27031 11033
rect 27154 11024 27160 11036
rect 27212 11024 27218 11076
rect 27338 11024 27344 11076
rect 27396 11064 27402 11076
rect 29748 11064 29776 11095
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 31754 11092 31760 11144
rect 31812 11092 31818 11144
rect 33689 11135 33747 11141
rect 33689 11132 33701 11135
rect 31864 11104 33701 11132
rect 29914 11064 29920 11076
rect 27396 11036 27752 11064
rect 27396 11024 27402 11036
rect 22002 10996 22008 11008
rect 18656 10968 22008 10996
rect 18656 10956 18662 10968
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 27617 10999 27675 11005
rect 27617 10996 27629 10999
rect 27304 10968 27629 10996
rect 27304 10956 27310 10968
rect 27617 10965 27629 10968
rect 27663 10965 27675 10999
rect 27724 10996 27752 11036
rect 28920 11036 29224 11064
rect 29748 11036 29920 11064
rect 28920 10996 28948 11036
rect 29086 10996 29092 11008
rect 27724 10968 28948 10996
rect 29047 10968 29092 10996
rect 27617 10959 27675 10965
rect 29086 10956 29092 10968
rect 29144 10956 29150 11008
rect 29196 10996 29224 11036
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 31110 11024 31116 11076
rect 31168 11064 31174 11076
rect 31864 11064 31892 11104
rect 33689 11101 33701 11104
rect 33735 11101 33747 11135
rect 33689 11095 33747 11101
rect 34054 11092 34060 11144
rect 34112 11132 34118 11144
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34112 11104 34897 11132
rect 34112 11092 34118 11104
rect 34885 11101 34897 11104
rect 34931 11132 34943 11135
rect 34974 11132 34980 11144
rect 34931 11104 34980 11132
rect 34931 11101 34943 11104
rect 34885 11095 34943 11101
rect 34974 11092 34980 11104
rect 35032 11092 35038 11144
rect 36924 11141 36952 11172
rect 35152 11135 35210 11141
rect 35152 11101 35164 11135
rect 35198 11132 35210 11135
rect 36909 11135 36967 11141
rect 35198 11104 36860 11132
rect 35198 11101 35210 11104
rect 35152 11095 35210 11101
rect 31168 11036 31892 11064
rect 31932 11067 31990 11073
rect 31168 11024 31174 11036
rect 31932 11033 31944 11067
rect 31978 11064 31990 11067
rect 35894 11064 35900 11076
rect 31978 11036 35900 11064
rect 31978 11033 31990 11036
rect 31932 11027 31990 11033
rect 35894 11024 35900 11036
rect 35952 11024 35958 11076
rect 35986 11024 35992 11076
rect 36044 11064 36050 11076
rect 36725 11067 36783 11073
rect 36725 11064 36737 11067
rect 36044 11036 36737 11064
rect 36044 11024 36050 11036
rect 36725 11033 36737 11036
rect 36771 11033 36783 11067
rect 36832 11064 36860 11104
rect 36909 11101 36921 11135
rect 36955 11101 36967 11135
rect 36909 11095 36967 11101
rect 37093 11135 37151 11141
rect 37093 11101 37105 11135
rect 37139 11132 37151 11135
rect 37734 11132 37740 11144
rect 37139 11104 37740 11132
rect 37139 11101 37151 11104
rect 37093 11095 37151 11101
rect 37734 11092 37740 11104
rect 37792 11092 37798 11144
rect 37550 11064 37556 11076
rect 36832 11036 37556 11064
rect 36725 11027 36783 11033
rect 37550 11024 37556 11036
rect 37608 11024 37614 11076
rect 37645 11067 37703 11073
rect 37645 11033 37657 11067
rect 37691 11064 37703 11067
rect 39114 11064 39120 11076
rect 37691 11036 39120 11064
rect 37691 11033 37703 11036
rect 37645 11027 37703 11033
rect 31202 10996 31208 11008
rect 29196 10968 31208 10996
rect 31202 10956 31208 10968
rect 31260 10956 31266 11008
rect 31478 10956 31484 11008
rect 31536 10996 31542 11008
rect 33318 10996 33324 11008
rect 31536 10968 33324 10996
rect 31536 10956 31542 10968
rect 33318 10956 33324 10968
rect 33376 10956 33382 11008
rect 33502 10996 33508 11008
rect 33463 10968 33508 10996
rect 33502 10956 33508 10968
rect 33560 10956 33566 11008
rect 33778 10956 33784 11008
rect 33836 10996 33842 11008
rect 37660 10996 37688 11027
rect 39114 11024 39120 11036
rect 39172 11024 39178 11076
rect 39224 11064 39252 11172
rect 41230 11160 41236 11172
rect 41288 11160 41294 11212
rect 41322 11160 41328 11212
rect 41380 11200 41386 11212
rect 42518 11200 42524 11212
rect 41380 11172 42524 11200
rect 41380 11160 41386 11172
rect 42518 11160 42524 11172
rect 42576 11160 42582 11212
rect 45664 11200 45692 11228
rect 42720 11172 43300 11200
rect 39301 11135 39359 11141
rect 39301 11101 39313 11135
rect 39347 11132 39359 11135
rect 40218 11132 40224 11144
rect 39347 11104 40224 11132
rect 39347 11101 39359 11104
rect 39301 11095 39359 11101
rect 40218 11092 40224 11104
rect 40276 11092 40282 11144
rect 40865 11135 40923 11141
rect 40865 11101 40877 11135
rect 40911 11132 40923 11135
rect 41414 11132 41420 11144
rect 40911 11104 41420 11132
rect 40911 11101 40923 11104
rect 40865 11095 40923 11101
rect 41414 11092 41420 11104
rect 41472 11092 41478 11144
rect 41782 11132 41788 11144
rect 41743 11104 41788 11132
rect 41782 11092 41788 11104
rect 41840 11092 41846 11144
rect 40126 11064 40132 11076
rect 39224 11036 39988 11064
rect 40087 11036 40132 11064
rect 37826 10996 37832 11008
rect 33836 10968 37832 10996
rect 33836 10956 33842 10968
rect 37826 10956 37832 10968
rect 37884 10956 37890 11008
rect 39960 10996 39988 11036
rect 40126 11024 40132 11036
rect 40184 11064 40190 11076
rect 42720 11064 42748 11172
rect 43272 11141 43300 11172
rect 44652 11172 45692 11200
rect 42797 11135 42855 11141
rect 42797 11101 42809 11135
rect 42843 11132 42855 11135
rect 43257 11135 43315 11141
rect 42843 11104 43208 11132
rect 42843 11101 42855 11104
rect 42797 11095 42855 11101
rect 40184 11036 42748 11064
rect 40184 11024 40190 11036
rect 40770 10996 40776 11008
rect 39960 10968 40776 10996
rect 40770 10956 40776 10968
rect 40828 10956 40834 11008
rect 41506 10956 41512 11008
rect 41564 10996 41570 11008
rect 42610 10996 42616 11008
rect 41564 10968 42616 10996
rect 41564 10956 41570 10968
rect 42610 10956 42616 10968
rect 42668 10956 42674 11008
rect 43180 10996 43208 11104
rect 43257 11101 43269 11135
rect 43303 11132 43315 11135
rect 44652 11132 44680 11172
rect 46216 11144 46244 11240
rect 47581 11237 47593 11271
rect 47627 11268 47639 11271
rect 48314 11268 48320 11280
rect 47627 11240 48320 11268
rect 47627 11237 47639 11240
rect 47581 11231 47639 11237
rect 48314 11228 48320 11240
rect 48372 11268 48378 11280
rect 48498 11268 48504 11280
rect 48372 11240 48504 11268
rect 48372 11228 48378 11240
rect 48498 11228 48504 11240
rect 48556 11228 48562 11280
rect 48590 11228 48596 11280
rect 48648 11268 48654 11280
rect 53101 11271 53159 11277
rect 48648 11240 49648 11268
rect 48648 11228 48654 11240
rect 47302 11160 47308 11212
rect 47360 11200 47366 11212
rect 49510 11200 49516 11212
rect 47360 11172 49516 11200
rect 47360 11160 47366 11172
rect 49510 11160 49516 11172
rect 49568 11160 49574 11212
rect 49620 11151 49648 11240
rect 53101 11237 53113 11271
rect 53147 11268 53159 11271
rect 54036 11268 54064 11308
rect 55398 11268 55404 11280
rect 53147 11240 54064 11268
rect 54956 11240 55404 11268
rect 53147 11237 53159 11240
rect 53101 11231 53159 11237
rect 49786 11160 49792 11212
rect 49844 11200 49850 11212
rect 51718 11200 51724 11212
rect 49844 11172 51724 11200
rect 49844 11160 49850 11172
rect 51718 11160 51724 11172
rect 51776 11160 51782 11212
rect 54956 11200 54984 11240
rect 55398 11228 55404 11240
rect 55456 11228 55462 11280
rect 56873 11271 56931 11277
rect 56873 11237 56885 11271
rect 56919 11237 56931 11271
rect 57808 11268 57836 11308
rect 57885 11305 57897 11339
rect 57931 11336 57943 11339
rect 59262 11336 59268 11348
rect 57931 11308 59268 11336
rect 57931 11305 57943 11308
rect 57885 11299 57943 11305
rect 59262 11296 59268 11308
rect 59320 11296 59326 11348
rect 59998 11336 60004 11348
rect 59959 11308 60004 11336
rect 59998 11296 60004 11308
rect 60056 11296 60062 11348
rect 62022 11296 62028 11348
rect 62080 11336 62086 11348
rect 62577 11339 62635 11345
rect 62577 11336 62589 11339
rect 62080 11308 62589 11336
rect 62080 11296 62086 11308
rect 62577 11305 62589 11308
rect 62623 11305 62635 11339
rect 62577 11299 62635 11305
rect 65889 11339 65947 11345
rect 65889 11305 65901 11339
rect 65935 11336 65947 11339
rect 68005 11339 68063 11345
rect 68005 11336 68017 11339
rect 65935 11308 68017 11336
rect 65935 11305 65947 11308
rect 65889 11299 65947 11305
rect 68005 11305 68017 11308
rect 68051 11336 68063 11339
rect 70210 11336 70216 11348
rect 68051 11308 70216 11336
rect 68051 11305 68063 11308
rect 68005 11299 68063 11305
rect 58802 11268 58808 11280
rect 57808 11240 58808 11268
rect 56873 11231 56931 11237
rect 56888 11200 56916 11231
rect 58802 11228 58808 11240
rect 58860 11228 58866 11280
rect 54864 11172 54984 11200
rect 55048 11172 55628 11200
rect 56888 11172 59860 11200
rect 49605 11145 49663 11151
rect 43303 11104 44680 11132
rect 45557 11135 45615 11141
rect 43303 11101 43315 11104
rect 43257 11095 43315 11101
rect 45557 11101 45569 11135
rect 45603 11132 45615 11135
rect 45646 11132 45652 11144
rect 45603 11104 45652 11132
rect 45603 11101 45615 11104
rect 45557 11095 45615 11101
rect 45646 11092 45652 11104
rect 45704 11092 45710 11144
rect 45738 11092 45744 11144
rect 45796 11132 45802 11144
rect 46198 11132 46204 11144
rect 45796 11104 45841 11132
rect 46159 11104 46204 11132
rect 45796 11092 45802 11104
rect 46198 11092 46204 11104
rect 46256 11092 46262 11144
rect 46290 11092 46296 11144
rect 46348 11132 46354 11144
rect 48590 11132 48596 11144
rect 46348 11104 48596 11132
rect 46348 11092 46354 11104
rect 48590 11092 48596 11104
rect 48648 11092 48654 11144
rect 48682 11092 48688 11144
rect 48740 11134 48746 11144
rect 48740 11132 48820 11134
rect 49142 11132 49148 11144
rect 48740 11104 49148 11132
rect 48740 11092 48746 11104
rect 49142 11092 49148 11104
rect 49200 11092 49206 11144
rect 49421 11135 49479 11141
rect 49421 11101 49433 11135
rect 49467 11101 49479 11135
rect 49605 11111 49617 11145
rect 49651 11111 49663 11145
rect 49605 11105 49663 11111
rect 50801 11135 50859 11141
rect 49421 11095 49479 11101
rect 50801 11101 50813 11135
rect 50847 11101 50859 11135
rect 50801 11095 50859 11101
rect 43346 11024 43352 11076
rect 43404 11064 43410 11076
rect 43502 11067 43560 11073
rect 43502 11064 43514 11067
rect 43404 11036 43514 11064
rect 43404 11024 43410 11036
rect 43502 11033 43514 11036
rect 43548 11033 43560 11067
rect 45462 11064 45468 11076
rect 43502 11027 43560 11033
rect 43640 11036 45468 11064
rect 43640 10996 43668 11036
rect 45462 11024 45468 11036
rect 45520 11024 45526 11076
rect 46468 11067 46526 11073
rect 46468 11033 46480 11067
rect 46514 11064 46526 11067
rect 46842 11064 46848 11076
rect 46514 11036 46848 11064
rect 46514 11033 46526 11036
rect 46468 11027 46526 11033
rect 46842 11024 46848 11036
rect 46900 11024 46906 11076
rect 48774 11064 48780 11076
rect 48516 11036 48780 11064
rect 43180 10968 43668 10996
rect 48406 10956 48412 11008
rect 48464 10996 48470 11008
rect 48516 11005 48544 11036
rect 48774 11024 48780 11036
rect 48832 11024 48838 11076
rect 49234 11024 49240 11076
rect 49292 11064 49298 11076
rect 49436 11064 49464 11095
rect 50816 11064 50844 11095
rect 50890 11092 50896 11144
rect 50948 11134 50954 11144
rect 50985 11135 51043 11141
rect 50985 11134 50997 11135
rect 50948 11106 50997 11134
rect 50948 11092 50954 11106
rect 50985 11101 50997 11106
rect 51031 11101 51043 11135
rect 54864 11132 54892 11172
rect 50985 11095 51043 11101
rect 51920 11104 54892 11132
rect 54941 11135 54999 11141
rect 51074 11064 51080 11076
rect 49292 11036 49464 11064
rect 49712 11036 50568 11064
rect 50816 11036 51080 11064
rect 49292 11024 49298 11036
rect 48501 10999 48559 11005
rect 48501 10996 48513 10999
rect 48464 10968 48513 10996
rect 48464 10956 48470 10968
rect 48501 10965 48513 10968
rect 48547 10965 48559 10999
rect 48501 10959 48559 10965
rect 48590 10956 48596 11008
rect 48648 10996 48654 11008
rect 49712 10996 49740 11036
rect 48648 10968 49740 10996
rect 49789 10999 49847 11005
rect 48648 10956 48654 10968
rect 49789 10965 49801 10999
rect 49835 10996 49847 10999
rect 50430 10996 50436 11008
rect 49835 10968 50436 10996
rect 49835 10965 49847 10968
rect 49789 10959 49847 10965
rect 50430 10956 50436 10968
rect 50488 10956 50494 11008
rect 50540 10996 50568 11036
rect 51074 11024 51080 11036
rect 51132 11024 51138 11076
rect 51169 11067 51227 11073
rect 51169 11033 51181 11067
rect 51215 11064 51227 11067
rect 51920 11064 51948 11104
rect 54941 11101 54953 11135
rect 54987 11132 54999 11135
rect 55048 11132 55076 11172
rect 55600 11144 55628 11172
rect 54987 11104 55076 11132
rect 54987 11101 54999 11104
rect 54941 11095 54999 11101
rect 55306 11092 55312 11144
rect 55364 11132 55370 11144
rect 55493 11135 55551 11141
rect 55493 11132 55505 11135
rect 55364 11104 55505 11132
rect 55364 11092 55370 11104
rect 55493 11101 55505 11104
rect 55539 11101 55551 11135
rect 55493 11095 55551 11101
rect 55582 11092 55588 11144
rect 55640 11092 55646 11144
rect 55760 11135 55818 11141
rect 55760 11101 55772 11135
rect 55806 11101 55818 11135
rect 57698 11132 57704 11144
rect 57659 11104 57704 11132
rect 55760 11095 55818 11101
rect 51215 11036 51948 11064
rect 51988 11067 52046 11073
rect 51215 11033 51227 11036
rect 51169 11027 51227 11033
rect 51988 11033 52000 11067
rect 52034 11064 52046 11067
rect 52546 11064 52552 11076
rect 52034 11036 52552 11064
rect 52034 11033 52046 11036
rect 51988 11027 52046 11033
rect 52546 11024 52552 11036
rect 52604 11024 52610 11076
rect 54674 11067 54732 11073
rect 54674 11064 54686 11067
rect 53852 11036 54686 11064
rect 53852 10996 53880 11036
rect 54674 11033 54686 11036
rect 54720 11033 54732 11067
rect 54674 11027 54732 11033
rect 55214 11024 55220 11076
rect 55272 11064 55278 11076
rect 55272 11036 55628 11064
rect 55272 11024 55278 11036
rect 50540 10968 53880 10996
rect 55600 10996 55628 11036
rect 55674 11024 55680 11076
rect 55732 11064 55738 11076
rect 55784 11064 55812 11095
rect 57698 11092 57704 11104
rect 57756 11092 57762 11144
rect 58158 11092 58164 11144
rect 58216 11132 58222 11144
rect 58437 11135 58495 11141
rect 58437 11132 58449 11135
rect 58216 11104 58449 11132
rect 58216 11092 58222 11104
rect 58437 11101 58449 11104
rect 58483 11101 58495 11135
rect 58618 11132 58624 11144
rect 58579 11104 58624 11132
rect 58437 11095 58495 11101
rect 58618 11092 58624 11104
rect 58676 11092 58682 11144
rect 58805 11135 58863 11141
rect 58805 11101 58817 11135
rect 58851 11132 58863 11135
rect 58986 11132 58992 11144
rect 58851 11104 58992 11132
rect 58851 11101 58863 11104
rect 58805 11095 58863 11101
rect 58986 11092 58992 11104
rect 59044 11092 59050 11144
rect 59832 11141 59860 11172
rect 62022 11160 62028 11212
rect 62080 11200 62086 11212
rect 62080 11172 64276 11200
rect 62080 11160 62086 11172
rect 59817 11135 59875 11141
rect 59817 11101 59829 11135
rect 59863 11101 59875 11135
rect 59817 11095 59875 11101
rect 60645 11135 60703 11141
rect 60645 11101 60657 11135
rect 60691 11132 60703 11135
rect 62114 11132 62120 11144
rect 60691 11104 62120 11132
rect 60691 11101 60703 11104
rect 60645 11095 60703 11101
rect 56134 11064 56140 11076
rect 55732 11036 55812 11064
rect 55876 11036 56140 11064
rect 55732 11024 55738 11036
rect 55876 10996 55904 11036
rect 56134 11024 56140 11036
rect 56192 11064 56198 11076
rect 60660 11064 60688 11095
rect 62114 11092 62120 11104
rect 62172 11092 62178 11144
rect 62758 11132 62764 11144
rect 62719 11104 62764 11132
rect 62758 11092 62764 11104
rect 62816 11092 62822 11144
rect 56192 11036 60688 11064
rect 60912 11067 60970 11073
rect 56192 11024 56198 11036
rect 60912 11033 60924 11067
rect 60958 11064 60970 11067
rect 63218 11064 63224 11076
rect 60958 11036 63224 11064
rect 60958 11033 60970 11036
rect 60912 11027 60970 11033
rect 63218 11024 63224 11036
rect 63276 11024 63282 11076
rect 64248 11064 64276 11172
rect 65242 11160 65248 11212
rect 65300 11200 65306 11212
rect 65904 11200 65932 11299
rect 70210 11296 70216 11308
rect 70268 11296 70274 11348
rect 70578 11296 70584 11348
rect 70636 11336 70642 11348
rect 81434 11336 81440 11348
rect 70636 11308 81440 11336
rect 70636 11296 70642 11308
rect 81434 11296 81440 11308
rect 81492 11296 81498 11348
rect 81526 11296 81532 11348
rect 81584 11336 81590 11348
rect 82449 11339 82507 11345
rect 82449 11336 82461 11339
rect 81584 11308 82461 11336
rect 81584 11296 81590 11308
rect 82449 11305 82461 11308
rect 82495 11305 82507 11339
rect 83550 11336 83556 11348
rect 82449 11299 82507 11305
rect 82556 11308 83556 11336
rect 66625 11271 66683 11277
rect 66625 11237 66637 11271
rect 66671 11237 66683 11271
rect 66625 11231 66683 11237
rect 65300 11172 65932 11200
rect 65300 11160 65306 11172
rect 64506 11092 64512 11144
rect 64564 11132 64570 11144
rect 66640 11132 66668 11231
rect 66714 11228 66720 11280
rect 66772 11268 66778 11280
rect 73249 11271 73307 11277
rect 66772 11240 69980 11268
rect 66772 11228 66778 11240
rect 66990 11160 66996 11212
rect 67048 11200 67054 11212
rect 69753 11203 69811 11209
rect 69753 11200 69765 11203
rect 67048 11172 69765 11200
rect 67048 11160 67054 11172
rect 69753 11169 69765 11172
rect 69799 11169 69811 11203
rect 69753 11163 69811 11169
rect 64564 11104 66668 11132
rect 66809 11135 66867 11141
rect 64564 11092 64570 11104
rect 66809 11101 66821 11135
rect 66855 11132 66867 11135
rect 68370 11132 68376 11144
rect 66855 11104 68376 11132
rect 66855 11101 66867 11104
rect 66809 11095 66867 11101
rect 68370 11092 68376 11104
rect 68428 11092 68434 11144
rect 68554 11092 68560 11144
rect 68612 11132 68618 11144
rect 69952 11141 69980 11240
rect 73249 11237 73261 11271
rect 73295 11268 73307 11271
rect 75638 11268 75644 11280
rect 73295 11240 75644 11268
rect 73295 11237 73307 11240
rect 73249 11231 73307 11237
rect 75638 11228 75644 11240
rect 75696 11228 75702 11280
rect 76561 11271 76619 11277
rect 76561 11237 76573 11271
rect 76607 11237 76619 11271
rect 76561 11231 76619 11237
rect 80701 11271 80759 11277
rect 80701 11237 80713 11271
rect 80747 11268 80759 11271
rect 81989 11271 82047 11277
rect 81989 11268 82001 11271
rect 80747 11240 82001 11268
rect 80747 11237 80759 11240
rect 80701 11231 80759 11237
rect 81989 11237 82001 11240
rect 82035 11268 82047 11271
rect 82556 11268 82584 11308
rect 83550 11296 83556 11308
rect 83608 11336 83614 11348
rect 87506 11336 87512 11348
rect 83608 11308 87512 11336
rect 83608 11296 83614 11308
rect 87506 11296 87512 11308
rect 87564 11296 87570 11348
rect 88521 11339 88579 11345
rect 88521 11305 88533 11339
rect 88567 11336 88579 11339
rect 107105 11339 107163 11345
rect 88567 11308 104756 11336
rect 88567 11305 88579 11308
rect 88521 11299 88579 11305
rect 82035 11240 82584 11268
rect 82035 11237 82047 11240
rect 81989 11231 82047 11237
rect 70302 11160 70308 11212
rect 70360 11200 70366 11212
rect 71409 11203 71467 11209
rect 71409 11200 71421 11203
rect 70360 11172 71421 11200
rect 70360 11160 70366 11172
rect 71409 11169 71421 11172
rect 71455 11200 71467 11203
rect 71866 11200 71872 11212
rect 71455 11172 71872 11200
rect 71455 11169 71467 11172
rect 71409 11163 71467 11169
rect 71866 11160 71872 11172
rect 71924 11160 71930 11212
rect 73614 11160 73620 11212
rect 73672 11200 73678 11212
rect 76576 11200 76604 11231
rect 84194 11228 84200 11280
rect 84252 11268 84258 11280
rect 86862 11268 86868 11280
rect 84252 11240 86868 11268
rect 84252 11228 84258 11240
rect 86862 11228 86868 11240
rect 86920 11228 86926 11280
rect 88702 11228 88708 11280
rect 88760 11268 88766 11280
rect 88981 11271 89039 11277
rect 88981 11268 88993 11271
rect 88760 11240 88993 11268
rect 88760 11228 88766 11240
rect 88981 11237 88993 11240
rect 89027 11237 89039 11271
rect 88981 11231 89039 11237
rect 90358 11228 90364 11280
rect 90416 11228 90422 11280
rect 90818 11268 90824 11280
rect 90779 11240 90824 11268
rect 90818 11228 90824 11240
rect 90876 11228 90882 11280
rect 92474 11268 92480 11280
rect 92435 11240 92480 11268
rect 92474 11228 92480 11240
rect 92532 11228 92538 11280
rect 94222 11228 94228 11280
rect 94280 11268 94286 11280
rect 95421 11271 95479 11277
rect 95421 11268 95433 11271
rect 94280 11240 95433 11268
rect 94280 11228 94286 11240
rect 95421 11237 95433 11240
rect 95467 11268 95479 11271
rect 95602 11268 95608 11280
rect 95467 11240 95608 11268
rect 95467 11237 95479 11240
rect 95421 11231 95479 11237
rect 95602 11228 95608 11240
rect 95660 11228 95666 11280
rect 96065 11271 96123 11277
rect 96065 11237 96077 11271
rect 96111 11268 96123 11271
rect 96430 11268 96436 11280
rect 96111 11240 96436 11268
rect 96111 11237 96123 11240
rect 96065 11231 96123 11237
rect 96430 11228 96436 11240
rect 96488 11228 96494 11280
rect 96798 11268 96804 11280
rect 96759 11240 96804 11268
rect 96798 11228 96804 11240
rect 96856 11228 96862 11280
rect 101674 11228 101680 11280
rect 101732 11268 101738 11280
rect 101953 11271 102011 11277
rect 101953 11268 101965 11271
rect 101732 11240 101965 11268
rect 101732 11228 101738 11240
rect 101953 11237 101965 11240
rect 101999 11237 102011 11271
rect 104728 11268 104756 11308
rect 107105 11305 107117 11339
rect 107151 11336 107163 11339
rect 107470 11336 107476 11348
rect 107151 11308 107476 11336
rect 107151 11305 107163 11308
rect 107105 11299 107163 11305
rect 107470 11296 107476 11308
rect 107528 11296 107534 11348
rect 107562 11296 107568 11348
rect 107620 11336 107626 11348
rect 107657 11339 107715 11345
rect 107657 11336 107669 11339
rect 107620 11308 107669 11336
rect 107620 11296 107626 11308
rect 107657 11305 107669 11308
rect 107703 11305 107715 11339
rect 108758 11336 108764 11348
rect 108719 11308 108764 11336
rect 107657 11299 107715 11305
rect 108758 11296 108764 11308
rect 108816 11296 108822 11348
rect 109586 11336 109592 11348
rect 109547 11308 109592 11336
rect 109586 11296 109592 11308
rect 109644 11296 109650 11348
rect 112070 11296 112076 11348
rect 112128 11336 112134 11348
rect 113818 11336 113824 11348
rect 112128 11308 113824 11336
rect 112128 11296 112134 11308
rect 113818 11296 113824 11308
rect 113876 11296 113882 11348
rect 114554 11296 114560 11348
rect 114612 11336 114618 11348
rect 115198 11336 115204 11348
rect 114612 11308 115204 11336
rect 114612 11296 114618 11308
rect 115198 11296 115204 11308
rect 115256 11296 115262 11348
rect 118418 11336 118424 11348
rect 115400 11308 118424 11336
rect 104728 11240 109034 11268
rect 101953 11231 102011 11237
rect 77938 11200 77944 11212
rect 73672 11172 76604 11200
rect 77899 11172 77944 11200
rect 73672 11160 73678 11172
rect 77938 11160 77944 11172
rect 77996 11200 78002 11212
rect 79321 11203 79379 11209
rect 79321 11200 79333 11203
rect 77996 11172 79333 11200
rect 77996 11160 78002 11172
rect 79321 11169 79333 11172
rect 79367 11169 79379 11203
rect 86678 11200 86684 11212
rect 79321 11163 79379 11169
rect 83752 11172 84056 11200
rect 69937 11135 69995 11141
rect 68612 11104 69520 11132
rect 68612 11092 68618 11104
rect 64248 11036 64736 11064
rect 55600 10968 55904 10996
rect 55950 10956 55956 11008
rect 56008 10996 56014 11008
rect 56686 10996 56692 11008
rect 56008 10968 56692 10996
rect 56008 10956 56014 10968
rect 56686 10956 56692 10968
rect 56744 10996 56750 11008
rect 59265 10999 59323 11005
rect 59265 10996 59277 10999
rect 56744 10968 59277 10996
rect 56744 10956 56750 10968
rect 59265 10965 59277 10968
rect 59311 10996 59323 10999
rect 61010 10996 61016 11008
rect 59311 10968 61016 10996
rect 59311 10965 59323 10968
rect 59265 10959 59323 10965
rect 61010 10956 61016 10968
rect 61068 10956 61074 11008
rect 62022 10996 62028 11008
rect 61983 10968 62028 10996
rect 62022 10956 62028 10968
rect 62080 10956 62086 11008
rect 63402 10996 63408 11008
rect 63363 10968 63408 10996
rect 63402 10956 63408 10968
rect 63460 10956 63466 11008
rect 63862 10996 63868 11008
rect 63823 10968 63868 10996
rect 63862 10956 63868 10968
rect 63920 10956 63926 11008
rect 64708 10996 64736 11036
rect 64782 11024 64788 11076
rect 64840 11064 64846 11076
rect 64978 11067 65036 11073
rect 64978 11064 64990 11067
rect 64840 11036 64990 11064
rect 64840 11024 64846 11036
rect 64978 11033 64990 11036
rect 65024 11033 65036 11067
rect 66714 11064 66720 11076
rect 64978 11027 65036 11033
rect 65076 11036 66720 11064
rect 65076 10996 65104 11036
rect 66714 11024 66720 11036
rect 66772 11024 66778 11076
rect 69290 11064 69296 11076
rect 69251 11036 69296 11064
rect 69290 11024 69296 11036
rect 69348 11024 69354 11076
rect 69492 11064 69520 11104
rect 69937 11101 69949 11135
rect 69983 11101 69995 11135
rect 69937 11095 69995 11101
rect 70026 11092 70032 11144
rect 70084 11132 70090 11144
rect 72136 11135 72194 11141
rect 70084 11104 70129 11132
rect 70084 11092 70090 11104
rect 72136 11101 72148 11135
rect 72182 11132 72194 11135
rect 72970 11132 72976 11144
rect 72182 11104 72976 11132
rect 72182 11101 72194 11104
rect 72136 11095 72194 11101
rect 72970 11092 72976 11104
rect 73028 11092 73034 11144
rect 75270 11132 75276 11144
rect 75231 11104 75276 11132
rect 75270 11092 75276 11104
rect 75328 11092 75334 11144
rect 76742 11092 76748 11144
rect 76800 11132 76806 11144
rect 78858 11132 78864 11144
rect 76800 11104 78864 11132
rect 76800 11092 76806 11104
rect 78858 11092 78864 11104
rect 78916 11092 78922 11144
rect 79336 11132 79364 11163
rect 81253 11135 81311 11141
rect 81253 11132 81265 11135
rect 79336 11104 81265 11132
rect 81253 11101 81265 11104
rect 81299 11132 81311 11135
rect 83752 11132 83780 11172
rect 81299 11104 83780 11132
rect 83829 11135 83887 11141
rect 81299 11101 81311 11104
rect 81253 11095 81311 11101
rect 83829 11101 83841 11135
rect 83875 11132 83887 11135
rect 83918 11132 83924 11144
rect 83875 11104 83924 11132
rect 83875 11101 83887 11104
rect 83829 11095 83887 11101
rect 83918 11092 83924 11104
rect 83976 11092 83982 11144
rect 84028 11132 84056 11172
rect 84672 11172 86684 11200
rect 84672 11132 84700 11172
rect 86678 11160 86684 11172
rect 86736 11200 86742 11212
rect 87141 11203 87199 11209
rect 87141 11200 87153 11203
rect 86736 11172 87153 11200
rect 86736 11160 86742 11172
rect 87141 11169 87153 11172
rect 87187 11169 87199 11203
rect 90376 11200 90404 11228
rect 98178 11200 98184 11212
rect 90376 11172 90772 11200
rect 98139 11172 98184 11200
rect 87141 11163 87199 11169
rect 84028 11104 84700 11132
rect 84749 11135 84807 11141
rect 84749 11101 84761 11135
rect 84795 11132 84807 11135
rect 85853 11135 85911 11141
rect 85853 11132 85865 11135
rect 84795 11104 85865 11132
rect 84795 11101 84807 11104
rect 84749 11095 84807 11101
rect 85853 11101 85865 11104
rect 85899 11132 85911 11135
rect 86497 11135 86555 11141
rect 86497 11132 86509 11135
rect 85899 11104 86509 11132
rect 85899 11101 85911 11104
rect 85853 11095 85911 11101
rect 86497 11101 86509 11104
rect 86543 11132 86555 11135
rect 90266 11132 90272 11144
rect 86543 11104 90272 11132
rect 86543 11101 86555 11104
rect 86497 11095 86555 11101
rect 90266 11092 90272 11104
rect 90324 11092 90330 11144
rect 90361 11135 90419 11141
rect 90361 11101 90373 11135
rect 90407 11132 90419 11135
rect 90634 11132 90640 11144
rect 90407 11104 90640 11132
rect 90407 11101 90419 11104
rect 90361 11095 90419 11101
rect 90634 11092 90640 11104
rect 90692 11092 90698 11144
rect 90744 11132 90772 11172
rect 98178 11160 98184 11172
rect 98236 11200 98242 11212
rect 99285 11203 99343 11209
rect 99285 11200 99297 11203
rect 98236 11172 99297 11200
rect 98236 11160 98242 11172
rect 99285 11169 99297 11172
rect 99331 11200 99343 11203
rect 102226 11200 102232 11212
rect 99331 11172 102232 11200
rect 99331 11169 99343 11172
rect 99285 11163 99343 11169
rect 102226 11160 102232 11172
rect 102284 11160 102290 11212
rect 103790 11200 103796 11212
rect 103256 11172 103560 11200
rect 103751 11172 103796 11200
rect 90744 11104 93164 11132
rect 72326 11064 72332 11076
rect 69492 11036 72332 11064
rect 72326 11024 72332 11036
rect 72384 11024 72390 11076
rect 74626 11064 74632 11076
rect 74587 11036 74632 11064
rect 74626 11024 74632 11036
rect 74684 11024 74690 11076
rect 77294 11024 77300 11076
rect 77352 11064 77358 11076
rect 77674 11067 77732 11073
rect 77674 11064 77686 11067
rect 77352 11036 77686 11064
rect 77352 11024 77358 11036
rect 77674 11033 77686 11036
rect 77720 11033 77732 11067
rect 77674 11027 77732 11033
rect 79588 11067 79646 11073
rect 79588 11033 79600 11067
rect 79634 11064 79646 11067
rect 82814 11064 82820 11076
rect 79634 11036 82820 11064
rect 79634 11033 79646 11036
rect 79588 11027 79646 11033
rect 82814 11024 82820 11036
rect 82872 11024 82878 11076
rect 83550 11024 83556 11076
rect 83608 11073 83614 11076
rect 83608 11067 83642 11073
rect 83630 11033 83642 11067
rect 83608 11027 83642 11033
rect 83608 11024 83614 11027
rect 85022 11024 85028 11076
rect 85080 11064 85086 11076
rect 85485 11067 85543 11073
rect 85485 11064 85497 11067
rect 85080 11036 85497 11064
rect 85080 11024 85086 11036
rect 85485 11033 85497 11036
rect 85531 11033 85543 11067
rect 85485 11027 85543 11033
rect 87408 11067 87466 11073
rect 87408 11033 87420 11067
rect 87454 11064 87466 11067
rect 88518 11064 88524 11076
rect 87454 11036 88524 11064
rect 87454 11033 87466 11036
rect 87408 11027 87466 11033
rect 88518 11024 88524 11036
rect 88576 11024 88582 11076
rect 90116 11067 90174 11073
rect 90116 11033 90128 11067
rect 90162 11064 90174 11067
rect 91557 11067 91615 11073
rect 91557 11064 91569 11067
rect 90162 11036 91569 11064
rect 90162 11033 90174 11036
rect 90116 11027 90174 11033
rect 91557 11033 91569 11036
rect 91603 11064 91615 11067
rect 93026 11064 93032 11076
rect 91603 11036 93032 11064
rect 91603 11033 91615 11036
rect 91557 11027 91615 11033
rect 93026 11024 93032 11036
rect 93084 11024 93090 11076
rect 93136 11064 93164 11104
rect 93210 11092 93216 11144
rect 93268 11132 93274 11144
rect 93857 11135 93915 11141
rect 93857 11132 93869 11135
rect 93268 11104 93869 11132
rect 93268 11092 93274 11104
rect 93857 11101 93869 11104
rect 93903 11132 93915 11135
rect 94869 11135 94927 11141
rect 94869 11132 94881 11135
rect 93903 11104 94881 11132
rect 93903 11101 93915 11104
rect 93857 11095 93915 11101
rect 94869 11101 94881 11104
rect 94915 11101 94927 11135
rect 94869 11095 94927 11101
rect 98730 11092 98736 11144
rect 98788 11132 98794 11144
rect 98825 11135 98883 11141
rect 98825 11132 98837 11135
rect 98788 11104 98837 11132
rect 98788 11092 98794 11104
rect 98825 11101 98837 11104
rect 98871 11101 98883 11135
rect 98825 11095 98883 11101
rect 101398 11092 101404 11144
rect 101456 11132 101462 11144
rect 103256 11132 103284 11172
rect 101456 11104 103284 11132
rect 103333 11135 103391 11141
rect 101456 11092 101462 11104
rect 103333 11101 103345 11135
rect 103379 11132 103391 11135
rect 103422 11132 103428 11144
rect 103379 11104 103428 11132
rect 103379 11101 103391 11104
rect 103333 11095 103391 11101
rect 103422 11092 103428 11104
rect 103480 11092 103486 11144
rect 103532 11132 103560 11172
rect 103790 11160 103796 11172
rect 103848 11160 103854 11212
rect 106277 11203 106335 11209
rect 106277 11169 106289 11203
rect 106323 11200 106335 11203
rect 106458 11200 106464 11212
rect 106323 11172 106464 11200
rect 106323 11169 106335 11172
rect 106277 11163 106335 11169
rect 106458 11160 106464 11172
rect 106516 11200 106522 11212
rect 106642 11200 106648 11212
rect 106516 11172 106648 11200
rect 106516 11160 106522 11172
rect 106642 11160 106648 11172
rect 106700 11160 106706 11212
rect 109006 11200 109034 11240
rect 109218 11228 109224 11280
rect 109276 11268 109282 11280
rect 109276 11240 109632 11268
rect 109276 11228 109282 11240
rect 109006 11172 109264 11200
rect 105814 11132 105820 11144
rect 103532 11104 105820 11132
rect 105814 11092 105820 11104
rect 105872 11092 105878 11144
rect 106734 11132 106740 11144
rect 106292 11104 106740 11132
rect 93612 11067 93670 11073
rect 93136 11036 93532 11064
rect 64708 10968 65104 10996
rect 68922 10956 68928 11008
rect 68980 10996 68986 11008
rect 70026 10996 70032 11008
rect 68980 10968 70032 10996
rect 68980 10956 68986 10968
rect 70026 10956 70032 10968
rect 70084 10956 70090 11008
rect 74077 10999 74135 11005
rect 74077 10965 74089 10999
rect 74123 10996 74135 10999
rect 74350 10996 74356 11008
rect 74123 10968 74356 10996
rect 74123 10965 74135 10968
rect 74077 10959 74135 10965
rect 74350 10956 74356 10968
rect 74408 10956 74414 11008
rect 75454 10996 75460 11008
rect 75415 10968 75460 10996
rect 75454 10956 75460 10968
rect 75512 10956 75518 11008
rect 77110 10956 77116 11008
rect 77168 10996 77174 11008
rect 81250 10996 81256 11008
rect 77168 10968 81256 10996
rect 77168 10956 77174 10968
rect 81250 10956 81256 10968
rect 81308 10956 81314 11008
rect 81342 10956 81348 11008
rect 81400 10996 81406 11008
rect 84562 10996 84568 11008
rect 81400 10968 84568 10996
rect 81400 10956 81406 10968
rect 84562 10956 84568 10968
rect 84620 10956 84626 11008
rect 84746 10956 84752 11008
rect 84804 10996 84810 11008
rect 84841 10999 84899 11005
rect 84841 10996 84853 10999
rect 84804 10968 84853 10996
rect 84804 10956 84810 10968
rect 84841 10965 84853 10968
rect 84887 10965 84899 10999
rect 84841 10959 84899 10965
rect 84930 10956 84936 11008
rect 84988 10996 84994 11008
rect 89714 10996 89720 11008
rect 84988 10968 89720 10996
rect 84988 10956 84994 10968
rect 89714 10956 89720 10968
rect 89772 10956 89778 11008
rect 90634 10956 90640 11008
rect 90692 10996 90698 11008
rect 92014 10996 92020 11008
rect 90692 10968 92020 10996
rect 90692 10956 90698 10968
rect 92014 10956 92020 10968
rect 92072 10956 92078 11008
rect 93504 10996 93532 11036
rect 93612 11033 93624 11067
rect 93658 11064 93670 11067
rect 94406 11064 94412 11076
rect 93658 11036 94412 11064
rect 93658 11033 93670 11036
rect 93612 11027 93670 11033
rect 94406 11024 94412 11036
rect 94464 11024 94470 11076
rect 97936 11067 97994 11073
rect 97936 11033 97948 11067
rect 97982 11064 97994 11067
rect 98270 11064 98276 11076
rect 97982 11036 98276 11064
rect 97982 11033 97994 11036
rect 97936 11027 97994 11033
rect 98270 11024 98276 11036
rect 98328 11024 98334 11076
rect 99837 11067 99895 11073
rect 99837 11033 99849 11067
rect 99883 11033 99895 11067
rect 103088 11067 103146 11073
rect 99837 11027 99895 11033
rect 101876 11036 102088 11064
rect 94774 10996 94780 11008
rect 93504 10968 94780 10996
rect 94774 10956 94780 10968
rect 94832 10956 94838 11008
rect 98638 10996 98644 11008
rect 98599 10968 98644 10996
rect 98638 10956 98644 10968
rect 98696 10956 98702 11008
rect 98822 10956 98828 11008
rect 98880 10996 98886 11008
rect 99466 10996 99472 11008
rect 98880 10968 99472 10996
rect 98880 10956 98886 10968
rect 99466 10956 99472 10968
rect 99524 10996 99530 11008
rect 99852 10996 99880 11027
rect 99524 10968 99880 10996
rect 99524 10956 99530 10968
rect 101122 10956 101128 11008
rect 101180 10996 101186 11008
rect 101876 10996 101904 11036
rect 101180 10968 101904 10996
rect 102060 10996 102088 11036
rect 103088 11033 103100 11067
rect 103134 11064 103146 11067
rect 103514 11064 103520 11076
rect 103134 11036 103520 11064
rect 103134 11033 103146 11036
rect 103088 11027 103146 11033
rect 103514 11024 103520 11036
rect 103572 11024 103578 11076
rect 104060 11067 104118 11073
rect 104060 11033 104072 11067
rect 104106 11064 104118 11067
rect 105722 11064 105728 11076
rect 104106 11036 105584 11064
rect 105683 11036 105728 11064
rect 104106 11033 104118 11036
rect 104060 11027 104118 11033
rect 103330 10996 103336 11008
rect 102060 10968 103336 10996
rect 101180 10956 101186 10968
rect 103330 10956 103336 10968
rect 103388 10956 103394 11008
rect 105170 10996 105176 11008
rect 105131 10968 105176 10996
rect 105170 10956 105176 10968
rect 105228 10956 105234 11008
rect 105556 10996 105584 11036
rect 105722 11024 105728 11036
rect 105780 11024 105786 11076
rect 106292 11064 106320 11104
rect 106734 11092 106740 11104
rect 106792 11092 106798 11144
rect 108298 11132 108304 11144
rect 108259 11104 108304 11132
rect 108298 11092 108304 11104
rect 108356 11132 108362 11144
rect 108574 11132 108580 11144
rect 108356 11104 108580 11132
rect 108356 11092 108362 11104
rect 108574 11092 108580 11104
rect 108632 11092 108638 11144
rect 108945 11135 109003 11141
rect 108945 11101 108957 11135
rect 108991 11101 109003 11135
rect 109126 11132 109132 11144
rect 109087 11104 109132 11132
rect 108945 11095 109003 11101
rect 105832 11036 106320 11064
rect 105832 10996 105860 11036
rect 106366 11024 106372 11076
rect 106424 11064 106430 11076
rect 107378 11064 107384 11076
rect 106424 11036 107384 11064
rect 106424 11024 106430 11036
rect 107378 11024 107384 11036
rect 107436 11024 107442 11076
rect 108960 11064 108988 11095
rect 109126 11092 109132 11104
rect 109184 11092 109190 11144
rect 109034 11064 109040 11076
rect 108960 11036 109040 11064
rect 109034 11024 109040 11036
rect 109092 11024 109098 11076
rect 109236 11064 109264 11172
rect 109604 11144 109632 11240
rect 111150 11228 111156 11280
rect 111208 11268 111214 11280
rect 111429 11271 111487 11277
rect 111429 11268 111441 11271
rect 111208 11240 111441 11268
rect 111208 11228 111214 11240
rect 111429 11237 111441 11240
rect 111475 11237 111487 11271
rect 111429 11231 111487 11237
rect 111058 11160 111064 11212
rect 111116 11200 111122 11212
rect 111116 11172 111748 11200
rect 111116 11160 111122 11172
rect 109586 11132 109592 11144
rect 109499 11104 109592 11132
rect 109586 11092 109592 11104
rect 109644 11132 109650 11144
rect 110969 11135 111027 11141
rect 110969 11132 110981 11135
rect 109644 11104 110981 11132
rect 109644 11092 109650 11104
rect 110969 11101 110981 11104
rect 111015 11101 111027 11135
rect 111610 11132 111616 11144
rect 111571 11104 111616 11132
rect 110969 11095 111027 11101
rect 111610 11092 111616 11104
rect 111668 11092 111674 11144
rect 111720 11132 111748 11172
rect 113174 11160 113180 11212
rect 113232 11200 113238 11212
rect 113358 11200 113364 11212
rect 113232 11172 113364 11200
rect 113232 11160 113238 11172
rect 113358 11160 113364 11172
rect 113416 11160 113422 11212
rect 115201 11203 115259 11209
rect 115201 11169 115213 11203
rect 115247 11200 115259 11203
rect 115290 11200 115296 11212
rect 115247 11172 115296 11200
rect 115247 11169 115259 11172
rect 115201 11163 115259 11169
rect 115290 11160 115296 11172
rect 115348 11160 115354 11212
rect 115400 11132 115428 11308
rect 118418 11296 118424 11308
rect 118476 11296 118482 11348
rect 119430 11336 119436 11348
rect 118528 11308 119436 11336
rect 115474 11228 115480 11280
rect 115532 11268 115538 11280
rect 115934 11268 115940 11280
rect 115532 11240 115940 11268
rect 115532 11228 115538 11240
rect 115934 11228 115940 11240
rect 115992 11228 115998 11280
rect 116578 11228 116584 11280
rect 116636 11268 116642 11280
rect 117317 11271 117375 11277
rect 117317 11268 117329 11271
rect 116636 11240 117329 11268
rect 116636 11228 116642 11240
rect 117317 11237 117329 11240
rect 117363 11237 117375 11271
rect 117317 11231 117375 11237
rect 117498 11228 117504 11280
rect 117556 11268 117562 11280
rect 118528 11268 118556 11308
rect 119430 11296 119436 11308
rect 119488 11296 119494 11348
rect 119614 11336 119620 11348
rect 119575 11308 119620 11336
rect 119614 11296 119620 11308
rect 119672 11336 119678 11348
rect 120994 11336 121000 11348
rect 119672 11308 121000 11336
rect 119672 11296 119678 11308
rect 120994 11296 121000 11308
rect 121052 11336 121058 11348
rect 123021 11339 123079 11345
rect 123021 11336 123033 11339
rect 121052 11308 123033 11336
rect 121052 11296 121058 11308
rect 123021 11305 123033 11308
rect 123067 11305 123079 11339
rect 129090 11336 129096 11348
rect 123021 11299 123079 11305
rect 123128 11308 128354 11336
rect 129051 11308 129096 11336
rect 117556 11240 118556 11268
rect 117556 11228 117562 11240
rect 118602 11228 118608 11280
rect 118660 11268 118666 11280
rect 123128 11268 123156 11308
rect 118660 11240 123156 11268
rect 124033 11271 124091 11277
rect 118660 11228 118666 11240
rect 124033 11237 124045 11271
rect 124079 11237 124091 11271
rect 124033 11231 124091 11237
rect 115750 11200 115756 11212
rect 115711 11172 115756 11200
rect 115750 11160 115756 11172
rect 115808 11160 115814 11212
rect 115842 11160 115848 11212
rect 115900 11200 115906 11212
rect 118329 11203 118387 11209
rect 118329 11200 118341 11203
rect 115900 11172 118341 11200
rect 115900 11160 115906 11172
rect 118329 11169 118341 11172
rect 118375 11169 118387 11203
rect 118329 11163 118387 11169
rect 118418 11160 118424 11212
rect 118476 11200 118482 11212
rect 122469 11203 122527 11209
rect 122469 11200 122481 11203
rect 118476 11172 122481 11200
rect 118476 11160 118482 11172
rect 117406 11132 117412 11144
rect 111720 11104 115428 11132
rect 115492 11104 117412 11132
rect 110414 11064 110420 11076
rect 109236 11036 110420 11064
rect 110414 11024 110420 11036
rect 110472 11064 110478 11076
rect 110724 11067 110782 11073
rect 110724 11064 110736 11067
rect 110472 11036 110736 11064
rect 110472 11024 110478 11036
rect 110724 11033 110736 11036
rect 110770 11064 110782 11067
rect 111702 11064 111708 11076
rect 110770 11036 111708 11064
rect 110770 11033 110782 11036
rect 110724 11027 110782 11033
rect 111702 11024 111708 11036
rect 111760 11024 111766 11076
rect 112162 11064 112168 11076
rect 112123 11036 112168 11064
rect 112162 11024 112168 11036
rect 112220 11024 112226 11076
rect 112809 11067 112867 11073
rect 112809 11064 112821 11067
rect 112272 11036 112821 11064
rect 105556 10968 105860 10996
rect 105906 10956 105912 11008
rect 105964 10996 105970 11008
rect 111058 10996 111064 11008
rect 105964 10968 111064 10996
rect 105964 10956 105970 10968
rect 111058 10956 111064 10968
rect 111116 10956 111122 11008
rect 111242 10956 111248 11008
rect 111300 10996 111306 11008
rect 112272 10996 112300 11036
rect 112809 11033 112821 11036
rect 112855 11064 112867 11067
rect 114956 11067 115014 11073
rect 112855 11036 114876 11064
rect 112855 11033 112867 11036
rect 112809 11027 112867 11033
rect 111300 10968 112300 10996
rect 114848 10996 114876 11036
rect 114956 11033 114968 11067
rect 115002 11064 115014 11067
rect 115382 11064 115388 11076
rect 115002 11036 115388 11064
rect 115002 11033 115014 11036
rect 114956 11027 115014 11033
rect 115382 11024 115388 11036
rect 115440 11024 115446 11076
rect 115492 10996 115520 11104
rect 117406 11092 117412 11104
rect 117464 11092 117470 11144
rect 117498 11092 117504 11144
rect 117556 11132 117562 11144
rect 117556 11104 117601 11132
rect 117556 11092 117562 11104
rect 117774 11092 117780 11144
rect 117832 11132 117838 11144
rect 118605 11135 118663 11141
rect 118605 11132 118617 11135
rect 117832 11104 118617 11132
rect 117832 11092 117838 11104
rect 118605 11101 118617 11104
rect 118651 11101 118663 11135
rect 120166 11132 120172 11144
rect 120127 11104 120172 11132
rect 118605 11095 118663 11101
rect 120166 11092 120172 11104
rect 120224 11092 120230 11144
rect 120920 11141 120948 11172
rect 122469 11169 122481 11172
rect 122515 11169 122527 11203
rect 122469 11163 122527 11169
rect 123018 11160 123024 11212
rect 123076 11200 123082 11212
rect 124048 11200 124076 11231
rect 125686 11228 125692 11280
rect 125744 11268 125750 11280
rect 126793 11271 126851 11277
rect 126793 11268 126805 11271
rect 125744 11240 126805 11268
rect 125744 11228 125750 11240
rect 126793 11237 126805 11240
rect 126839 11237 126851 11271
rect 128326 11268 128354 11308
rect 129090 11296 129096 11308
rect 129148 11296 129154 11348
rect 129274 11296 129280 11348
rect 129332 11336 129338 11348
rect 132221 11339 132279 11345
rect 129332 11308 130516 11336
rect 129332 11296 129338 11308
rect 130488 11268 130516 11308
rect 132221 11305 132233 11339
rect 132267 11336 132279 11339
rect 132770 11336 132776 11348
rect 132267 11308 132776 11336
rect 132267 11305 132279 11308
rect 132221 11299 132279 11305
rect 132770 11296 132776 11308
rect 132828 11296 132834 11348
rect 133046 11296 133052 11348
rect 133104 11336 133110 11348
rect 134518 11336 134524 11348
rect 133104 11308 134380 11336
rect 134479 11308 134524 11336
rect 133104 11296 133110 11308
rect 134352 11268 134380 11308
rect 134518 11296 134524 11308
rect 134576 11296 134582 11348
rect 134702 11296 134708 11348
rect 134760 11336 134766 11348
rect 137002 11336 137008 11348
rect 134760 11308 137008 11336
rect 134760 11296 134766 11308
rect 137002 11296 137008 11308
rect 137060 11296 137066 11348
rect 138474 11296 138480 11348
rect 138532 11336 138538 11348
rect 139762 11336 139768 11348
rect 138532 11308 139768 11336
rect 138532 11296 138538 11308
rect 139762 11296 139768 11308
rect 139820 11296 139826 11348
rect 141068 11308 141280 11336
rect 128326 11240 129504 11268
rect 130488 11240 132632 11268
rect 134352 11240 138612 11268
rect 126793 11231 126851 11237
rect 123076 11172 124076 11200
rect 123076 11160 123082 11172
rect 120905 11135 120963 11141
rect 120905 11101 120917 11135
rect 120951 11101 120963 11135
rect 120905 11095 120963 11101
rect 120994 11092 121000 11144
rect 121052 11132 121058 11144
rect 121549 11135 121607 11141
rect 121052 11104 121097 11132
rect 121052 11092 121058 11104
rect 121549 11101 121561 11135
rect 121595 11132 121607 11135
rect 121914 11132 121920 11144
rect 121595 11104 121920 11132
rect 121595 11101 121607 11104
rect 121549 11095 121607 11101
rect 121914 11092 121920 11104
rect 121972 11132 121978 11144
rect 122558 11132 122564 11144
rect 121972 11104 122564 11132
rect 121972 11092 121978 11104
rect 122558 11092 122564 11104
rect 122616 11092 122622 11144
rect 122650 11092 122656 11144
rect 122708 11132 122714 11144
rect 124766 11132 124772 11144
rect 122708 11104 124772 11132
rect 122708 11092 122714 11104
rect 124766 11092 124772 11104
rect 124824 11092 124830 11144
rect 125146 11135 125204 11141
rect 125146 11101 125158 11135
rect 125192 11101 125204 11135
rect 125146 11095 125204 11101
rect 117222 11064 117228 11076
rect 116228 11036 117228 11064
rect 114848 10968 115520 10996
rect 111300 10956 111306 10968
rect 115934 10956 115940 11008
rect 115992 10996 115998 11008
rect 116228 11005 116256 11036
rect 117222 11024 117228 11036
rect 117280 11024 117286 11076
rect 117314 11024 117320 11076
rect 117372 11064 117378 11076
rect 119154 11064 119160 11076
rect 117372 11036 119160 11064
rect 117372 11024 117378 11036
rect 119154 11024 119160 11036
rect 119212 11024 119218 11076
rect 119614 11024 119620 11076
rect 119672 11064 119678 11076
rect 120721 11067 120779 11073
rect 120721 11064 120733 11067
rect 119672 11036 120733 11064
rect 119672 11024 119678 11036
rect 120721 11033 120733 11036
rect 120767 11033 120779 11067
rect 120721 11027 120779 11033
rect 121656 11036 121960 11064
rect 116213 10999 116271 11005
rect 116213 10996 116225 10999
rect 115992 10968 116225 10996
rect 115992 10956 115998 10968
rect 116213 10965 116225 10968
rect 116259 10965 116271 10999
rect 116213 10959 116271 10965
rect 116302 10956 116308 11008
rect 116360 10996 116366 11008
rect 121656 10996 121684 11036
rect 116360 10968 121684 10996
rect 121733 10999 121791 11005
rect 116360 10956 116366 10968
rect 121733 10965 121745 10999
rect 121779 10996 121791 10999
rect 121822 10996 121828 11008
rect 121779 10968 121828 10996
rect 121779 10965 121791 10968
rect 121733 10959 121791 10965
rect 121822 10956 121828 10968
rect 121880 10956 121886 11008
rect 121932 10996 121960 11036
rect 122098 11024 122104 11076
rect 122156 11064 122162 11076
rect 125152 11064 125180 11095
rect 125401 11092 125407 11144
rect 125459 11132 125465 11144
rect 125459 11104 125504 11132
rect 125459 11092 125465 11104
rect 125594 11092 125600 11144
rect 125652 11132 125658 11144
rect 126149 11135 126207 11141
rect 126149 11132 126161 11135
rect 125652 11104 126161 11132
rect 125652 11092 125658 11104
rect 126149 11101 126161 11104
rect 126195 11101 126207 11135
rect 126149 11095 126207 11101
rect 126238 11092 126244 11144
rect 126296 11132 126302 11144
rect 127802 11132 127808 11144
rect 126296 11104 126341 11132
rect 127763 11104 127808 11132
rect 126296 11092 126302 11104
rect 127802 11092 127808 11104
rect 127860 11092 127866 11144
rect 128078 11132 128084 11144
rect 128039 11104 128084 11132
rect 128078 11092 128084 11104
rect 128136 11092 128142 11144
rect 128262 11092 128268 11144
rect 128320 11132 128326 11144
rect 129366 11132 129372 11144
rect 128320 11104 129372 11132
rect 128320 11092 128326 11104
rect 129366 11092 129372 11104
rect 129424 11092 129430 11144
rect 129476 11132 129504 11240
rect 131853 11203 131911 11209
rect 131853 11169 131865 11203
rect 131899 11200 131911 11203
rect 132494 11200 132500 11212
rect 131899 11172 132500 11200
rect 131899 11169 131911 11172
rect 131853 11163 131911 11169
rect 132494 11160 132500 11172
rect 132552 11160 132558 11212
rect 130194 11132 130200 11144
rect 130252 11141 130258 11144
rect 129476 11104 130200 11132
rect 130194 11092 130200 11104
rect 130252 11095 130264 11141
rect 130473 11135 130531 11141
rect 130473 11101 130485 11135
rect 130519 11132 130531 11135
rect 130930 11132 130936 11144
rect 130519 11104 130936 11132
rect 130519 11101 130531 11104
rect 130473 11095 130531 11101
rect 130252 11092 130258 11095
rect 130930 11092 130936 11104
rect 130988 11092 130994 11144
rect 132037 11135 132095 11141
rect 132037 11101 132049 11135
rect 132083 11101 132095 11135
rect 132037 11095 132095 11101
rect 125226 11064 125232 11076
rect 122156 11036 123064 11064
rect 125152 11036 125232 11064
rect 122156 11024 122162 11036
rect 122926 10996 122932 11008
rect 121932 10968 122932 10996
rect 122926 10956 122932 10968
rect 122984 10956 122990 11008
rect 123036 10996 123064 11036
rect 125226 11024 125232 11036
rect 125284 11064 125290 11076
rect 125686 11064 125692 11076
rect 125284 11036 125692 11064
rect 125284 11024 125290 11036
rect 125686 11024 125692 11036
rect 125744 11024 125750 11076
rect 125778 11024 125784 11076
rect 125836 11064 125842 11076
rect 125965 11067 126023 11073
rect 125965 11064 125977 11067
rect 125836 11036 125977 11064
rect 125836 11024 125842 11036
rect 125965 11033 125977 11036
rect 126011 11033 126023 11067
rect 125965 11027 126023 11033
rect 126882 11024 126888 11076
rect 126940 11064 126946 11076
rect 130378 11064 130384 11076
rect 126940 11036 130384 11064
rect 126940 11024 126946 11036
rect 130378 11024 130384 11036
rect 130436 11024 130442 11076
rect 130746 11024 130752 11076
rect 130804 11064 130810 11076
rect 131301 11067 131359 11073
rect 131301 11064 131313 11067
rect 130804 11036 131313 11064
rect 130804 11024 130810 11036
rect 131301 11033 131313 11036
rect 131347 11064 131359 11067
rect 132052 11064 132080 11095
rect 131347 11036 132080 11064
rect 132604 11064 132632 11240
rect 133138 11200 133144 11212
rect 133099 11172 133144 11200
rect 133138 11160 133144 11172
rect 133196 11160 133202 11212
rect 137278 11160 137284 11212
rect 137336 11200 137342 11212
rect 137373 11203 137431 11209
rect 137373 11200 137385 11203
rect 137336 11172 137385 11200
rect 137336 11160 137342 11172
rect 137373 11169 137385 11172
rect 137419 11200 137431 11203
rect 138584 11200 138612 11240
rect 138658 11228 138664 11280
rect 138716 11268 138722 11280
rect 139489 11271 139547 11277
rect 139489 11268 139501 11271
rect 138716 11240 139501 11268
rect 138716 11228 138722 11240
rect 139489 11237 139501 11240
rect 139535 11237 139547 11271
rect 139489 11231 139547 11237
rect 141068 11200 141096 11308
rect 141252 11268 141280 11308
rect 141510 11296 141516 11348
rect 141568 11336 141574 11348
rect 147122 11336 147128 11348
rect 141568 11308 147128 11336
rect 141568 11296 141574 11308
rect 147122 11296 147128 11308
rect 147180 11296 147186 11348
rect 147306 11336 147312 11348
rect 147267 11308 147312 11336
rect 147306 11296 147312 11308
rect 147364 11296 147370 11348
rect 147490 11296 147496 11348
rect 147548 11336 147554 11348
rect 147766 11336 147772 11348
rect 147548 11308 147772 11336
rect 147548 11296 147554 11308
rect 147766 11296 147772 11308
rect 147824 11296 147830 11348
rect 149241 11339 149299 11345
rect 149241 11305 149253 11339
rect 149287 11336 149299 11339
rect 149330 11336 149336 11348
rect 149287 11308 149336 11336
rect 149287 11305 149299 11308
rect 149241 11299 149299 11305
rect 149330 11296 149336 11308
rect 149388 11296 149394 11348
rect 149974 11336 149980 11348
rect 149440 11308 149980 11336
rect 143810 11268 143816 11280
rect 141252 11240 143816 11268
rect 143810 11228 143816 11240
rect 143868 11228 143874 11280
rect 137419 11172 138520 11200
rect 138584 11172 141096 11200
rect 141160 11172 141464 11200
rect 137419 11169 137431 11172
rect 137373 11163 137431 11169
rect 133230 11092 133236 11144
rect 133288 11132 133294 11144
rect 138290 11132 138296 11144
rect 133288 11104 138296 11132
rect 133288 11092 133294 11104
rect 138290 11092 138296 11104
rect 138348 11092 138354 11144
rect 138492 11132 138520 11172
rect 139486 11132 139492 11144
rect 138492 11104 139492 11132
rect 139486 11092 139492 11104
rect 139544 11092 139550 11144
rect 140590 11132 140596 11144
rect 139596 11104 140596 11132
rect 133408 11067 133466 11073
rect 132604 11036 133368 11064
rect 131347 11033 131359 11036
rect 131301 11027 131359 11033
rect 123662 10996 123668 11008
rect 123036 10968 123668 10996
rect 123662 10956 123668 10968
rect 123720 10956 123726 11008
rect 125042 10956 125048 11008
rect 125100 10996 125106 11008
rect 129366 10996 129372 11008
rect 125100 10968 129372 10996
rect 125100 10956 125106 10968
rect 129366 10956 129372 10968
rect 129424 10996 129430 11008
rect 130562 10996 130568 11008
rect 129424 10968 130568 10996
rect 129424 10956 129430 10968
rect 130562 10956 130568 10968
rect 130620 10956 130626 11008
rect 133340 10996 133368 11036
rect 133408 11033 133420 11067
rect 133454 11064 133466 11067
rect 133690 11064 133696 11076
rect 133454 11036 133696 11064
rect 133454 11033 133466 11036
rect 133408 11027 133466 11033
rect 133690 11024 133696 11036
rect 133748 11024 133754 11076
rect 134702 11064 134708 11076
rect 133800 11036 134708 11064
rect 133800 10996 133828 11036
rect 134702 11024 134708 11036
rect 134760 11024 134766 11076
rect 135530 11064 135536 11076
rect 135491 11036 135536 11064
rect 135530 11024 135536 11036
rect 135588 11024 135594 11076
rect 135806 11024 135812 11076
rect 135864 11064 135870 11076
rect 136082 11064 136088 11076
rect 135864 11036 136088 11064
rect 135864 11024 135870 11036
rect 136082 11024 136088 11036
rect 136140 11024 136146 11076
rect 136821 11067 136879 11073
rect 136821 11033 136833 11067
rect 136867 11064 136879 11067
rect 139596 11064 139624 11104
rect 140590 11092 140596 11104
rect 140648 11132 140654 11144
rect 141160 11132 141188 11172
rect 140648 11104 141188 11132
rect 141237 11135 141295 11141
rect 140648 11092 140654 11104
rect 141237 11101 141249 11135
rect 141283 11134 141295 11135
rect 141326 11134 141332 11144
rect 141283 11106 141332 11134
rect 141283 11101 141295 11106
rect 141237 11095 141295 11101
rect 141326 11092 141332 11106
rect 141384 11092 141390 11144
rect 141436 11141 141464 11172
rect 141602 11160 141608 11212
rect 141660 11200 141666 11212
rect 144822 11200 144828 11212
rect 141660 11172 143856 11200
rect 144783 11172 144828 11200
rect 141660 11160 141666 11172
rect 141421 11135 141479 11141
rect 141421 11101 141433 11135
rect 141467 11101 141479 11135
rect 141421 11095 141479 11101
rect 142157 11135 142215 11141
rect 142157 11101 142169 11135
rect 142203 11101 142215 11135
rect 142157 11095 142215 11101
rect 142341 11135 142399 11141
rect 142341 11101 142353 11135
rect 142387 11132 142399 11135
rect 142982 11132 142988 11144
rect 142387 11104 142988 11132
rect 142387 11101 142399 11104
rect 142341 11095 142399 11101
rect 136867 11036 139624 11064
rect 139765 11067 139823 11073
rect 136867 11033 136879 11036
rect 136821 11027 136879 11033
rect 139765 11033 139777 11067
rect 139811 11064 139823 11067
rect 140409 11067 140467 11073
rect 140409 11064 140421 11067
rect 139811 11036 140421 11064
rect 139811 11033 139823 11036
rect 139765 11027 139823 11033
rect 140409 11033 140421 11036
rect 140455 11064 140467 11067
rect 140682 11064 140688 11076
rect 140455 11036 140688 11064
rect 140455 11033 140467 11036
rect 140409 11027 140467 11033
rect 140682 11024 140688 11036
rect 140740 11024 140746 11076
rect 141050 11064 141056 11076
rect 141011 11036 141056 11064
rect 141050 11024 141056 11036
rect 141108 11024 141114 11076
rect 141602 11024 141608 11076
rect 141660 11064 141666 11076
rect 141973 11067 142031 11073
rect 141973 11064 141985 11067
rect 141660 11036 141985 11064
rect 141660 11024 141666 11036
rect 141973 11033 141985 11036
rect 142019 11033 142031 11067
rect 142172 11064 142200 11095
rect 142982 11092 142988 11104
rect 143040 11092 143046 11144
rect 143828 11132 143856 11172
rect 144822 11160 144828 11172
rect 144880 11160 144886 11212
rect 144914 11160 144920 11212
rect 144972 11160 144978 11212
rect 147324 11200 147352 11296
rect 148597 11203 148655 11209
rect 148597 11200 148609 11203
rect 147324 11172 148609 11200
rect 148597 11169 148609 11172
rect 148643 11169 148655 11203
rect 148597 11163 148655 11169
rect 144932 11132 144960 11160
rect 143828 11104 144960 11132
rect 146570 11092 146576 11144
rect 146628 11132 146634 11144
rect 146665 11135 146723 11141
rect 146665 11132 146677 11135
rect 146628 11104 146677 11132
rect 146628 11092 146634 11104
rect 146665 11101 146677 11104
rect 146711 11101 146723 11135
rect 146665 11095 146723 11101
rect 146846 11092 146852 11144
rect 146904 11132 146910 11144
rect 147125 11135 147183 11141
rect 147125 11132 147137 11135
rect 146904 11104 147137 11132
rect 146904 11092 146910 11104
rect 147125 11101 147137 11104
rect 147171 11101 147183 11135
rect 147125 11095 147183 11101
rect 147646 11104 148364 11132
rect 143994 11064 144000 11076
rect 142172 11036 144000 11064
rect 141973 11027 142031 11033
rect 143994 11024 144000 11036
rect 144052 11024 144058 11076
rect 144546 11024 144552 11076
rect 144604 11073 144610 11076
rect 144604 11064 144616 11073
rect 146420 11067 146478 11073
rect 144604 11036 144649 11064
rect 144604 11027 144616 11036
rect 146420 11033 146432 11067
rect 146466 11064 146478 11067
rect 147646 11064 147674 11104
rect 148226 11064 148232 11076
rect 146466 11036 147674 11064
rect 148187 11036 148232 11064
rect 146466 11033 146478 11036
rect 146420 11027 146478 11033
rect 144604 11024 144610 11027
rect 148226 11024 148232 11036
rect 148284 11024 148290 11076
rect 148336 11064 148364 11104
rect 148410 11092 148416 11144
rect 148468 11132 148474 11144
rect 148468 11104 148513 11132
rect 148468 11092 148474 11104
rect 149440 11064 149468 11308
rect 149974 11296 149980 11308
rect 150032 11296 150038 11348
rect 150434 11296 150440 11348
rect 150492 11336 150498 11348
rect 150802 11336 150808 11348
rect 150492 11308 150808 11336
rect 150492 11296 150498 11308
rect 150802 11296 150808 11308
rect 150860 11296 150866 11348
rect 150986 11296 150992 11348
rect 151044 11336 151050 11348
rect 151081 11339 151139 11345
rect 151081 11336 151093 11339
rect 151044 11308 151093 11336
rect 151044 11296 151050 11308
rect 151081 11305 151093 11308
rect 151127 11305 151139 11339
rect 151081 11299 151139 11305
rect 153194 11296 153200 11348
rect 153252 11336 153258 11348
rect 153381 11339 153439 11345
rect 153381 11336 153393 11339
rect 153252 11308 153393 11336
rect 153252 11296 153258 11308
rect 153381 11305 153393 11308
rect 153427 11305 153439 11339
rect 153381 11299 153439 11305
rect 153470 11296 153476 11348
rect 153528 11336 153534 11348
rect 153528 11308 155448 11336
rect 153528 11296 153534 11308
rect 150621 11203 150679 11209
rect 150621 11169 150633 11203
rect 150667 11200 150679 11203
rect 151354 11200 151360 11212
rect 150667 11172 151360 11200
rect 150667 11169 150679 11172
rect 150621 11163 150679 11169
rect 149606 11092 149612 11144
rect 149664 11132 149670 11144
rect 150636 11132 150664 11163
rect 151354 11160 151360 11172
rect 151412 11160 151418 11212
rect 152458 11200 152464 11212
rect 152419 11172 152464 11200
rect 152458 11160 152464 11172
rect 152516 11160 152522 11212
rect 155218 11200 155224 11212
rect 154684 11172 155224 11200
rect 149664 11104 150664 11132
rect 149664 11092 149670 11104
rect 151262 11092 151268 11144
rect 151320 11132 151326 11144
rect 154494 11135 154552 11141
rect 154494 11132 154506 11135
rect 151320 11104 154506 11132
rect 151320 11092 151326 11104
rect 154494 11101 154506 11104
rect 154540 11132 154552 11135
rect 154684 11132 154712 11172
rect 155218 11160 155224 11172
rect 155276 11160 155282 11212
rect 155420 11141 155448 11308
rect 155678 11296 155684 11348
rect 155736 11336 155742 11348
rect 156046 11336 156052 11348
rect 155736 11308 156052 11336
rect 155736 11296 155742 11308
rect 156046 11296 156052 11308
rect 156104 11296 156110 11348
rect 156877 11339 156935 11345
rect 156877 11305 156889 11339
rect 156923 11336 156935 11339
rect 159450 11336 159456 11348
rect 156923 11308 159456 11336
rect 156923 11305 156935 11308
rect 156877 11299 156935 11305
rect 159450 11296 159456 11308
rect 159508 11296 159514 11348
rect 157521 11271 157579 11277
rect 157521 11237 157533 11271
rect 157567 11268 157579 11271
rect 158346 11268 158352 11280
rect 157567 11240 158352 11268
rect 157567 11237 157579 11240
rect 157521 11231 157579 11237
rect 158346 11228 158352 11240
rect 158404 11228 158410 11280
rect 155494 11160 155500 11212
rect 155552 11200 155558 11212
rect 155552 11172 157104 11200
rect 155552 11160 155558 11172
rect 154540 11104 154712 11132
rect 154761 11135 154819 11141
rect 154540 11101 154552 11104
rect 154494 11095 154552 11101
rect 154761 11101 154773 11135
rect 154807 11101 154819 11135
rect 154761 11095 154819 11101
rect 155405 11135 155463 11141
rect 155405 11101 155417 11135
rect 155451 11101 155463 11135
rect 155405 11095 155463 11101
rect 155589 11135 155647 11141
rect 155589 11101 155601 11135
rect 155635 11132 155647 11135
rect 155954 11132 155960 11144
rect 155635 11104 155960 11132
rect 155635 11101 155647 11104
rect 155589 11095 155647 11101
rect 148336 11036 149468 11064
rect 149514 11024 149520 11076
rect 149572 11064 149578 11076
rect 150354 11067 150412 11073
rect 150354 11064 150366 11067
rect 149572 11036 150366 11064
rect 149572 11024 149578 11036
rect 150354 11033 150366 11036
rect 150400 11033 150412 11067
rect 150354 11027 150412 11033
rect 152194 11067 152252 11073
rect 152194 11033 152206 11067
rect 152240 11064 152252 11067
rect 152240 11036 153976 11064
rect 152240 11033 152252 11036
rect 152194 11027 152252 11033
rect 133340 10968 133828 10996
rect 134426 10956 134432 11008
rect 134484 10996 134490 11008
rect 134978 10996 134984 11008
rect 134484 10968 134984 10996
rect 134484 10956 134490 10968
rect 134978 10956 134984 10968
rect 135036 10956 135042 11008
rect 135070 10956 135076 11008
rect 135128 10996 135134 11008
rect 141326 10996 141332 11008
rect 135128 10968 141332 10996
rect 135128 10956 135134 10968
rect 141326 10956 141332 10968
rect 141384 10956 141390 11008
rect 143166 10956 143172 11008
rect 143224 10996 143230 11008
rect 143442 10996 143448 11008
rect 143224 10968 143448 10996
rect 143224 10956 143230 10968
rect 143442 10956 143448 10968
rect 143500 10956 143506 11008
rect 145282 10996 145288 11008
rect 145243 10968 145288 10996
rect 145282 10956 145288 10968
rect 145340 10956 145346 11008
rect 145374 10956 145380 11008
rect 145432 10996 145438 11008
rect 149330 10996 149336 11008
rect 145432 10968 149336 10996
rect 145432 10956 145438 10968
rect 149330 10956 149336 10968
rect 149388 10956 149394 11008
rect 151538 10956 151544 11008
rect 151596 10996 151602 11008
rect 152200 10996 152228 11027
rect 151596 10968 152228 10996
rect 153948 10996 153976 11036
rect 154022 11024 154028 11076
rect 154080 11064 154086 11076
rect 154390 11064 154396 11076
rect 154080 11036 154396 11064
rect 154080 11024 154086 11036
rect 154390 11024 154396 11036
rect 154448 11064 154454 11076
rect 154776 11064 154804 11095
rect 155954 11092 155960 11104
rect 156012 11132 156018 11144
rect 156049 11135 156107 11141
rect 156049 11132 156061 11135
rect 156012 11104 156061 11132
rect 156012 11092 156018 11104
rect 156049 11101 156061 11104
rect 156095 11101 156107 11135
rect 156230 11132 156236 11144
rect 156191 11104 156236 11132
rect 156049 11095 156107 11101
rect 156230 11092 156236 11104
rect 156288 11092 156294 11144
rect 157076 11141 157104 11172
rect 157061 11135 157119 11141
rect 157061 11101 157073 11135
rect 157107 11101 157119 11135
rect 157061 11095 157119 11101
rect 157705 11135 157763 11141
rect 157705 11101 157717 11135
rect 157751 11132 157763 11135
rect 158622 11132 158628 11144
rect 157751 11104 158628 11132
rect 157751 11101 157763 11104
rect 157705 11095 157763 11101
rect 158622 11092 158628 11104
rect 158680 11092 158686 11144
rect 154448 11036 154804 11064
rect 154448 11024 154454 11036
rect 154850 11024 154856 11076
rect 154908 11064 154914 11076
rect 155221 11067 155279 11073
rect 155221 11064 155233 11067
rect 154908 11036 155233 11064
rect 154908 11024 154914 11036
rect 155221 11033 155233 11036
rect 155267 11033 155279 11067
rect 156138 11064 156144 11076
rect 155221 11027 155279 11033
rect 155328 11036 156144 11064
rect 155328 10996 155356 11036
rect 156138 11024 156144 11036
rect 156196 11024 156202 11076
rect 156414 11064 156420 11076
rect 156375 11036 156420 11064
rect 156414 11024 156420 11036
rect 156472 11024 156478 11076
rect 153948 10968 155356 10996
rect 151596 10956 151602 10968
rect 155402 10956 155408 11008
rect 155460 10996 155466 11008
rect 157426 10996 157432 11008
rect 155460 10968 157432 10996
rect 155460 10956 155466 10968
rect 157426 10956 157432 10968
rect 157484 10956 157490 11008
rect 1104 10906 159043 10928
rect 1104 10854 40394 10906
rect 40446 10854 40458 10906
rect 40510 10854 40522 10906
rect 40574 10854 40586 10906
rect 40638 10854 40650 10906
rect 40702 10854 79839 10906
rect 79891 10854 79903 10906
rect 79955 10854 79967 10906
rect 80019 10854 80031 10906
rect 80083 10854 80095 10906
rect 80147 10854 119284 10906
rect 119336 10854 119348 10906
rect 119400 10854 119412 10906
rect 119464 10854 119476 10906
rect 119528 10854 119540 10906
rect 119592 10854 158729 10906
rect 158781 10854 158793 10906
rect 158845 10854 158857 10906
rect 158909 10854 158921 10906
rect 158973 10854 158985 10906
rect 159037 10854 159043 10906
rect 1104 10832 159043 10854
rect 5718 10792 5724 10804
rect 5679 10764 5724 10792
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 12308 10764 13829 10792
rect 12308 10752 12314 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 13817 10755 13875 10761
rect 4056 10727 4114 10733
rect 4056 10693 4068 10727
rect 4102 10724 4114 10727
rect 4154 10724 4160 10736
rect 4102 10696 4160 10724
rect 4102 10693 4114 10696
rect 4056 10687 4114 10693
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8386 10656 8392 10668
rect 8343 10628 8392 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 11072 10656 11100 10752
rect 12066 10733 12072 10736
rect 12060 10724 12072 10733
rect 12027 10696 12072 10724
rect 12060 10687 12072 10696
rect 12066 10684 12072 10687
rect 12124 10684 12130 10736
rect 13832 10724 13860 10755
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 18598 10792 18604 10804
rect 15396 10764 18604 10792
rect 15396 10724 15424 10764
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 18785 10795 18843 10801
rect 18785 10761 18797 10795
rect 18831 10761 18843 10795
rect 18785 10755 18843 10761
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19426 10792 19432 10804
rect 19383 10764 19432 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 13832 10696 15424 10724
rect 16942 10684 16948 10736
rect 17000 10724 17006 10736
rect 17650 10727 17708 10733
rect 17650 10724 17662 10727
rect 17000 10696 17662 10724
rect 17000 10684 17006 10696
rect 17650 10693 17662 10696
rect 17696 10693 17708 10727
rect 17650 10687 17708 10693
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11072 10628 11805 10656
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 13630 10656 13636 10668
rect 13591 10628 13636 10656
rect 11793 10619 11851 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 15378 10656 15384 10668
rect 14691 10628 15384 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 16574 10656 16580 10668
rect 15519 10628 16580 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17034 10656 17040 10668
rect 16899 10628 17040 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 17034 10616 17040 10628
rect 17092 10656 17098 10668
rect 17405 10660 17463 10665
rect 17328 10659 17463 10660
rect 17328 10656 17417 10659
rect 17092 10632 17417 10656
rect 17092 10628 17356 10632
rect 17092 10616 17098 10628
rect 17405 10625 17417 10632
rect 17451 10625 17463 10659
rect 18800 10656 18828 10755
rect 19426 10752 19432 10764
rect 19484 10792 19490 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19484 10764 19809 10792
rect 19484 10752 19490 10764
rect 19797 10761 19809 10764
rect 19843 10792 19855 10795
rect 20530 10792 20536 10804
rect 19843 10764 20536 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22097 10795 22155 10801
rect 22097 10792 22109 10795
rect 22060 10764 22109 10792
rect 22060 10752 22066 10764
rect 22097 10761 22109 10764
rect 22143 10792 22155 10795
rect 24857 10795 24915 10801
rect 24857 10792 24869 10795
rect 22143 10764 24869 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 24857 10761 24869 10764
rect 24903 10792 24915 10795
rect 25130 10792 25136 10804
rect 24903 10764 25136 10792
rect 24903 10761 24915 10764
rect 24857 10755 24915 10761
rect 25130 10752 25136 10764
rect 25188 10752 25194 10804
rect 26602 10792 26608 10804
rect 26563 10764 26608 10792
rect 26602 10752 26608 10764
rect 26660 10752 26666 10804
rect 27614 10792 27620 10804
rect 27172 10764 27620 10792
rect 25501 10727 25559 10733
rect 25501 10693 25513 10727
rect 25547 10724 25559 10727
rect 27172 10724 27200 10764
rect 27614 10752 27620 10764
rect 27672 10752 27678 10804
rect 27706 10752 27712 10804
rect 27764 10792 27770 10804
rect 27801 10795 27859 10801
rect 27801 10792 27813 10795
rect 27764 10764 27813 10792
rect 27764 10752 27770 10764
rect 27801 10761 27813 10764
rect 27847 10761 27859 10795
rect 27801 10755 27859 10761
rect 29086 10752 29092 10804
rect 29144 10792 29150 10804
rect 30098 10792 30104 10804
rect 29144 10764 30104 10792
rect 29144 10752 29150 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 30190 10752 30196 10804
rect 30248 10792 30254 10804
rect 33226 10792 33232 10804
rect 30248 10764 33232 10792
rect 30248 10752 30254 10764
rect 33226 10752 33232 10764
rect 33284 10752 33290 10804
rect 33318 10752 33324 10804
rect 33376 10792 33382 10804
rect 36909 10795 36967 10801
rect 36909 10792 36921 10795
rect 33376 10764 36921 10792
rect 33376 10752 33382 10764
rect 36909 10761 36921 10764
rect 36955 10761 36967 10795
rect 36909 10755 36967 10761
rect 37553 10795 37611 10801
rect 37553 10761 37565 10795
rect 37599 10792 37611 10795
rect 37642 10792 37648 10804
rect 37599 10764 37648 10792
rect 37599 10761 37611 10764
rect 37553 10755 37611 10761
rect 37642 10752 37648 10764
rect 37700 10752 37706 10804
rect 40034 10792 40040 10804
rect 39995 10764 40040 10792
rect 40034 10752 40040 10764
rect 40092 10752 40098 10804
rect 40402 10752 40408 10804
rect 40460 10792 40466 10804
rect 41506 10792 41512 10804
rect 40460 10764 41512 10792
rect 40460 10752 40466 10764
rect 41506 10752 41512 10764
rect 41564 10752 41570 10804
rect 42610 10752 42616 10804
rect 42668 10792 42674 10804
rect 44818 10792 44824 10804
rect 42668 10764 44824 10792
rect 42668 10752 42674 10764
rect 44818 10752 44824 10764
rect 44876 10752 44882 10804
rect 44910 10752 44916 10804
rect 44968 10792 44974 10804
rect 45097 10795 45155 10801
rect 45097 10792 45109 10795
rect 44968 10764 45109 10792
rect 44968 10752 44974 10764
rect 45097 10761 45109 10764
rect 45143 10761 45155 10795
rect 45097 10755 45155 10761
rect 45833 10795 45891 10801
rect 45833 10761 45845 10795
rect 45879 10792 45891 10795
rect 46106 10792 46112 10804
rect 45879 10764 46112 10792
rect 45879 10761 45891 10764
rect 45833 10755 45891 10761
rect 46106 10752 46112 10764
rect 46164 10752 46170 10804
rect 48498 10752 48504 10804
rect 48556 10792 48562 10804
rect 49418 10792 49424 10804
rect 48556 10764 49424 10792
rect 48556 10752 48562 10764
rect 49418 10752 49424 10764
rect 49476 10752 49482 10804
rect 49789 10795 49847 10801
rect 49789 10761 49801 10795
rect 49835 10761 49847 10795
rect 49789 10755 49847 10761
rect 51077 10795 51135 10801
rect 51077 10761 51089 10795
rect 51123 10792 51135 10795
rect 52638 10792 52644 10804
rect 51123 10764 52644 10792
rect 51123 10761 51135 10764
rect 51077 10755 51135 10761
rect 25547 10696 27200 10724
rect 25547 10693 25559 10696
rect 25501 10687 25559 10693
rect 27246 10684 27252 10736
rect 27304 10724 27310 10736
rect 33502 10724 33508 10736
rect 27304 10696 29224 10724
rect 27304 10684 27310 10696
rect 28350 10656 28356 10668
rect 17405 10619 17463 10625
rect 17512 10628 18460 10656
rect 18800 10628 28356 10656
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 17512 10588 17540 10628
rect 9171 10560 10088 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 10060 10464 10088 10560
rect 13188 10560 17540 10588
rect 18432 10588 18460 10628
rect 28350 10616 28356 10628
rect 28408 10616 28414 10668
rect 29196 10665 29224 10696
rect 29932 10696 33508 10724
rect 28925 10659 28983 10665
rect 28925 10625 28937 10659
rect 28971 10656 28983 10659
rect 29181 10659 29239 10665
rect 28971 10628 29132 10656
rect 28971 10625 28983 10628
rect 28925 10619 28983 10625
rect 22186 10588 22192 10600
rect 18432 10560 22192 10588
rect 13188 10529 13216 10560
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 23014 10588 23020 10600
rect 22927 10560 23020 10588
rect 23014 10548 23020 10560
rect 23072 10588 23078 10600
rect 27338 10588 27344 10600
rect 23072 10560 27344 10588
rect 23072 10548 23078 10560
rect 27338 10548 27344 10560
rect 27396 10548 27402 10600
rect 29104 10588 29132 10628
rect 29181 10625 29193 10659
rect 29227 10656 29239 10659
rect 29546 10656 29552 10668
rect 29227 10628 29552 10656
rect 29227 10625 29239 10628
rect 29181 10619 29239 10625
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 29932 10588 29960 10696
rect 33502 10684 33508 10696
rect 33560 10684 33566 10736
rect 38841 10727 38899 10733
rect 38841 10724 38853 10727
rect 34348 10696 38853 10724
rect 30098 10616 30104 10668
rect 30156 10656 30162 10668
rect 30265 10659 30323 10665
rect 30265 10656 30277 10659
rect 30156 10628 30277 10656
rect 30156 10616 30162 10628
rect 30265 10625 30277 10628
rect 30311 10625 30323 10659
rect 32953 10659 33011 10665
rect 32953 10656 32965 10659
rect 30265 10619 30323 10625
rect 31036 10628 31754 10656
rect 29104 10560 29960 10588
rect 30006 10548 30012 10600
rect 30064 10588 30070 10600
rect 30064 10560 30109 10588
rect 30064 10548 30070 10560
rect 13173 10523 13231 10529
rect 13173 10489 13185 10523
rect 13219 10489 13231 10523
rect 13173 10483 13231 10489
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 15654 10520 15660 10532
rect 14875 10492 15660 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 15764 10492 16988 10520
rect 5166 10452 5172 10464
rect 5127 10424 5172 10452
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 8113 10455 8171 10461
rect 8113 10421 8125 10455
rect 8159 10452 8171 10455
rect 8202 10452 8208 10464
rect 8159 10424 8208 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 9490 10452 9496 10464
rect 9451 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 15764 10452 15792 10492
rect 13688 10424 15792 10452
rect 16117 10455 16175 10461
rect 13688 10412 13694 10424
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16666 10452 16672 10464
rect 16163 10424 16672 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16960 10452 16988 10492
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 18564 10492 27384 10520
rect 18564 10480 18570 10492
rect 19978 10452 19984 10464
rect 16960 10424 19984 10452
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 21358 10452 21364 10464
rect 21319 10424 21364 10452
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 23750 10452 23756 10464
rect 23711 10424 23756 10452
rect 23750 10412 23756 10424
rect 23808 10412 23814 10464
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 25961 10455 26019 10461
rect 25961 10452 25973 10455
rect 25648 10424 25973 10452
rect 25648 10412 25654 10424
rect 25961 10421 25973 10424
rect 26007 10452 26019 10455
rect 26970 10452 26976 10464
rect 26007 10424 26976 10452
rect 26007 10421 26019 10424
rect 25961 10415 26019 10421
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 27246 10452 27252 10464
rect 27207 10424 27252 10452
rect 27246 10412 27252 10424
rect 27304 10412 27310 10464
rect 27356 10452 27384 10492
rect 31036 10452 31064 10628
rect 31202 10548 31208 10600
rect 31260 10588 31266 10600
rect 31260 10560 31432 10588
rect 31260 10548 31266 10560
rect 31404 10529 31432 10560
rect 31389 10523 31447 10529
rect 31389 10489 31401 10523
rect 31435 10489 31447 10523
rect 31726 10520 31754 10628
rect 32416 10628 32965 10656
rect 32416 10529 32444 10628
rect 32953 10625 32965 10628
rect 32999 10625 33011 10659
rect 33870 10656 33876 10668
rect 33831 10628 33876 10656
rect 32953 10619 33011 10625
rect 33870 10616 33876 10628
rect 33928 10616 33934 10668
rect 33594 10548 33600 10600
rect 33652 10588 33658 10600
rect 33689 10591 33747 10597
rect 33689 10588 33701 10591
rect 33652 10560 33701 10588
rect 33652 10548 33658 10560
rect 33689 10557 33701 10560
rect 33735 10557 33747 10591
rect 33689 10551 33747 10557
rect 32401 10523 32459 10529
rect 32401 10520 32413 10523
rect 31726 10492 32413 10520
rect 31389 10483 31447 10489
rect 32401 10489 32413 10492
rect 32447 10489 32459 10523
rect 34348 10520 34376 10696
rect 38841 10693 38853 10696
rect 38887 10693 38899 10727
rect 40052 10724 40080 10752
rect 45922 10724 45928 10736
rect 40052 10696 44036 10724
rect 38841 10687 38899 10693
rect 35785 10659 35843 10665
rect 35785 10656 35797 10659
rect 34992 10628 35797 10656
rect 34422 10548 34428 10600
rect 34480 10588 34486 10600
rect 34992 10597 35020 10628
rect 35785 10625 35797 10628
rect 35831 10625 35843 10659
rect 38856 10656 38884 10687
rect 40218 10656 40224 10668
rect 38856 10628 40224 10656
rect 35785 10619 35843 10625
rect 40218 10616 40224 10628
rect 40276 10616 40282 10668
rect 40497 10659 40555 10665
rect 40497 10625 40509 10659
rect 40543 10656 40555 10659
rect 41138 10656 41144 10668
rect 40543 10628 41144 10656
rect 40543 10625 40555 10628
rect 40497 10619 40555 10625
rect 41138 10616 41144 10628
rect 41196 10616 41202 10668
rect 41322 10656 41328 10668
rect 41283 10628 41328 10656
rect 41322 10616 41328 10628
rect 41380 10616 41386 10668
rect 44008 10665 44036 10696
rect 44468 10696 45928 10724
rect 44468 10665 44496 10696
rect 45922 10684 45928 10696
rect 45980 10684 45986 10736
rect 46014 10684 46020 10736
rect 46072 10724 46078 10736
rect 48590 10724 48596 10736
rect 46072 10696 48596 10724
rect 46072 10684 46078 10696
rect 48590 10684 48596 10696
rect 48648 10684 48654 10736
rect 49804 10724 49832 10755
rect 52638 10752 52644 10764
rect 52696 10752 52702 10804
rect 55674 10792 55680 10804
rect 55635 10764 55680 10792
rect 55674 10752 55680 10764
rect 55732 10752 55738 10804
rect 56318 10752 56324 10804
rect 56376 10752 56382 10804
rect 57517 10795 57575 10801
rect 57517 10761 57529 10795
rect 57563 10792 57575 10795
rect 57698 10792 57704 10804
rect 57563 10764 57704 10792
rect 57563 10761 57575 10764
rect 57517 10755 57575 10761
rect 57698 10752 57704 10764
rect 57756 10752 57762 10804
rect 58250 10752 58256 10804
rect 58308 10792 58314 10804
rect 59170 10792 59176 10804
rect 58308 10764 59176 10792
rect 58308 10752 58314 10764
rect 59170 10752 59176 10764
rect 59228 10752 59234 10804
rect 60645 10795 60703 10801
rect 60645 10761 60657 10795
rect 60691 10792 60703 10795
rect 81066 10792 81072 10804
rect 60691 10764 80054 10792
rect 81027 10764 81072 10792
rect 60691 10761 60703 10764
rect 60645 10755 60703 10761
rect 53558 10724 53564 10736
rect 49804 10696 53564 10724
rect 53558 10684 53564 10696
rect 53616 10684 53622 10736
rect 55214 10724 55220 10736
rect 54312 10696 55220 10724
rect 41877 10659 41935 10665
rect 41877 10625 41889 10659
rect 41923 10625 41935 10659
rect 41877 10619 41935 10625
rect 43737 10659 43795 10665
rect 43737 10625 43749 10659
rect 43783 10656 43795 10659
rect 43993 10659 44051 10665
rect 43783 10628 43944 10656
rect 43783 10625 43795 10628
rect 43737 10619 43795 10625
rect 34977 10591 35035 10597
rect 34977 10588 34989 10591
rect 34480 10560 34989 10588
rect 34480 10548 34486 10560
rect 34977 10557 34989 10560
rect 35023 10557 35035 10591
rect 34977 10551 35035 10557
rect 35250 10548 35256 10600
rect 35308 10588 35314 10600
rect 35529 10591 35587 10597
rect 35529 10588 35541 10591
rect 35308 10560 35541 10588
rect 35308 10548 35314 10560
rect 35529 10557 35541 10560
rect 35575 10557 35587 10591
rect 40236 10588 40264 10616
rect 41782 10588 41788 10600
rect 40236 10560 41788 10588
rect 35529 10551 35587 10557
rect 41782 10548 41788 10560
rect 41840 10588 41846 10600
rect 41892 10588 41920 10619
rect 41840 10560 41920 10588
rect 43916 10588 43944 10628
rect 43993 10625 44005 10659
rect 44039 10656 44051 10659
rect 44453 10659 44511 10665
rect 44453 10656 44465 10659
rect 44039 10628 44465 10656
rect 44039 10625 44051 10628
rect 43993 10619 44051 10625
rect 44453 10625 44465 10628
rect 44499 10625 44511 10659
rect 44453 10619 44511 10625
rect 45281 10659 45339 10665
rect 45281 10625 45293 10659
rect 45327 10625 45339 10659
rect 45281 10619 45339 10625
rect 44910 10588 44916 10600
rect 43916 10560 44916 10588
rect 41840 10548 41846 10560
rect 44910 10548 44916 10560
rect 44968 10548 44974 10600
rect 32401 10483 32459 10489
rect 33060 10492 34376 10520
rect 27356 10424 31064 10452
rect 31294 10412 31300 10464
rect 31352 10452 31358 10464
rect 33060 10452 33088 10492
rect 40034 10480 40040 10532
rect 40092 10520 40098 10532
rect 41141 10523 41199 10529
rect 41141 10520 41153 10523
rect 40092 10492 41153 10520
rect 40092 10480 40098 10492
rect 41141 10489 41153 10492
rect 41187 10489 41199 10523
rect 41141 10483 41199 10489
rect 41230 10480 41236 10532
rect 41288 10520 41294 10532
rect 41288 10492 43116 10520
rect 41288 10480 41294 10492
rect 31352 10424 33088 10452
rect 33137 10455 33195 10461
rect 31352 10412 31358 10424
rect 33137 10421 33149 10455
rect 33183 10452 33195 10455
rect 33778 10452 33784 10464
rect 33183 10424 33784 10452
rect 33183 10421 33195 10424
rect 33137 10415 33195 10421
rect 33778 10412 33784 10424
rect 33836 10412 33842 10464
rect 34057 10455 34115 10461
rect 34057 10421 34069 10455
rect 34103 10452 34115 10455
rect 36446 10452 36452 10464
rect 34103 10424 36452 10452
rect 34103 10421 34115 10424
rect 34057 10415 34115 10421
rect 36446 10412 36452 10424
rect 36504 10412 36510 10464
rect 39390 10452 39396 10464
rect 39351 10424 39396 10452
rect 39390 10412 39396 10424
rect 39448 10452 39454 10464
rect 40126 10452 40132 10464
rect 39448 10424 40132 10452
rect 39448 10412 39454 10424
rect 40126 10412 40132 10424
rect 40184 10412 40190 10464
rect 40681 10455 40739 10461
rect 40681 10421 40693 10455
rect 40727 10452 40739 10455
rect 40954 10452 40960 10464
rect 40727 10424 40960 10452
rect 40727 10421 40739 10424
rect 40681 10415 40739 10421
rect 40954 10412 40960 10424
rect 41012 10412 41018 10464
rect 41690 10412 41696 10464
rect 41748 10452 41754 10464
rect 41969 10455 42027 10461
rect 41969 10452 41981 10455
rect 41748 10424 41981 10452
rect 41748 10412 41754 10424
rect 41969 10421 41981 10424
rect 42015 10421 42027 10455
rect 42610 10452 42616 10464
rect 42571 10424 42616 10452
rect 41969 10415 42027 10421
rect 42610 10412 42616 10424
rect 42668 10412 42674 10464
rect 43088 10452 43116 10492
rect 45186 10452 45192 10464
rect 43088 10424 45192 10452
rect 45186 10412 45192 10424
rect 45244 10412 45250 10464
rect 45296 10452 45324 10619
rect 45370 10616 45376 10668
rect 45428 10656 45434 10668
rect 46946 10659 47004 10665
rect 46946 10656 46958 10659
rect 45428 10628 46958 10656
rect 45428 10616 45434 10628
rect 46946 10625 46958 10628
rect 46992 10625 47004 10659
rect 47210 10656 47216 10668
rect 47171 10628 47216 10656
rect 46946 10619 47004 10625
rect 47210 10616 47216 10628
rect 47268 10616 47274 10668
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 48406 10656 48412 10668
rect 48367 10628 48412 10656
rect 48406 10616 48412 10628
rect 48464 10616 48470 10668
rect 48676 10659 48734 10665
rect 48676 10625 48688 10659
rect 48722 10656 48734 10659
rect 49878 10656 49884 10668
rect 48722 10628 49884 10656
rect 48722 10625 48734 10628
rect 48676 10619 48734 10625
rect 49878 10616 49884 10628
rect 49936 10616 49942 10668
rect 50430 10656 50436 10668
rect 50391 10628 50436 10656
rect 50430 10616 50436 10628
rect 50488 10616 50494 10668
rect 50890 10656 50896 10668
rect 50851 10628 50896 10656
rect 50890 10616 50896 10628
rect 50948 10616 50954 10668
rect 51813 10659 51871 10665
rect 51813 10656 51825 10659
rect 51046 10628 51825 10656
rect 49418 10548 49424 10600
rect 49476 10588 49482 10600
rect 51046 10588 51074 10628
rect 51813 10625 51825 10628
rect 51859 10625 51871 10659
rect 51813 10619 51871 10625
rect 51902 10616 51908 10668
rect 51960 10656 51966 10668
rect 51960 10628 52005 10656
rect 51960 10616 51966 10628
rect 52638 10616 52644 10668
rect 52696 10656 52702 10668
rect 54312 10665 54340 10696
rect 55214 10684 55220 10696
rect 55272 10684 55278 10736
rect 54297 10659 54355 10665
rect 54297 10656 54309 10659
rect 52696 10628 54309 10656
rect 52696 10616 52702 10628
rect 54297 10625 54309 10628
rect 54343 10625 54355 10659
rect 54297 10619 54355 10625
rect 54564 10659 54622 10665
rect 54564 10625 54576 10659
rect 54610 10656 54622 10659
rect 56042 10656 56048 10668
rect 54610 10628 56048 10656
rect 54610 10625 54622 10628
rect 54564 10619 54622 10625
rect 56042 10616 56048 10628
rect 56100 10616 56106 10668
rect 56336 10656 56364 10752
rect 56502 10684 56508 10736
rect 56560 10724 56566 10736
rect 58066 10724 58072 10736
rect 56560 10696 58072 10724
rect 56560 10684 56566 10696
rect 58066 10684 58072 10696
rect 58124 10684 58130 10736
rect 59280 10696 60412 10724
rect 56393 10659 56451 10665
rect 56393 10656 56405 10659
rect 56336 10628 56405 10656
rect 56393 10625 56405 10628
rect 56439 10656 56451 10659
rect 58342 10656 58348 10668
rect 56439 10628 58348 10656
rect 56439 10625 56451 10628
rect 56393 10619 56451 10625
rect 58342 10616 58348 10628
rect 58400 10616 58406 10668
rect 58805 10659 58863 10665
rect 58621 10649 58679 10655
rect 58621 10615 58633 10649
rect 58667 10615 58679 10649
rect 58805 10625 58817 10659
rect 58851 10656 58863 10659
rect 58851 10628 59032 10656
rect 58851 10625 58863 10628
rect 58805 10619 58863 10625
rect 58621 10609 58679 10615
rect 49476 10560 51074 10588
rect 49476 10548 49482 10560
rect 51166 10548 51172 10600
rect 51224 10588 51230 10600
rect 52917 10591 52975 10597
rect 51224 10560 52224 10588
rect 51224 10548 51230 10560
rect 49510 10480 49516 10532
rect 49568 10520 49574 10532
rect 50249 10523 50307 10529
rect 50249 10520 50261 10523
rect 49568 10492 50261 10520
rect 49568 10480 49574 10492
rect 50249 10489 50261 10492
rect 50295 10489 50307 10523
rect 50249 10483 50307 10489
rect 50430 10480 50436 10532
rect 50488 10520 50494 10532
rect 51629 10523 51687 10529
rect 51629 10520 51641 10523
rect 50488 10492 51641 10520
rect 50488 10480 50494 10492
rect 51629 10489 51641 10492
rect 51675 10489 51687 10523
rect 52196 10520 52224 10560
rect 52917 10557 52929 10591
rect 52963 10557 52975 10591
rect 52917 10551 52975 10557
rect 52932 10520 52960 10551
rect 53006 10548 53012 10600
rect 53064 10588 53070 10600
rect 53193 10591 53251 10597
rect 53193 10588 53205 10591
rect 53064 10560 53205 10588
rect 53064 10548 53070 10560
rect 53193 10557 53205 10560
rect 53239 10557 53251 10591
rect 53193 10551 53251 10557
rect 52196 10492 52960 10520
rect 51629 10483 51687 10489
rect 47854 10452 47860 10464
rect 45296 10424 47860 10452
rect 47854 10412 47860 10424
rect 47912 10412 47918 10464
rect 47949 10455 48007 10461
rect 47949 10421 47961 10455
rect 47995 10452 48007 10455
rect 48038 10452 48044 10464
rect 47995 10424 48044 10452
rect 47995 10421 48007 10424
rect 47949 10415 48007 10421
rect 48038 10412 48044 10424
rect 48096 10412 48102 10464
rect 53208 10452 53236 10551
rect 55306 10548 55312 10600
rect 55364 10588 55370 10600
rect 55766 10588 55772 10600
rect 55364 10560 55772 10588
rect 55364 10548 55370 10560
rect 55766 10548 55772 10560
rect 55824 10588 55830 10600
rect 56137 10591 56195 10597
rect 56137 10588 56149 10591
rect 55824 10560 56149 10588
rect 55824 10548 55830 10560
rect 56137 10557 56149 10560
rect 56183 10557 56195 10591
rect 56137 10551 56195 10557
rect 58636 10532 58664 10609
rect 59004 10588 59032 10628
rect 59078 10616 59084 10668
rect 59136 10656 59142 10668
rect 59280 10665 59308 10696
rect 59265 10659 59323 10665
rect 59265 10656 59277 10659
rect 59136 10628 59277 10656
rect 59136 10616 59142 10628
rect 59265 10625 59277 10628
rect 59311 10625 59323 10659
rect 59265 10619 59323 10625
rect 59532 10659 59590 10665
rect 59532 10625 59544 10659
rect 59578 10656 59590 10659
rect 59998 10656 60004 10668
rect 59578 10628 60004 10656
rect 59578 10625 59590 10628
rect 59532 10619 59590 10625
rect 59998 10616 60004 10628
rect 60056 10616 60062 10668
rect 60384 10656 60412 10696
rect 60734 10684 60740 10736
rect 60792 10724 60798 10736
rect 61350 10727 61408 10733
rect 61350 10724 61362 10727
rect 60792 10696 61362 10724
rect 60792 10684 60798 10696
rect 61350 10693 61362 10696
rect 61396 10693 61408 10727
rect 61350 10687 61408 10693
rect 64230 10684 64236 10736
rect 64288 10724 64294 10736
rect 68557 10727 68615 10733
rect 68557 10724 68569 10727
rect 64288 10696 68569 10724
rect 64288 10684 64294 10696
rect 68557 10693 68569 10696
rect 68603 10724 68615 10727
rect 69290 10724 69296 10736
rect 68603 10696 69296 10724
rect 68603 10693 68615 10696
rect 68557 10687 68615 10693
rect 69290 10684 69296 10696
rect 69348 10684 69354 10736
rect 72697 10727 72755 10733
rect 69400 10696 72556 10724
rect 60642 10656 60648 10668
rect 60384 10628 60648 10656
rect 60642 10616 60648 10628
rect 60700 10656 60706 10668
rect 61105 10659 61163 10665
rect 61105 10656 61117 10659
rect 60700 10628 61117 10656
rect 60700 10616 60706 10628
rect 61105 10625 61117 10628
rect 61151 10625 61163 10659
rect 63862 10656 63868 10668
rect 63775 10628 63868 10656
rect 61105 10619 61163 10625
rect 63862 10616 63868 10628
rect 63920 10616 63926 10668
rect 64138 10616 64144 10668
rect 64196 10656 64202 10668
rect 64509 10659 64567 10665
rect 64509 10656 64521 10659
rect 64196 10628 64521 10656
rect 64196 10616 64202 10628
rect 64509 10625 64521 10628
rect 64555 10625 64567 10659
rect 64509 10619 64567 10625
rect 66921 10659 66979 10665
rect 66921 10625 66933 10659
rect 66967 10656 66979 10659
rect 68922 10656 68928 10668
rect 66967 10628 68928 10656
rect 66967 10625 66979 10628
rect 66921 10619 66979 10625
rect 68922 10616 68928 10628
rect 68980 10656 68986 10668
rect 69400 10656 69428 10696
rect 68980 10628 69428 10656
rect 69928 10659 69986 10665
rect 68980 10616 68986 10628
rect 69928 10625 69940 10659
rect 69974 10656 69986 10659
rect 70486 10656 70492 10668
rect 69974 10628 70492 10656
rect 69974 10625 69986 10628
rect 69928 10619 69986 10625
rect 70486 10616 70492 10628
rect 70544 10616 70550 10668
rect 72528 10665 72556 10696
rect 72697 10693 72709 10727
rect 72743 10724 72755 10727
rect 74442 10724 74448 10736
rect 72743 10696 74448 10724
rect 72743 10693 72755 10696
rect 72697 10687 72755 10693
rect 74442 10684 74448 10696
rect 74500 10684 74506 10736
rect 78950 10724 78956 10736
rect 74552 10696 78956 10724
rect 72513 10659 72571 10665
rect 72513 10625 72525 10659
rect 72559 10625 72571 10659
rect 72513 10619 72571 10625
rect 72602 10616 72608 10668
rect 72660 10656 72666 10668
rect 73709 10659 73767 10665
rect 73709 10656 73721 10659
rect 72660 10628 73721 10656
rect 72660 10616 72666 10628
rect 73709 10625 73721 10628
rect 73755 10625 73767 10659
rect 73709 10619 73767 10625
rect 73893 10659 73951 10665
rect 73893 10625 73905 10659
rect 73939 10656 73951 10659
rect 74552 10656 74580 10696
rect 78950 10684 78956 10696
rect 79008 10684 79014 10736
rect 79134 10724 79140 10736
rect 79095 10696 79140 10724
rect 79134 10684 79140 10696
rect 79192 10724 79198 10736
rect 79870 10724 79876 10736
rect 79192 10696 79876 10724
rect 79192 10684 79198 10696
rect 79870 10684 79876 10696
rect 79928 10733 79934 10736
rect 79928 10727 79992 10733
rect 79928 10693 79946 10727
rect 79980 10693 79992 10727
rect 80026 10724 80054 10764
rect 81066 10752 81072 10764
rect 81124 10752 81130 10804
rect 84930 10792 84936 10804
rect 81176 10764 84936 10792
rect 81176 10724 81204 10764
rect 84930 10752 84936 10764
rect 84988 10752 84994 10804
rect 86678 10752 86684 10804
rect 86736 10792 86742 10804
rect 87693 10795 87751 10801
rect 87693 10792 87705 10795
rect 86736 10764 87705 10792
rect 86736 10752 86742 10764
rect 83826 10724 83832 10736
rect 80026 10696 81204 10724
rect 82096 10696 83832 10724
rect 79928 10687 79992 10693
rect 79928 10684 79934 10687
rect 73939 10628 74580 10656
rect 73939 10625 73951 10628
rect 73893 10619 73951 10625
rect 74626 10616 74632 10668
rect 74684 10656 74690 10668
rect 75926 10659 75984 10665
rect 75926 10656 75938 10659
rect 74684 10628 75938 10656
rect 74684 10616 74690 10628
rect 75926 10625 75938 10628
rect 75972 10625 75984 10659
rect 76190 10656 76196 10668
rect 76151 10628 76196 10656
rect 75926 10619 75984 10625
rect 76190 10616 76196 10628
rect 76248 10656 76254 10668
rect 76466 10656 76472 10668
rect 76248 10628 76472 10656
rect 76248 10616 76254 10628
rect 76466 10616 76472 10628
rect 76524 10616 76530 10668
rect 76742 10656 76748 10668
rect 76703 10628 76748 10656
rect 76742 10616 76748 10628
rect 76800 10616 76806 10668
rect 77012 10659 77070 10665
rect 77012 10625 77024 10659
rect 77058 10656 77070 10659
rect 77846 10656 77852 10668
rect 77058 10628 77852 10656
rect 77058 10625 77070 10628
rect 77012 10619 77070 10625
rect 77846 10616 77852 10628
rect 77904 10616 77910 10668
rect 82096 10665 82124 10696
rect 83826 10684 83832 10696
rect 83884 10684 83890 10736
rect 86436 10727 86494 10733
rect 86436 10693 86448 10727
rect 86482 10724 86494 10727
rect 87230 10724 87236 10736
rect 86482 10696 87236 10724
rect 86482 10693 86494 10696
rect 86436 10687 86494 10693
rect 87230 10684 87236 10696
rect 87288 10684 87294 10736
rect 82081 10659 82139 10665
rect 82081 10625 82093 10659
rect 82127 10625 82139 10659
rect 82081 10619 82139 10625
rect 82725 10659 82783 10665
rect 82725 10625 82737 10659
rect 82771 10654 82783 10659
rect 86681 10659 86739 10665
rect 82771 10626 82860 10654
rect 82771 10625 82783 10626
rect 82725 10619 82783 10625
rect 59170 10588 59176 10600
rect 59004 10560 59176 10588
rect 59170 10548 59176 10560
rect 59228 10548 59234 10600
rect 62206 10548 62212 10600
rect 62264 10588 62270 10600
rect 63402 10588 63408 10600
rect 62264 10560 63408 10588
rect 62264 10548 62270 10560
rect 63402 10548 63408 10560
rect 63460 10588 63466 10600
rect 63681 10591 63739 10597
rect 63681 10588 63693 10591
rect 63460 10560 63693 10588
rect 63460 10548 63466 10560
rect 63681 10557 63693 10560
rect 63727 10557 63739 10591
rect 63880 10588 63908 10616
rect 67174 10588 67180 10600
rect 63880 10560 65288 10588
rect 67135 10560 67180 10588
rect 63681 10551 63739 10557
rect 57422 10480 57428 10532
rect 57480 10520 57486 10532
rect 57480 10492 58572 10520
rect 57480 10480 57486 10492
rect 55306 10452 55312 10464
rect 53208 10424 55312 10452
rect 55306 10412 55312 10424
rect 55364 10412 55370 10464
rect 58066 10412 58072 10464
rect 58124 10452 58130 10464
rect 58437 10455 58495 10461
rect 58437 10452 58449 10455
rect 58124 10424 58449 10452
rect 58124 10412 58130 10424
rect 58437 10421 58449 10424
rect 58483 10421 58495 10455
rect 58544 10452 58572 10492
rect 58618 10480 58624 10532
rect 58676 10480 58682 10532
rect 62482 10520 62488 10532
rect 62443 10492 62488 10520
rect 62482 10480 62488 10492
rect 62540 10480 62546 10532
rect 62022 10452 62028 10464
rect 58544 10424 62028 10452
rect 58437 10415 58495 10421
rect 62022 10412 62028 10424
rect 62080 10412 62086 10464
rect 64049 10455 64107 10461
rect 64049 10421 64061 10455
rect 64095 10452 64107 10455
rect 64598 10452 64604 10464
rect 64095 10424 64604 10452
rect 64095 10421 64107 10424
rect 64049 10415 64107 10421
rect 64598 10412 64604 10424
rect 64656 10412 64662 10464
rect 64690 10412 64696 10464
rect 64748 10452 64754 10464
rect 65260 10461 65288 10560
rect 67174 10548 67180 10560
rect 67232 10548 67238 10600
rect 69661 10591 69719 10597
rect 69661 10588 69673 10591
rect 69124 10560 69673 10588
rect 65794 10520 65800 10532
rect 65755 10492 65800 10520
rect 65794 10480 65800 10492
rect 65852 10480 65858 10532
rect 65245 10455 65303 10461
rect 64748 10424 64793 10452
rect 64748 10412 64754 10424
rect 65245 10421 65257 10455
rect 65291 10452 65303 10455
rect 66254 10452 66260 10464
rect 65291 10424 66260 10452
rect 65291 10421 65303 10424
rect 65245 10415 65303 10421
rect 66254 10412 66260 10424
rect 66312 10412 66318 10464
rect 67818 10452 67824 10464
rect 67779 10424 67824 10452
rect 67818 10412 67824 10424
rect 67876 10412 67882 10464
rect 68370 10412 68376 10464
rect 68428 10452 68434 10464
rect 68738 10452 68744 10464
rect 68428 10424 68744 10452
rect 68428 10412 68434 10424
rect 68738 10412 68744 10424
rect 68796 10452 68802 10464
rect 69124 10461 69152 10560
rect 69661 10557 69673 10560
rect 69707 10557 69719 10591
rect 69661 10551 69719 10557
rect 71774 10548 71780 10600
rect 71832 10588 71838 10600
rect 72329 10591 72387 10597
rect 72329 10588 72341 10591
rect 71832 10560 72341 10588
rect 71832 10548 71838 10560
rect 72329 10557 72341 10560
rect 72375 10557 72387 10591
rect 72329 10551 72387 10557
rect 73525 10591 73583 10597
rect 73525 10557 73537 10591
rect 73571 10588 73583 10591
rect 74350 10588 74356 10600
rect 73571 10560 74356 10588
rect 73571 10557 73583 10560
rect 73525 10551 73583 10557
rect 74350 10548 74356 10560
rect 74408 10588 74414 10600
rect 74408 10560 75224 10588
rect 74408 10548 74414 10560
rect 71041 10523 71099 10529
rect 71041 10489 71053 10523
rect 71087 10520 71099 10523
rect 74718 10520 74724 10532
rect 71087 10492 74724 10520
rect 71087 10489 71099 10492
rect 71041 10483 71099 10489
rect 74718 10480 74724 10492
rect 74776 10480 74782 10532
rect 69109 10455 69167 10461
rect 69109 10452 69121 10455
rect 68796 10424 69121 10452
rect 68796 10412 68802 10424
rect 69109 10421 69121 10424
rect 69155 10421 69167 10455
rect 71774 10452 71780 10464
rect 71735 10424 71780 10452
rect 69109 10415 69167 10421
rect 71774 10412 71780 10424
rect 71832 10412 71838 10464
rect 74810 10452 74816 10464
rect 74771 10424 74816 10452
rect 74810 10412 74816 10424
rect 74868 10412 74874 10464
rect 75196 10452 75224 10560
rect 78858 10548 78864 10600
rect 78916 10588 78922 10600
rect 79686 10588 79692 10600
rect 78916 10560 79692 10588
rect 78916 10548 78922 10560
rect 79686 10548 79692 10560
rect 79744 10548 79750 10600
rect 82538 10588 82544 10600
rect 82499 10560 82544 10588
rect 82538 10548 82544 10560
rect 82596 10548 82602 10600
rect 82832 10588 82860 10626
rect 86681 10625 86693 10659
rect 86727 10656 86739 10659
rect 87340 10656 87368 10764
rect 87693 10761 87705 10764
rect 87739 10792 87751 10795
rect 89717 10795 89775 10801
rect 89717 10792 89729 10795
rect 87739 10764 89729 10792
rect 87739 10761 87751 10764
rect 87693 10755 87751 10761
rect 89717 10761 89729 10764
rect 89763 10792 89775 10795
rect 93210 10792 93216 10804
rect 89763 10764 93216 10792
rect 89763 10761 89775 10764
rect 89717 10755 89775 10761
rect 93210 10752 93216 10764
rect 93268 10752 93274 10804
rect 94406 10752 94412 10804
rect 94464 10792 94470 10804
rect 94464 10764 100708 10792
rect 94464 10752 94470 10764
rect 88334 10684 88340 10736
rect 88392 10724 88398 10736
rect 98822 10724 98828 10736
rect 88392 10696 98828 10724
rect 88392 10684 88398 10696
rect 98822 10684 98828 10696
rect 98880 10684 98886 10736
rect 98932 10696 100616 10724
rect 86727 10628 87368 10656
rect 86727 10625 86739 10628
rect 86681 10619 86739 10625
rect 87690 10616 87696 10668
rect 87748 10656 87754 10668
rect 87748 10628 88380 10656
rect 87748 10616 87754 10628
rect 82998 10588 83004 10600
rect 82832 10560 83004 10588
rect 82998 10548 83004 10560
rect 83056 10548 83062 10600
rect 83366 10548 83372 10600
rect 83424 10588 83430 10600
rect 84838 10588 84844 10600
rect 83424 10560 84844 10588
rect 83424 10548 83430 10560
rect 84838 10548 84844 10560
rect 84896 10548 84902 10600
rect 86862 10548 86868 10600
rect 86920 10588 86926 10600
rect 88352 10588 88380 10628
rect 88426 10616 88432 10668
rect 88484 10656 88490 10668
rect 89073 10659 89131 10665
rect 89073 10656 89085 10659
rect 88484 10628 89085 10656
rect 88484 10616 88490 10628
rect 89073 10625 89085 10628
rect 89119 10656 89131 10659
rect 89162 10656 89168 10668
rect 89119 10628 89168 10656
rect 89119 10625 89131 10628
rect 89073 10619 89131 10625
rect 89162 10616 89168 10628
rect 89220 10616 89226 10668
rect 89257 10659 89315 10665
rect 89257 10625 89269 10659
rect 89303 10656 89315 10659
rect 90450 10656 90456 10668
rect 89303 10628 90456 10656
rect 89303 10625 89315 10628
rect 89257 10619 89315 10625
rect 90450 10616 90456 10628
rect 90508 10616 90514 10668
rect 91761 10659 91819 10665
rect 91761 10625 91773 10659
rect 91807 10656 91819 10659
rect 94314 10656 94320 10668
rect 91807 10628 94320 10656
rect 91807 10625 91819 10628
rect 91761 10619 91819 10625
rect 94314 10616 94320 10628
rect 94372 10616 94378 10668
rect 94774 10616 94780 10668
rect 94832 10656 94838 10668
rect 98932 10656 98960 10696
rect 94832 10628 98960 10656
rect 94832 10616 94838 10628
rect 88886 10588 88892 10600
rect 86920 10560 87552 10588
rect 88352 10560 88892 10588
rect 86920 10548 86926 10560
rect 78125 10523 78183 10529
rect 78125 10489 78137 10523
rect 78171 10520 78183 10523
rect 87230 10520 87236 10532
rect 78171 10492 79640 10520
rect 78171 10489 78183 10492
rect 78125 10483 78183 10489
rect 76374 10452 76380 10464
rect 75196 10424 76380 10452
rect 76374 10412 76380 10424
rect 76432 10412 76438 10464
rect 79612 10452 79640 10492
rect 81728 10492 85436 10520
rect 87191 10492 87236 10520
rect 81728 10452 81756 10492
rect 81894 10452 81900 10464
rect 79612 10424 81756 10452
rect 81855 10424 81900 10452
rect 81894 10412 81900 10424
rect 81952 10412 81958 10464
rect 82909 10455 82967 10461
rect 82909 10421 82921 10455
rect 82955 10452 82967 10455
rect 83826 10452 83832 10464
rect 82955 10424 83832 10452
rect 82955 10421 82967 10424
rect 82909 10415 82967 10421
rect 83826 10412 83832 10424
rect 83884 10412 83890 10464
rect 84562 10412 84568 10464
rect 84620 10452 84626 10464
rect 85298 10452 85304 10464
rect 84620 10424 85304 10452
rect 84620 10412 84626 10424
rect 85298 10412 85304 10424
rect 85356 10412 85362 10464
rect 85408 10452 85436 10492
rect 87230 10480 87236 10492
rect 87288 10480 87294 10532
rect 87524 10520 87552 10560
rect 88886 10548 88892 10560
rect 88944 10548 88950 10600
rect 92014 10588 92020 10600
rect 91975 10560 92020 10588
rect 92014 10548 92020 10560
rect 92072 10588 92078 10600
rect 92290 10588 92296 10600
rect 92072 10560 92296 10588
rect 92072 10548 92078 10560
rect 92290 10548 92296 10560
rect 92348 10548 92354 10600
rect 93026 10548 93032 10600
rect 93084 10588 93090 10600
rect 98822 10588 98828 10600
rect 93084 10560 98828 10588
rect 93084 10548 93090 10560
rect 98822 10548 98828 10560
rect 98880 10548 98886 10600
rect 100588 10588 100616 10696
rect 100680 10656 100708 10764
rect 100846 10752 100852 10804
rect 100904 10792 100910 10804
rect 102134 10792 102140 10804
rect 100904 10764 102140 10792
rect 100904 10752 100910 10764
rect 102134 10752 102140 10764
rect 102192 10752 102198 10804
rect 102226 10752 102232 10804
rect 102284 10792 102290 10804
rect 103517 10795 103575 10801
rect 102284 10764 102456 10792
rect 102284 10752 102290 10764
rect 101984 10727 102042 10733
rect 101984 10693 101996 10727
rect 102030 10724 102042 10727
rect 102318 10724 102324 10736
rect 102030 10696 102324 10724
rect 102030 10693 102042 10696
rect 101984 10687 102042 10693
rect 102318 10684 102324 10696
rect 102376 10684 102382 10736
rect 102229 10659 102287 10665
rect 100680 10628 102180 10656
rect 102152 10588 102180 10628
rect 102229 10625 102241 10659
rect 102275 10656 102287 10659
rect 102428 10656 102456 10764
rect 103517 10761 103529 10795
rect 103563 10792 103575 10795
rect 103790 10792 103796 10804
rect 103563 10764 103796 10792
rect 103563 10761 103575 10764
rect 103517 10755 103575 10761
rect 103790 10752 103796 10764
rect 103848 10752 103854 10804
rect 106461 10795 106519 10801
rect 106461 10761 106473 10795
rect 106507 10792 106519 10795
rect 107746 10792 107752 10804
rect 106507 10764 107752 10792
rect 106507 10761 106519 10764
rect 106461 10755 106519 10761
rect 107746 10752 107752 10764
rect 107804 10752 107810 10804
rect 108669 10795 108727 10801
rect 108669 10761 108681 10795
rect 108715 10792 108727 10795
rect 108942 10792 108948 10804
rect 108715 10764 108948 10792
rect 108715 10761 108727 10764
rect 108669 10755 108727 10761
rect 102781 10727 102839 10733
rect 102781 10693 102793 10727
rect 102827 10724 102839 10727
rect 103422 10724 103428 10736
rect 102827 10696 103428 10724
rect 102827 10693 102839 10696
rect 102781 10687 102839 10693
rect 102796 10656 102824 10687
rect 103422 10684 103428 10696
rect 103480 10724 103486 10736
rect 104342 10724 104348 10736
rect 103480 10696 104348 10724
rect 103480 10684 103486 10696
rect 104342 10684 104348 10696
rect 104400 10724 104406 10736
rect 104529 10727 104587 10733
rect 104529 10724 104541 10727
rect 104400 10696 104541 10724
rect 104400 10684 104406 10696
rect 104529 10693 104541 10696
rect 104575 10724 104587 10727
rect 107562 10724 107568 10736
rect 104575 10696 107568 10724
rect 104575 10693 104587 10696
rect 104529 10687 104587 10693
rect 103330 10656 103336 10668
rect 102275 10628 102824 10656
rect 103243 10628 103336 10656
rect 102275 10625 102287 10628
rect 102229 10619 102287 10625
rect 103330 10616 103336 10628
rect 103388 10656 103394 10668
rect 105096 10665 105124 10696
rect 107562 10684 107568 10696
rect 107620 10684 107626 10736
rect 108684 10724 108712 10755
rect 108942 10752 108948 10764
rect 109000 10752 109006 10804
rect 109034 10752 109040 10804
rect 109092 10792 109098 10804
rect 110598 10792 110604 10804
rect 109092 10764 110604 10792
rect 109092 10752 109098 10764
rect 110598 10752 110604 10764
rect 110656 10752 110662 10804
rect 110874 10752 110880 10804
rect 110932 10792 110938 10804
rect 111518 10792 111524 10804
rect 110932 10764 111524 10792
rect 110932 10752 110938 10764
rect 111518 10752 111524 10764
rect 111576 10792 111582 10804
rect 112625 10795 112683 10801
rect 112625 10792 112637 10795
rect 111576 10764 112637 10792
rect 111576 10752 111582 10764
rect 112625 10761 112637 10764
rect 112671 10792 112683 10795
rect 112714 10792 112720 10804
rect 112671 10764 112720 10792
rect 112671 10761 112683 10764
rect 112625 10755 112683 10761
rect 112714 10752 112720 10764
rect 112772 10752 112778 10804
rect 112898 10752 112904 10804
rect 112956 10792 112962 10804
rect 113637 10795 113695 10801
rect 113637 10792 113649 10795
rect 112956 10764 113649 10792
rect 112956 10752 112962 10764
rect 113637 10761 113649 10764
rect 113683 10761 113695 10795
rect 113637 10755 113695 10761
rect 114833 10795 114891 10801
rect 114833 10761 114845 10795
rect 114879 10792 114891 10795
rect 115290 10792 115296 10804
rect 114879 10764 115296 10792
rect 114879 10761 114891 10764
rect 114833 10755 114891 10761
rect 115290 10752 115296 10764
rect 115348 10752 115354 10804
rect 115658 10752 115664 10804
rect 115716 10792 115722 10804
rect 115937 10795 115995 10801
rect 115937 10792 115949 10795
rect 115716 10764 115949 10792
rect 115716 10752 115722 10764
rect 115937 10761 115949 10764
rect 115983 10761 115995 10795
rect 115937 10755 115995 10761
rect 116210 10752 116216 10804
rect 116268 10792 116274 10804
rect 116268 10764 117104 10792
rect 116268 10752 116274 10764
rect 116946 10724 116952 10736
rect 107764 10696 108712 10724
rect 108776 10696 116952 10724
rect 105081 10659 105139 10665
rect 103388 10628 104572 10656
rect 103388 10616 103394 10628
rect 104544 10600 104572 10628
rect 105081 10625 105093 10659
rect 105127 10625 105139 10659
rect 105081 10619 105139 10625
rect 105348 10659 105406 10665
rect 105348 10625 105360 10659
rect 105394 10656 105406 10659
rect 107013 10659 107071 10665
rect 107013 10656 107025 10659
rect 105394 10628 107025 10656
rect 105394 10625 105406 10628
rect 105348 10619 105406 10625
rect 107013 10625 107025 10628
rect 107059 10656 107071 10659
rect 107470 10656 107476 10668
rect 107059 10628 107476 10656
rect 107059 10625 107071 10628
rect 107013 10619 107071 10625
rect 107470 10616 107476 10628
rect 107528 10616 107534 10668
rect 107764 10665 107792 10696
rect 107749 10659 107807 10665
rect 107749 10625 107761 10659
rect 107795 10625 107807 10659
rect 107749 10619 107807 10625
rect 107933 10659 107991 10665
rect 107933 10625 107945 10659
rect 107979 10625 107991 10659
rect 107933 10619 107991 10625
rect 104066 10588 104072 10600
rect 100588 10560 101260 10588
rect 102152 10560 104072 10588
rect 90637 10523 90695 10529
rect 90637 10520 90649 10523
rect 87524 10492 90649 10520
rect 90637 10489 90649 10492
rect 90683 10489 90695 10523
rect 101122 10520 101128 10532
rect 90637 10483 90695 10489
rect 92032 10492 101128 10520
rect 88334 10452 88340 10464
rect 85408 10424 88340 10452
rect 88334 10412 88340 10424
rect 88392 10412 88398 10464
rect 88429 10455 88487 10461
rect 88429 10421 88441 10455
rect 88475 10452 88487 10455
rect 88518 10452 88524 10464
rect 88475 10424 88524 10452
rect 88475 10421 88487 10424
rect 88429 10415 88487 10421
rect 88518 10412 88524 10424
rect 88576 10412 88582 10464
rect 90266 10412 90272 10464
rect 90324 10452 90330 10464
rect 92032 10452 92060 10492
rect 101122 10480 101128 10492
rect 101180 10480 101186 10532
rect 92750 10452 92756 10464
rect 90324 10424 92060 10452
rect 92711 10424 92756 10452
rect 90324 10412 90330 10424
rect 92750 10412 92756 10424
rect 92808 10412 92814 10464
rect 93946 10412 93952 10464
rect 94004 10452 94010 10464
rect 94317 10455 94375 10461
rect 94317 10452 94329 10455
rect 94004 10424 94329 10452
rect 94004 10412 94010 10424
rect 94317 10421 94329 10424
rect 94363 10421 94375 10455
rect 94866 10452 94872 10464
rect 94827 10424 94872 10452
rect 94317 10415 94375 10421
rect 94866 10412 94872 10424
rect 94924 10412 94930 10464
rect 95326 10412 95332 10464
rect 95384 10452 95390 10464
rect 95421 10455 95479 10461
rect 95421 10452 95433 10455
rect 95384 10424 95433 10452
rect 95384 10412 95390 10424
rect 95421 10421 95433 10424
rect 95467 10421 95479 10455
rect 95421 10415 95479 10421
rect 95510 10412 95516 10464
rect 95568 10452 95574 10464
rect 95973 10455 96031 10461
rect 95973 10452 95985 10455
rect 95568 10424 95985 10452
rect 95568 10412 95574 10424
rect 95973 10421 95985 10424
rect 96019 10421 96031 10455
rect 95973 10415 96031 10421
rect 96709 10455 96767 10461
rect 96709 10421 96721 10455
rect 96755 10452 96767 10455
rect 97074 10452 97080 10464
rect 96755 10424 97080 10452
rect 96755 10421 96767 10424
rect 96709 10415 96767 10421
rect 97074 10412 97080 10424
rect 97132 10412 97138 10464
rect 98270 10452 98276 10464
rect 98231 10424 98276 10452
rect 98270 10412 98276 10424
rect 98328 10412 98334 10464
rect 98362 10412 98368 10464
rect 98420 10452 98426 10464
rect 100846 10452 100852 10464
rect 98420 10424 100852 10452
rect 98420 10412 98426 10424
rect 100846 10412 100852 10424
rect 100904 10412 100910 10464
rect 101232 10452 101260 10560
rect 104066 10548 104072 10560
rect 104124 10548 104130 10600
rect 104526 10548 104532 10600
rect 104584 10548 104590 10600
rect 107838 10548 107844 10600
rect 107896 10588 107902 10600
rect 107948 10588 107976 10619
rect 108206 10616 108212 10668
rect 108264 10656 108270 10668
rect 108776 10656 108804 10696
rect 116946 10684 116952 10696
rect 117004 10684 117010 10736
rect 117076 10733 117104 10764
rect 117682 10752 117688 10804
rect 117740 10792 117746 10804
rect 117777 10795 117835 10801
rect 117777 10792 117789 10795
rect 117740 10764 117789 10792
rect 117740 10752 117746 10764
rect 117777 10761 117789 10764
rect 117823 10761 117835 10795
rect 122650 10792 122656 10804
rect 117777 10755 117835 10761
rect 118160 10764 122656 10792
rect 117072 10727 117130 10733
rect 117072 10693 117084 10727
rect 117118 10693 117130 10727
rect 117072 10687 117130 10693
rect 108264 10628 108804 10656
rect 108264 10616 108270 10628
rect 110598 10616 110604 10668
rect 110656 10656 110662 10668
rect 110874 10656 110880 10668
rect 110656 10628 110880 10656
rect 110656 10616 110662 10628
rect 110874 10616 110880 10628
rect 110932 10616 110938 10668
rect 110966 10616 110972 10668
rect 111024 10656 111030 10668
rect 111426 10656 111432 10668
rect 111024 10628 111432 10656
rect 111024 10616 111030 10628
rect 111426 10616 111432 10628
rect 111484 10616 111490 10668
rect 111518 10616 111524 10668
rect 111576 10656 111582 10668
rect 111576 10628 111621 10656
rect 111576 10616 111582 10628
rect 111794 10616 111800 10668
rect 111852 10656 111858 10668
rect 113726 10656 113732 10668
rect 111852 10628 113732 10656
rect 111852 10616 111858 10628
rect 113726 10616 113732 10628
rect 113784 10616 113790 10668
rect 113821 10659 113879 10665
rect 113821 10625 113833 10659
rect 113867 10656 113879 10659
rect 114554 10656 114560 10668
rect 113867 10628 114560 10656
rect 113867 10625 113879 10628
rect 113821 10619 113879 10625
rect 114554 10616 114560 10628
rect 114612 10616 114618 10668
rect 117866 10656 117872 10668
rect 114664 10628 117872 10656
rect 107896 10560 107976 10588
rect 107896 10548 107902 10560
rect 109126 10548 109132 10600
rect 109184 10588 109190 10600
rect 109681 10591 109739 10597
rect 109681 10588 109693 10591
rect 109184 10560 109693 10588
rect 109184 10548 109190 10560
rect 109681 10557 109693 10560
rect 109727 10588 109739 10591
rect 110414 10588 110420 10600
rect 109727 10560 110420 10588
rect 109727 10557 109739 10560
rect 109681 10551 109739 10557
rect 110414 10548 110420 10560
rect 110472 10548 110478 10600
rect 110690 10548 110696 10600
rect 110748 10588 110754 10600
rect 114664 10588 114692 10628
rect 117866 10616 117872 10628
rect 117924 10616 117930 10668
rect 110748 10560 114692 10588
rect 110748 10548 110754 10560
rect 115658 10548 115664 10600
rect 115716 10588 115722 10600
rect 116210 10588 116216 10600
rect 115716 10560 116216 10588
rect 115716 10548 115722 10560
rect 116210 10548 116216 10560
rect 116268 10548 116274 10600
rect 117314 10588 117320 10600
rect 117275 10560 117320 10588
rect 117314 10548 117320 10560
rect 117372 10548 117378 10600
rect 107470 10480 107476 10532
rect 107528 10520 107534 10532
rect 107528 10492 108896 10520
rect 107528 10480 107534 10492
rect 107838 10452 107844 10464
rect 101232 10424 107844 10452
rect 107838 10412 107844 10424
rect 107896 10412 107902 10464
rect 108117 10455 108175 10461
rect 108117 10421 108129 10455
rect 108163 10452 108175 10455
rect 108482 10452 108488 10464
rect 108163 10424 108488 10452
rect 108163 10421 108175 10424
rect 108117 10415 108175 10421
rect 108482 10412 108488 10424
rect 108540 10412 108546 10464
rect 108868 10452 108896 10492
rect 111610 10480 111616 10532
rect 111668 10520 111674 10532
rect 118160 10520 118188 10764
rect 122650 10752 122656 10764
rect 122708 10752 122714 10804
rect 122926 10752 122932 10804
rect 122984 10792 122990 10804
rect 125321 10795 125379 10801
rect 125321 10792 125333 10795
rect 122984 10764 125333 10792
rect 122984 10752 122990 10764
rect 125321 10761 125333 10764
rect 125367 10792 125379 10795
rect 125686 10792 125692 10804
rect 125367 10764 125692 10792
rect 125367 10761 125379 10764
rect 125321 10755 125379 10761
rect 125686 10752 125692 10764
rect 125744 10752 125750 10804
rect 126701 10795 126759 10801
rect 126701 10761 126713 10795
rect 126747 10761 126759 10795
rect 130194 10792 130200 10804
rect 130155 10764 130200 10792
rect 126701 10755 126759 10761
rect 120166 10684 120172 10736
rect 120224 10724 120230 10736
rect 126716 10724 126744 10755
rect 130194 10752 130200 10764
rect 130252 10752 130258 10804
rect 136174 10792 136180 10804
rect 130304 10764 136180 10792
rect 120224 10696 126744 10724
rect 120224 10684 120230 10696
rect 126790 10684 126796 10736
rect 126848 10724 126854 10736
rect 130304 10724 130332 10764
rect 136174 10752 136180 10764
rect 136232 10752 136238 10804
rect 136729 10795 136787 10801
rect 136729 10761 136741 10795
rect 136775 10792 136787 10795
rect 136910 10792 136916 10804
rect 136775 10764 136916 10792
rect 136775 10761 136787 10764
rect 136729 10755 136787 10761
rect 136910 10752 136916 10764
rect 136968 10752 136974 10804
rect 137646 10752 137652 10804
rect 137704 10792 137710 10804
rect 138658 10792 138664 10804
rect 137704 10764 138664 10792
rect 137704 10752 137710 10764
rect 138658 10752 138664 10764
rect 138716 10752 138722 10804
rect 138750 10752 138756 10804
rect 138808 10792 138814 10804
rect 139121 10795 139179 10801
rect 139121 10792 139133 10795
rect 138808 10764 139133 10792
rect 138808 10752 138814 10764
rect 139121 10761 139133 10764
rect 139167 10761 139179 10795
rect 139121 10755 139179 10761
rect 139854 10752 139860 10804
rect 139912 10792 139918 10804
rect 140774 10792 140780 10804
rect 139912 10764 140780 10792
rect 139912 10752 139918 10764
rect 140774 10752 140780 10764
rect 140832 10752 140838 10804
rect 140961 10795 141019 10801
rect 140961 10761 140973 10795
rect 141007 10761 141019 10795
rect 140961 10755 141019 10761
rect 126848 10696 130332 10724
rect 131568 10727 131626 10733
rect 126848 10684 126854 10696
rect 131568 10693 131580 10727
rect 131614 10724 131626 10727
rect 140976 10724 141004 10755
rect 141326 10752 141332 10804
rect 141384 10792 141390 10804
rect 147306 10792 147312 10804
rect 141384 10764 147312 10792
rect 141384 10752 141390 10764
rect 147306 10752 147312 10764
rect 147364 10752 147370 10804
rect 148778 10792 148784 10804
rect 147416 10764 148784 10792
rect 131614 10696 141004 10724
rect 131614 10693 131626 10696
rect 131568 10687 131626 10693
rect 141234 10684 141240 10736
rect 141292 10724 141298 10736
rect 141789 10727 141847 10733
rect 141789 10724 141801 10727
rect 141292 10696 141801 10724
rect 141292 10684 141298 10696
rect 141789 10693 141801 10696
rect 141835 10724 141847 10727
rect 144825 10727 144883 10733
rect 144825 10724 144837 10727
rect 141835 10696 144837 10724
rect 141835 10693 141847 10696
rect 141789 10687 141847 10693
rect 144825 10693 144837 10696
rect 144871 10693 144883 10727
rect 144825 10687 144883 10693
rect 144914 10684 144920 10736
rect 144972 10724 144978 10736
rect 145898 10727 145956 10733
rect 145898 10724 145910 10727
rect 144972 10696 145910 10724
rect 144972 10684 144978 10696
rect 145898 10693 145910 10696
rect 145944 10693 145956 10727
rect 147416 10724 147444 10764
rect 148778 10752 148784 10764
rect 148836 10752 148842 10804
rect 148873 10795 148931 10801
rect 148873 10761 148885 10795
rect 148919 10792 148931 10795
rect 150250 10792 150256 10804
rect 148919 10764 150256 10792
rect 148919 10761 148931 10764
rect 148873 10755 148931 10761
rect 150250 10752 150256 10764
rect 150308 10752 150314 10804
rect 150710 10752 150716 10804
rect 150768 10792 150774 10804
rect 150805 10795 150863 10801
rect 150805 10792 150817 10795
rect 150768 10764 150817 10792
rect 150768 10752 150774 10764
rect 150805 10761 150817 10764
rect 150851 10761 150863 10795
rect 150805 10755 150863 10761
rect 150894 10752 150900 10804
rect 150952 10792 150958 10804
rect 152550 10792 152556 10804
rect 150952 10764 152556 10792
rect 150952 10752 150958 10764
rect 152550 10752 152556 10764
rect 152608 10752 152614 10804
rect 153930 10752 153936 10804
rect 153988 10792 153994 10804
rect 154574 10792 154580 10804
rect 153988 10764 154580 10792
rect 153988 10752 153994 10764
rect 154574 10752 154580 10764
rect 154632 10752 154638 10804
rect 155310 10792 155316 10804
rect 155271 10764 155316 10792
rect 155310 10752 155316 10764
rect 155368 10752 155374 10804
rect 155678 10752 155684 10804
rect 155736 10792 155742 10804
rect 157613 10795 157671 10801
rect 157613 10792 157625 10795
rect 155736 10764 157625 10792
rect 155736 10752 155742 10764
rect 157613 10761 157625 10764
rect 157659 10761 157671 10795
rect 158254 10792 158260 10804
rect 158215 10764 158260 10792
rect 157613 10755 157671 10761
rect 158254 10752 158260 10764
rect 158312 10752 158318 10804
rect 155402 10724 155408 10736
rect 145898 10687 145956 10693
rect 146036 10696 147444 10724
rect 147692 10696 150756 10724
rect 118602 10616 118608 10668
rect 118660 10656 118666 10668
rect 118901 10659 118959 10665
rect 118901 10656 118913 10659
rect 118660 10628 118913 10656
rect 118660 10616 118666 10628
rect 118901 10625 118913 10628
rect 118947 10656 118959 10659
rect 120534 10656 120540 10668
rect 118947 10628 120120 10656
rect 120495 10628 120540 10656
rect 118947 10625 118959 10628
rect 118901 10619 118959 10625
rect 119154 10588 119160 10600
rect 119115 10560 119160 10588
rect 119154 10548 119160 10560
rect 119212 10548 119218 10600
rect 120092 10588 120120 10628
rect 120534 10616 120540 10628
rect 120592 10616 120598 10668
rect 122098 10616 122104 10668
rect 122156 10665 122162 10668
rect 122156 10656 122168 10665
rect 122156 10628 122201 10656
rect 122156 10619 122168 10628
rect 122156 10616 122162 10619
rect 122282 10616 122288 10668
rect 122340 10656 122346 10668
rect 123021 10659 123079 10665
rect 123021 10656 123033 10659
rect 122340 10628 123033 10656
rect 122340 10616 122346 10628
rect 123021 10625 123033 10628
rect 123067 10625 123079 10659
rect 123021 10619 123079 10625
rect 123754 10616 123760 10668
rect 123812 10656 123818 10668
rect 124217 10659 124275 10665
rect 124217 10656 124229 10659
rect 123812 10628 124229 10656
rect 123812 10616 123818 10628
rect 124217 10625 124229 10628
rect 124263 10656 124275 10659
rect 125226 10656 125232 10668
rect 124263 10628 125232 10656
rect 124263 10625 124275 10628
rect 124217 10619 124275 10625
rect 125226 10616 125232 10628
rect 125284 10616 125290 10668
rect 125686 10616 125692 10668
rect 125744 10646 125750 10668
rect 125873 10659 125931 10665
rect 125873 10646 125885 10659
rect 125744 10625 125885 10646
rect 125919 10625 125931 10659
rect 125744 10619 125931 10625
rect 126057 10659 126115 10665
rect 126057 10625 126069 10659
rect 126103 10656 126115 10659
rect 126146 10656 126152 10668
rect 126103 10628 126152 10656
rect 126103 10625 126115 10628
rect 126057 10619 126115 10625
rect 125744 10618 125916 10619
rect 125744 10616 125750 10618
rect 126146 10616 126152 10628
rect 126204 10616 126210 10668
rect 126882 10656 126888 10668
rect 126843 10628 126888 10656
rect 126882 10616 126888 10628
rect 126940 10616 126946 10668
rect 126974 10616 126980 10668
rect 127032 10656 127038 10668
rect 127989 10659 128047 10665
rect 127989 10656 128001 10659
rect 127032 10628 128001 10656
rect 127032 10616 127038 10628
rect 127989 10625 128001 10628
rect 128035 10625 128047 10659
rect 127989 10619 128047 10625
rect 128078 10616 128084 10668
rect 128136 10656 128142 10668
rect 128354 10656 128360 10668
rect 128136 10628 128360 10656
rect 128136 10616 128142 10628
rect 128354 10616 128360 10628
rect 128412 10616 128418 10668
rect 128446 10616 128452 10668
rect 128504 10656 128510 10668
rect 128541 10659 128599 10665
rect 128541 10656 128553 10659
rect 128504 10628 128553 10656
rect 128504 10616 128510 10628
rect 128541 10625 128553 10628
rect 128587 10625 128599 10659
rect 128541 10619 128599 10625
rect 128817 10659 128875 10665
rect 128817 10625 128829 10659
rect 128863 10656 128875 10659
rect 128906 10656 128912 10668
rect 128863 10628 128912 10656
rect 128863 10625 128875 10628
rect 128817 10619 128875 10625
rect 128906 10616 128912 10628
rect 128964 10616 128970 10668
rect 130562 10616 130568 10668
rect 130620 10656 130626 10668
rect 130841 10659 130899 10665
rect 130841 10656 130853 10659
rect 130620 10628 130853 10656
rect 130620 10616 130626 10628
rect 130841 10625 130853 10628
rect 130887 10656 130899 10659
rect 130887 10628 132356 10656
rect 130887 10625 130899 10628
rect 130841 10619 130899 10625
rect 122374 10588 122380 10600
rect 120092 10560 121132 10588
rect 122335 10560 122380 10588
rect 111668 10492 116440 10520
rect 111668 10480 111674 10492
rect 110598 10452 110604 10464
rect 108868 10424 110604 10452
rect 110598 10412 110604 10424
rect 110656 10412 110662 10464
rect 110782 10452 110788 10464
rect 110743 10424 110788 10452
rect 110782 10412 110788 10424
rect 110840 10412 110846 10464
rect 111245 10455 111303 10461
rect 111245 10421 111257 10455
rect 111291 10452 111303 10455
rect 111334 10452 111340 10464
rect 111291 10424 111340 10452
rect 111291 10421 111303 10424
rect 111245 10415 111303 10421
rect 111334 10412 111340 10424
rect 111392 10412 111398 10464
rect 111426 10412 111432 10464
rect 111484 10452 111490 10464
rect 112165 10455 112223 10461
rect 112165 10452 112177 10455
rect 111484 10424 112177 10452
rect 111484 10412 111490 10424
rect 112165 10421 112177 10424
rect 112211 10452 112223 10455
rect 113450 10452 113456 10464
rect 112211 10424 113456 10452
rect 112211 10421 112223 10424
rect 112165 10415 112223 10421
rect 113450 10412 113456 10424
rect 113508 10412 113514 10464
rect 113818 10412 113824 10464
rect 113876 10452 113882 10464
rect 115293 10455 115351 10461
rect 115293 10452 115305 10455
rect 113876 10424 115305 10452
rect 113876 10412 113882 10424
rect 115293 10421 115305 10424
rect 115339 10452 115351 10455
rect 115842 10452 115848 10464
rect 115339 10424 115848 10452
rect 115339 10421 115351 10424
rect 115293 10415 115351 10421
rect 115842 10412 115848 10424
rect 115900 10412 115906 10464
rect 116412 10452 116440 10492
rect 117332 10492 118188 10520
rect 117332 10452 117360 10492
rect 116412 10424 117360 10452
rect 117866 10412 117872 10464
rect 117924 10452 117930 10464
rect 120166 10452 120172 10464
rect 117924 10424 120172 10452
rect 117924 10412 117930 10424
rect 120166 10412 120172 10424
rect 120224 10412 120230 10464
rect 120350 10452 120356 10464
rect 120311 10424 120356 10452
rect 120350 10412 120356 10424
rect 120408 10412 120414 10464
rect 120994 10452 121000 10464
rect 120955 10424 121000 10452
rect 120994 10412 121000 10424
rect 121052 10412 121058 10464
rect 121104 10452 121132 10560
rect 122374 10548 122380 10560
rect 122432 10548 122438 10600
rect 125594 10588 125600 10600
rect 122475 10560 125600 10588
rect 122475 10452 122503 10560
rect 125594 10548 125600 10560
rect 125652 10548 125658 10600
rect 131301 10591 131359 10597
rect 131301 10557 131313 10591
rect 131347 10557 131359 10591
rect 132328 10588 132356 10628
rect 132402 10616 132408 10668
rect 132460 10656 132466 10668
rect 132460 10628 136864 10656
rect 132460 10616 132466 10628
rect 136726 10588 136732 10600
rect 132328 10560 136732 10588
rect 131301 10551 131359 10557
rect 122558 10480 122564 10532
rect 122616 10520 122622 10532
rect 122616 10492 125732 10520
rect 122616 10480 122622 10492
rect 121104 10424 122503 10452
rect 122834 10412 122840 10464
rect 122892 10452 122898 10464
rect 122929 10455 122987 10461
rect 122929 10452 122941 10455
rect 122892 10424 122941 10452
rect 122892 10412 122898 10424
rect 122929 10421 122941 10424
rect 122975 10421 122987 10455
rect 123662 10452 123668 10464
rect 123623 10424 123668 10452
rect 122929 10415 122987 10421
rect 123662 10412 123668 10424
rect 123720 10412 123726 10464
rect 123754 10412 123760 10464
rect 123812 10452 123818 10464
rect 125594 10452 125600 10464
rect 123812 10424 125600 10452
rect 123812 10412 123818 10424
rect 125594 10412 125600 10424
rect 125652 10412 125658 10464
rect 125704 10452 125732 10492
rect 127066 10480 127072 10532
rect 127124 10520 127130 10532
rect 127805 10523 127863 10529
rect 127805 10520 127817 10523
rect 127124 10492 127817 10520
rect 127124 10480 127130 10492
rect 127805 10489 127817 10492
rect 127851 10489 127863 10523
rect 127805 10483 127863 10489
rect 126146 10452 126152 10464
rect 125704 10424 126152 10452
rect 126146 10412 126152 10424
rect 126204 10412 126210 10464
rect 126241 10455 126299 10461
rect 126241 10421 126253 10455
rect 126287 10452 126299 10455
rect 127526 10452 127532 10464
rect 126287 10424 127532 10452
rect 126287 10421 126299 10424
rect 126241 10415 126299 10421
rect 127526 10412 127532 10424
rect 127584 10412 127590 10464
rect 128170 10412 128176 10464
rect 128228 10452 128234 10464
rect 130194 10452 130200 10464
rect 128228 10424 130200 10452
rect 128228 10412 128234 10424
rect 130194 10412 130200 10424
rect 130252 10412 130258 10464
rect 130286 10412 130292 10464
rect 130344 10452 130350 10464
rect 131316 10452 131344 10551
rect 136726 10548 136732 10560
rect 136784 10548 136790 10600
rect 136836 10588 136864 10628
rect 138014 10616 138020 10668
rect 138072 10656 138078 10668
rect 138405 10659 138463 10665
rect 138405 10656 138417 10659
rect 138072 10628 138417 10656
rect 138072 10616 138078 10628
rect 138405 10625 138417 10628
rect 138451 10625 138463 10659
rect 138405 10619 138463 10625
rect 138661 10659 138719 10665
rect 138661 10625 138673 10659
rect 138707 10656 138719 10659
rect 138707 10628 138796 10656
rect 138707 10625 138719 10628
rect 138661 10619 138719 10625
rect 137646 10588 137652 10600
rect 136836 10560 137652 10588
rect 137646 10548 137652 10560
rect 137704 10548 137710 10600
rect 138768 10588 138796 10628
rect 140314 10616 140320 10668
rect 140372 10656 140378 10668
rect 141142 10656 141148 10668
rect 140372 10628 140636 10656
rect 141103 10628 141148 10656
rect 140372 10616 140378 10628
rect 139486 10588 139492 10600
rect 138768 10560 139492 10588
rect 139486 10548 139492 10560
rect 139544 10588 139550 10600
rect 139673 10591 139731 10597
rect 139673 10588 139685 10591
rect 139544 10560 139685 10588
rect 139544 10548 139550 10560
rect 139673 10557 139685 10560
rect 139719 10588 139731 10591
rect 140498 10588 140504 10600
rect 139719 10560 140504 10588
rect 139719 10557 139731 10560
rect 139673 10551 139731 10557
rect 140498 10548 140504 10560
rect 140556 10548 140562 10600
rect 140608 10588 140636 10628
rect 141142 10616 141148 10628
rect 141200 10616 141206 10668
rect 141326 10616 141332 10668
rect 141384 10656 141390 10668
rect 143997 10659 144055 10665
rect 143997 10656 144009 10659
rect 141384 10628 144009 10656
rect 141384 10616 141390 10628
rect 143997 10625 144009 10628
rect 144043 10625 144055 10659
rect 144178 10656 144184 10668
rect 144139 10628 144184 10656
rect 143997 10619 144055 10625
rect 144178 10616 144184 10628
rect 144236 10616 144242 10668
rect 144730 10656 144736 10668
rect 144288 10628 144736 10656
rect 144288 10588 144316 10628
rect 144730 10616 144736 10628
rect 144788 10616 144794 10668
rect 145190 10616 145196 10668
rect 145248 10656 145254 10668
rect 145653 10659 145711 10665
rect 145653 10656 145665 10659
rect 145248 10628 145665 10656
rect 145248 10616 145254 10628
rect 145653 10625 145665 10628
rect 145699 10625 145711 10659
rect 146036 10656 146064 10696
rect 145653 10619 145711 10625
rect 145760 10628 146064 10656
rect 140608 10560 144316 10588
rect 144365 10591 144423 10597
rect 144365 10557 144377 10591
rect 144411 10588 144423 10591
rect 145760 10588 145788 10628
rect 146938 10616 146944 10668
rect 146996 10656 147002 10668
rect 147692 10656 147720 10696
rect 150728 10680 150756 10696
rect 150912 10696 155408 10724
rect 146996 10628 147720 10656
rect 147760 10659 147818 10665
rect 146996 10616 147002 10628
rect 147760 10625 147772 10659
rect 147806 10656 147818 10659
rect 147806 10628 149376 10656
rect 147806 10625 147818 10628
rect 147760 10619 147818 10625
rect 144411 10560 145788 10588
rect 144411 10557 144423 10560
rect 144365 10551 144423 10557
rect 133233 10523 133291 10529
rect 133233 10520 133245 10523
rect 132236 10492 133245 10520
rect 132236 10452 132264 10492
rect 133233 10489 133245 10492
rect 133279 10520 133291 10523
rect 135625 10523 135683 10529
rect 133279 10492 134840 10520
rect 133279 10489 133291 10492
rect 133233 10483 133291 10489
rect 130344 10424 132264 10452
rect 132681 10455 132739 10461
rect 130344 10412 130350 10424
rect 132681 10421 132693 10455
rect 132727 10452 132739 10455
rect 133046 10452 133052 10464
rect 132727 10424 133052 10452
rect 132727 10421 132739 10424
rect 132681 10415 132739 10421
rect 133046 10412 133052 10424
rect 133104 10412 133110 10464
rect 133690 10452 133696 10464
rect 133651 10424 133696 10452
rect 133690 10412 133696 10424
rect 133748 10412 133754 10464
rect 134812 10461 134840 10492
rect 135625 10489 135637 10523
rect 135671 10520 135683 10523
rect 135671 10492 137416 10520
rect 135671 10489 135683 10492
rect 135625 10483 135683 10489
rect 134797 10455 134855 10461
rect 134797 10421 134809 10455
rect 134843 10452 134855 10455
rect 134978 10452 134984 10464
rect 134843 10424 134984 10452
rect 134843 10421 134855 10424
rect 134797 10415 134855 10421
rect 134978 10412 134984 10424
rect 135036 10452 135042 10464
rect 135530 10452 135536 10464
rect 135036 10424 135536 10452
rect 135036 10412 135042 10424
rect 135530 10412 135536 10424
rect 135588 10412 135594 10464
rect 136177 10455 136235 10461
rect 136177 10421 136189 10455
rect 136223 10452 136235 10455
rect 136542 10452 136548 10464
rect 136223 10424 136548 10452
rect 136223 10421 136235 10424
rect 136177 10415 136235 10421
rect 136542 10412 136548 10424
rect 136600 10412 136606 10464
rect 136634 10412 136640 10464
rect 136692 10452 136698 10464
rect 137281 10455 137339 10461
rect 137281 10452 137293 10455
rect 136692 10424 137293 10452
rect 136692 10412 136698 10424
rect 137281 10421 137293 10424
rect 137327 10421 137339 10455
rect 137388 10452 137416 10492
rect 138658 10480 138664 10532
rect 138716 10520 138722 10532
rect 138716 10492 143212 10520
rect 138716 10480 138722 10492
rect 139854 10452 139860 10464
rect 137388 10424 139860 10452
rect 137281 10415 137339 10421
rect 139854 10412 139860 10424
rect 139912 10412 139918 10464
rect 139946 10412 139952 10464
rect 140004 10452 140010 10464
rect 141326 10452 141332 10464
rect 140004 10424 141332 10452
rect 140004 10412 140010 10424
rect 141326 10412 141332 10424
rect 141384 10412 141390 10464
rect 142890 10412 142896 10464
rect 142948 10452 142954 10464
rect 143077 10455 143135 10461
rect 143077 10452 143089 10455
rect 142948 10424 143089 10452
rect 142948 10412 142954 10424
rect 143077 10421 143089 10424
rect 143123 10421 143135 10455
rect 143184 10452 143212 10492
rect 143534 10480 143540 10532
rect 143592 10520 143598 10532
rect 144380 10520 144408 10551
rect 146662 10548 146668 10600
rect 146720 10588 146726 10600
rect 147493 10591 147551 10597
rect 147493 10588 147505 10591
rect 146720 10560 147505 10588
rect 146720 10548 146726 10560
rect 147493 10557 147505 10560
rect 147539 10557 147551 10591
rect 149348 10588 149376 10628
rect 149422 10616 149428 10668
rect 149480 10656 149486 10668
rect 149609 10659 149667 10665
rect 149480 10628 149525 10656
rect 149480 10616 149486 10628
rect 149609 10625 149621 10659
rect 149655 10656 149667 10659
rect 150158 10656 150164 10668
rect 149655 10628 150164 10656
rect 149655 10625 149667 10628
rect 149609 10619 149667 10625
rect 150158 10616 150164 10628
rect 150216 10616 150222 10668
rect 150253 10659 150311 10665
rect 150253 10625 150265 10659
rect 150299 10656 150311 10659
rect 150728 10656 150848 10680
rect 150912 10656 150940 10696
rect 155402 10684 155408 10696
rect 155460 10684 155466 10736
rect 150299 10628 150572 10656
rect 150728 10652 150940 10656
rect 150820 10628 150940 10652
rect 150299 10625 150311 10628
rect 150253 10619 150311 10625
rect 150434 10588 150440 10600
rect 149348 10560 150440 10588
rect 147493 10551 147551 10557
rect 150434 10548 150440 10560
rect 150492 10548 150498 10600
rect 150544 10588 150572 10628
rect 151630 10616 151636 10668
rect 151688 10656 151694 10668
rect 151918 10659 151976 10665
rect 151918 10656 151930 10659
rect 151688 10628 151930 10656
rect 151688 10616 151694 10628
rect 151918 10625 151930 10628
rect 151964 10625 151976 10659
rect 151918 10619 151976 10625
rect 152090 10616 152096 10668
rect 152148 10656 152154 10668
rect 152185 10659 152243 10665
rect 152185 10656 152197 10659
rect 152148 10628 152197 10656
rect 152148 10616 152154 10628
rect 152185 10625 152197 10628
rect 152231 10656 152243 10659
rect 152458 10656 152464 10668
rect 152231 10628 152464 10656
rect 152231 10625 152243 10628
rect 152185 10619 152243 10625
rect 152458 10616 152464 10628
rect 152516 10616 152522 10668
rect 153758 10659 153816 10665
rect 153758 10656 153770 10659
rect 152568 10628 153770 10656
rect 152568 10588 152596 10628
rect 153758 10625 153770 10628
rect 153804 10656 153816 10659
rect 154390 10656 154396 10668
rect 153804 10628 154396 10656
rect 153804 10625 153816 10628
rect 153758 10619 153816 10625
rect 154390 10616 154396 10628
rect 154448 10616 154454 10668
rect 154666 10656 154672 10668
rect 154627 10628 154672 10656
rect 154666 10616 154672 10628
rect 154724 10616 154730 10668
rect 155957 10659 156015 10665
rect 155957 10625 155969 10659
rect 156003 10625 156015 10659
rect 156138 10656 156144 10668
rect 156099 10628 156144 10656
rect 155957 10619 156015 10625
rect 154022 10588 154028 10600
rect 150544 10560 150756 10588
rect 149974 10520 149980 10532
rect 143592 10492 144408 10520
rect 146772 10492 147536 10520
rect 143592 10480 143598 10492
rect 146772 10452 146800 10492
rect 143184 10424 146800 10452
rect 143077 10415 143135 10421
rect 146846 10412 146852 10464
rect 146904 10452 146910 10464
rect 147030 10452 147036 10464
rect 146904 10424 147036 10452
rect 146904 10412 146910 10424
rect 147030 10412 147036 10424
rect 147088 10412 147094 10464
rect 147508 10452 147536 10492
rect 148980 10492 149980 10520
rect 148980 10452 149008 10492
rect 149974 10480 149980 10492
rect 150032 10480 150038 10532
rect 150728 10520 150756 10560
rect 152209 10560 152596 10588
rect 153983 10560 154028 10588
rect 150894 10520 150900 10532
rect 150728 10492 150900 10520
rect 150894 10480 150900 10492
rect 150952 10480 150958 10532
rect 147508 10424 149008 10452
rect 149054 10412 149060 10464
rect 149112 10452 149118 10464
rect 150069 10455 150127 10461
rect 150069 10452 150081 10455
rect 149112 10424 150081 10452
rect 149112 10412 149118 10424
rect 150069 10421 150081 10424
rect 150115 10421 150127 10455
rect 150069 10415 150127 10421
rect 150250 10412 150256 10464
rect 150308 10452 150314 10464
rect 152209 10452 152237 10560
rect 154022 10548 154028 10560
rect 154080 10548 154086 10600
rect 154206 10548 154212 10600
rect 154264 10588 154270 10600
rect 154853 10591 154911 10597
rect 154853 10588 154865 10591
rect 154264 10560 154865 10588
rect 154264 10548 154270 10560
rect 154853 10557 154865 10560
rect 154899 10557 154911 10591
rect 154853 10551 154911 10557
rect 155972 10588 156000 10619
rect 156138 10616 156144 10628
rect 156196 10616 156202 10668
rect 156966 10656 156972 10668
rect 156927 10628 156972 10656
rect 156966 10616 156972 10628
rect 157024 10616 157030 10668
rect 157797 10659 157855 10665
rect 157797 10625 157809 10659
rect 157843 10656 157855 10659
rect 159082 10656 159088 10668
rect 157843 10628 159088 10656
rect 157843 10625 157855 10628
rect 157797 10619 157855 10625
rect 159082 10616 159088 10628
rect 159140 10616 159146 10668
rect 156785 10591 156843 10597
rect 156785 10588 156797 10591
rect 155972 10560 156797 10588
rect 152642 10520 152648 10532
rect 152603 10492 152648 10520
rect 152642 10480 152648 10492
rect 152700 10480 152706 10532
rect 154298 10480 154304 10532
rect 154356 10520 154362 10532
rect 155972 10520 156000 10560
rect 156785 10557 156797 10560
rect 156831 10557 156843 10591
rect 156785 10551 156843 10557
rect 154356 10492 156000 10520
rect 156325 10523 156383 10529
rect 154356 10480 154362 10492
rect 156325 10489 156337 10523
rect 156371 10520 156383 10523
rect 158438 10520 158444 10532
rect 156371 10492 158444 10520
rect 156371 10489 156383 10492
rect 156325 10483 156383 10489
rect 158438 10480 158444 10492
rect 158496 10480 158502 10532
rect 150308 10424 152237 10452
rect 150308 10412 150314 10424
rect 152274 10412 152280 10464
rect 152332 10452 152338 10464
rect 154485 10455 154543 10461
rect 154485 10452 154497 10455
rect 152332 10424 154497 10452
rect 152332 10412 152338 10424
rect 154485 10421 154497 10424
rect 154531 10421 154543 10455
rect 154485 10415 154543 10421
rect 155218 10412 155224 10464
rect 155276 10452 155282 10464
rect 155402 10452 155408 10464
rect 155276 10424 155408 10452
rect 155276 10412 155282 10424
rect 155402 10412 155408 10424
rect 155460 10452 155466 10464
rect 155862 10452 155868 10464
rect 155460 10424 155868 10452
rect 155460 10412 155466 10424
rect 155862 10412 155868 10424
rect 155920 10412 155926 10464
rect 157150 10452 157156 10464
rect 157111 10424 157156 10452
rect 157150 10412 157156 10424
rect 157208 10412 157214 10464
rect 1104 10362 158884 10384
rect 1104 10310 20672 10362
rect 20724 10310 20736 10362
rect 20788 10310 20800 10362
rect 20852 10310 20864 10362
rect 20916 10310 20928 10362
rect 20980 10310 60117 10362
rect 60169 10310 60181 10362
rect 60233 10310 60245 10362
rect 60297 10310 60309 10362
rect 60361 10310 60373 10362
rect 60425 10310 99562 10362
rect 99614 10310 99626 10362
rect 99678 10310 99690 10362
rect 99742 10310 99754 10362
rect 99806 10310 99818 10362
rect 99870 10310 139007 10362
rect 139059 10310 139071 10362
rect 139123 10310 139135 10362
rect 139187 10310 139199 10362
rect 139251 10310 139263 10362
rect 139315 10310 158884 10362
rect 1104 10288 158884 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 1995 10220 5672 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 5644 10180 5672 10220
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5776 10220 5825 10248
rect 5776 10208 5782 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 5813 10211 5871 10217
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 19472 10248
rect 9548 10208 9554 10220
rect 12621 10183 12679 10189
rect 12621 10180 12633 10183
rect 5644 10152 12633 10180
rect 12621 10149 12633 10152
rect 12667 10180 12679 10183
rect 13630 10180 13636 10192
rect 12667 10152 13636 10180
rect 12667 10149 12679 10152
rect 12621 10143 12679 10149
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 16758 10180 16764 10192
rect 15703 10152 16764 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 16758 10140 16764 10152
rect 16816 10180 16822 10192
rect 17310 10180 17316 10192
rect 16816 10152 17316 10180
rect 16816 10140 16822 10152
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 14182 10112 14188 10124
rect 12406 10084 14188 10112
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 3844 10016 3985 10044
rect 3844 10004 3850 10016
rect 3973 10013 3985 10016
rect 4019 10044 4031 10047
rect 5718 10044 5724 10056
rect 4019 10016 5724 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 10336 10016 11437 10044
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 1673 9979 1731 9985
rect 1673 9976 1685 9979
rect 1636 9948 1685 9976
rect 1636 9936 1642 9948
rect 1673 9945 1685 9948
rect 1719 9945 1731 9979
rect 1673 9939 1731 9945
rect 4240 9979 4298 9985
rect 4240 9945 4252 9979
rect 4286 9976 4298 9979
rect 4982 9976 4988 9988
rect 4286 9948 4988 9976
rect 4286 9945 4298 9948
rect 4240 9939 4298 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 10336 9985 10364 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 12406 10044 12434 10084
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 16942 10112 16948 10124
rect 16408 10084 16948 10112
rect 13078 10044 13084 10056
rect 11655 10016 12434 10044
rect 13039 10016 13084 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 10321 9979 10379 9985
rect 10321 9976 10333 9979
rect 8260 9948 10333 9976
rect 8260 9936 8266 9948
rect 10321 9945 10333 9948
rect 10367 9945 10379 9979
rect 10321 9939 10379 9945
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9976 11023 9979
rect 11624 9976 11652 10007
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 14274 10044 14280 10056
rect 14187 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10044 14338 10056
rect 15102 10044 15108 10056
rect 14332 10016 15108 10044
rect 14332 10004 14338 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 16408 10053 16436 10084
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17034 10072 17040 10124
rect 17092 10112 17098 10124
rect 18138 10112 18144 10124
rect 17092 10084 18144 10112
rect 17092 10072 17098 10084
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16666 10044 16672 10056
rect 16623 10016 16672 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 19334 10044 19340 10056
rect 17359 10016 19340 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19444 10053 19472 10220
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 23750 10248 23756 10260
rect 20128 10220 23756 10248
rect 20128 10208 20134 10220
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24578 10208 24584 10260
rect 24636 10248 24642 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 24636 10220 25421 10248
rect 24636 10208 24642 10220
rect 25409 10217 25421 10220
rect 25455 10217 25467 10251
rect 27246 10248 27252 10260
rect 25409 10211 25467 10217
rect 25976 10220 27252 10248
rect 25424 10112 25452 10211
rect 25976 10121 26004 10220
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 27338 10208 27344 10260
rect 27396 10248 27402 10260
rect 29181 10251 29239 10257
rect 27396 10220 28764 10248
rect 27396 10208 27402 10220
rect 25961 10115 26019 10121
rect 25961 10112 25973 10115
rect 25424 10084 25973 10112
rect 25961 10081 25973 10084
rect 26007 10081 26019 10115
rect 27264 10112 27292 10208
rect 28736 10180 28764 10220
rect 29181 10217 29193 10251
rect 29227 10248 29239 10251
rect 30834 10248 30840 10260
rect 29227 10220 30840 10248
rect 29227 10217 29239 10220
rect 29181 10211 29239 10217
rect 30834 10208 30840 10220
rect 30892 10208 30898 10260
rect 39390 10248 39396 10260
rect 31220 10220 39396 10248
rect 30190 10180 30196 10192
rect 28736 10152 30196 10180
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 27801 10115 27859 10121
rect 27801 10112 27813 10115
rect 27264 10084 27813 10112
rect 25961 10075 26019 10081
rect 27801 10081 27813 10084
rect 27847 10081 27859 10115
rect 27801 10075 27859 10081
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 25130 10004 25136 10056
rect 25188 10044 25194 10056
rect 29454 10044 29460 10056
rect 25188 10016 29460 10044
rect 25188 10004 25194 10016
rect 29454 10004 29460 10016
rect 29512 10004 29518 10056
rect 29546 10004 29552 10056
rect 29604 10044 29610 10056
rect 31220 10053 31248 10220
rect 39390 10208 39396 10220
rect 39448 10208 39454 10260
rect 40313 10251 40371 10257
rect 40313 10217 40325 10251
rect 40359 10248 40371 10251
rect 40402 10248 40408 10260
rect 40359 10220 40408 10248
rect 40359 10217 40371 10220
rect 40313 10211 40371 10217
rect 40402 10208 40408 10220
rect 40460 10208 40466 10260
rect 40770 10208 40776 10260
rect 40828 10248 40834 10260
rect 41046 10248 41052 10260
rect 40828 10220 41052 10248
rect 40828 10208 40834 10220
rect 41046 10208 41052 10220
rect 41104 10208 41110 10260
rect 41414 10208 41420 10260
rect 41472 10248 41478 10260
rect 44450 10248 44456 10260
rect 41472 10220 41517 10248
rect 41892 10220 44456 10248
rect 41472 10208 41478 10220
rect 33226 10140 33232 10192
rect 33284 10180 33290 10192
rect 36262 10180 36268 10192
rect 33284 10152 36268 10180
rect 33284 10140 33290 10152
rect 36262 10140 36268 10152
rect 36320 10140 36326 10192
rect 37645 10183 37703 10189
rect 37645 10149 37657 10183
rect 37691 10180 37703 10183
rect 41230 10180 41236 10192
rect 37691 10152 41236 10180
rect 37691 10149 37703 10152
rect 37645 10143 37703 10149
rect 41230 10140 41236 10152
rect 41288 10140 41294 10192
rect 41892 10180 41920 10220
rect 44450 10208 44456 10220
rect 44508 10208 44514 10260
rect 44637 10251 44695 10257
rect 44637 10217 44649 10251
rect 44683 10248 44695 10251
rect 46014 10248 46020 10260
rect 44683 10220 46020 10248
rect 44683 10217 44695 10220
rect 44637 10211 44695 10217
rect 46014 10208 46020 10220
rect 46072 10208 46078 10260
rect 46109 10251 46167 10257
rect 46109 10217 46121 10251
rect 46155 10248 46167 10251
rect 46566 10248 46572 10260
rect 46155 10220 46572 10248
rect 46155 10217 46167 10220
rect 46109 10211 46167 10217
rect 46566 10208 46572 10220
rect 46624 10208 46630 10260
rect 47486 10248 47492 10260
rect 46676 10220 47492 10248
rect 46676 10180 46704 10220
rect 47486 10208 47492 10220
rect 47544 10208 47550 10260
rect 47857 10251 47915 10257
rect 47857 10217 47869 10251
rect 47903 10248 47915 10251
rect 48682 10248 48688 10260
rect 47903 10220 48688 10248
rect 47903 10217 47915 10220
rect 47857 10211 47915 10217
rect 48682 10208 48688 10220
rect 48740 10208 48746 10260
rect 50338 10208 50344 10260
rect 50396 10248 50402 10260
rect 50433 10251 50491 10257
rect 50433 10248 50445 10251
rect 50396 10220 50445 10248
rect 50396 10208 50402 10220
rect 50433 10217 50445 10220
rect 50479 10217 50491 10251
rect 51258 10248 51264 10260
rect 51219 10220 51264 10248
rect 50433 10211 50491 10217
rect 51258 10208 51264 10220
rect 51316 10208 51322 10260
rect 52181 10251 52239 10257
rect 52181 10217 52193 10251
rect 52227 10248 52239 10251
rect 52454 10248 52460 10260
rect 52227 10220 52460 10248
rect 52227 10217 52239 10220
rect 52181 10211 52239 10217
rect 52454 10208 52460 10220
rect 52512 10208 52518 10260
rect 64230 10248 64236 10260
rect 52564 10220 64236 10248
rect 48774 10180 48780 10192
rect 41386 10152 41920 10180
rect 45572 10152 46704 10180
rect 46768 10152 48780 10180
rect 38562 10072 38568 10124
rect 38620 10112 38626 10124
rect 38841 10115 38899 10121
rect 38841 10112 38853 10115
rect 38620 10084 38853 10112
rect 38620 10072 38626 10084
rect 38841 10081 38853 10084
rect 38887 10081 38899 10115
rect 41386 10112 41414 10152
rect 45572 10121 45600 10152
rect 38841 10075 38899 10081
rect 40788 10084 41414 10112
rect 45557 10115 45615 10121
rect 31205 10047 31263 10053
rect 31205 10044 31217 10047
rect 29604 10016 31217 10044
rect 29604 10004 29610 10016
rect 31205 10013 31217 10016
rect 31251 10013 31263 10047
rect 31205 10007 31263 10013
rect 31294 10004 31300 10056
rect 31352 10044 31358 10056
rect 31849 10047 31907 10053
rect 31849 10044 31861 10047
rect 31352 10016 31861 10044
rect 31352 10004 31358 10016
rect 31849 10013 31861 10016
rect 31895 10013 31907 10047
rect 32766 10044 32772 10056
rect 32727 10016 32772 10044
rect 31849 10007 31907 10013
rect 32766 10004 32772 10016
rect 32824 10004 32830 10056
rect 33413 10047 33471 10053
rect 33413 10013 33425 10047
rect 33459 10013 33471 10047
rect 33413 10007 33471 10013
rect 33505 10047 33563 10053
rect 33505 10013 33517 10047
rect 33551 10013 33563 10047
rect 33505 10007 33563 10013
rect 33689 10047 33747 10053
rect 33689 10013 33701 10047
rect 33735 10044 33747 10047
rect 35342 10044 35348 10056
rect 33735 10016 35348 10044
rect 33735 10013 33747 10016
rect 33689 10007 33747 10013
rect 11011 9948 11652 9976
rect 11011 9945 11023 9948
rect 10965 9939 11023 9945
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 14522 9979 14580 9985
rect 14522 9976 14534 9979
rect 12584 9948 14534 9976
rect 12584 9936 12590 9948
rect 14522 9945 14534 9948
rect 14568 9945 14580 9979
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 14522 9939 14580 9945
rect 14660 9948 16221 9976
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5442 9908 5448 9920
rect 5399 9880 5448 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 8386 9908 8392 9920
rect 8347 9880 8392 9908
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 11790 9908 11796 9920
rect 11751 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 13262 9908 13268 9920
rect 13223 9880 13268 9908
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14660 9908 14688 9948
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 18506 9976 18512 9988
rect 16908 9948 18512 9976
rect 16908 9936 16914 9948
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 26206 9979 26264 9985
rect 26206 9976 26218 9979
rect 19628 9948 26218 9976
rect 17126 9908 17132 9920
rect 13596 9880 14688 9908
rect 17087 9880 17132 9908
rect 13596 9868 13602 9880
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17865 9911 17923 9917
rect 17865 9877 17877 9911
rect 17911 9908 17923 9911
rect 18417 9911 18475 9917
rect 18417 9908 18429 9911
rect 17911 9880 18429 9908
rect 17911 9877 17923 9880
rect 17865 9871 17923 9877
rect 18417 9877 18429 9880
rect 18463 9908 18475 9911
rect 19334 9908 19340 9920
rect 18463 9880 19340 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 19628 9917 19656 9948
rect 26206 9945 26218 9948
rect 26252 9945 26264 9979
rect 26206 9939 26264 9945
rect 28068 9979 28126 9985
rect 28068 9945 28080 9979
rect 28114 9976 28126 9979
rect 30960 9979 31018 9985
rect 28114 9948 30880 9976
rect 28114 9945 28126 9948
rect 28068 9939 28126 9945
rect 19613 9911 19671 9917
rect 19613 9877 19625 9911
rect 19659 9877 19671 9911
rect 20070 9908 20076 9920
rect 20031 9880 20076 9908
rect 19613 9871 19671 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 25682 9868 25688 9920
rect 25740 9908 25746 9920
rect 27341 9911 27399 9917
rect 27341 9908 27353 9911
rect 25740 9880 27353 9908
rect 25740 9868 25746 9880
rect 27341 9877 27353 9880
rect 27387 9908 27399 9911
rect 28994 9908 29000 9920
rect 27387 9880 29000 9908
rect 27387 9877 27399 9880
rect 27341 9871 27399 9877
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 29270 9868 29276 9920
rect 29328 9908 29334 9920
rect 29825 9911 29883 9917
rect 29825 9908 29837 9911
rect 29328 9880 29837 9908
rect 29328 9868 29334 9880
rect 29825 9877 29837 9880
rect 29871 9908 29883 9911
rect 30098 9908 30104 9920
rect 29871 9880 30104 9908
rect 29871 9877 29883 9880
rect 29825 9871 29883 9877
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 30852 9908 30880 9948
rect 30960 9945 30972 9979
rect 31006 9976 31018 9979
rect 31570 9976 31576 9988
rect 31006 9948 31576 9976
rect 31006 9945 31018 9948
rect 30960 9939 31018 9945
rect 31570 9936 31576 9948
rect 31628 9936 31634 9988
rect 31726 9948 32628 9976
rect 31726 9908 31754 9948
rect 32030 9908 32036 9920
rect 30852 9880 31754 9908
rect 31991 9880 32036 9908
rect 32030 9868 32036 9880
rect 32088 9868 32094 9920
rect 32600 9917 32628 9948
rect 32585 9911 32643 9917
rect 32585 9877 32597 9911
rect 32631 9877 32643 9911
rect 33428 9908 33456 10007
rect 33520 9976 33548 10007
rect 35342 10004 35348 10016
rect 35400 10004 35406 10056
rect 35894 10004 35900 10056
rect 35952 10044 35958 10056
rect 40788 10053 40816 10084
rect 45557 10081 45569 10115
rect 45603 10081 45615 10115
rect 45557 10075 45615 10081
rect 36265 10047 36323 10053
rect 36265 10044 36277 10047
rect 35952 10016 36277 10044
rect 35952 10004 35958 10016
rect 36265 10013 36277 10016
rect 36311 10013 36323 10047
rect 38105 10047 38163 10053
rect 38105 10044 38117 10047
rect 36265 10007 36323 10013
rect 36464 10016 38117 10044
rect 33520 9948 34284 9976
rect 33594 9908 33600 9920
rect 33428 9880 33600 9908
rect 32585 9871 32643 9877
rect 33594 9868 33600 9880
rect 33652 9908 33658 9920
rect 34149 9911 34207 9917
rect 34149 9908 34161 9911
rect 33652 9880 34161 9908
rect 33652 9868 33658 9880
rect 34149 9877 34161 9880
rect 34195 9877 34207 9911
rect 34256 9908 34284 9948
rect 34514 9936 34520 9988
rect 34572 9976 34578 9988
rect 36464 9976 36492 10016
rect 38105 10013 38117 10016
rect 38151 10013 38163 10047
rect 38105 10007 38163 10013
rect 40773 10047 40831 10053
rect 40773 10013 40785 10047
rect 40819 10013 40831 10047
rect 40773 10007 40831 10013
rect 34572 9948 36492 9976
rect 36532 9979 36590 9985
rect 34572 9936 34578 9948
rect 36532 9945 36544 9979
rect 36578 9976 36590 9979
rect 36630 9976 36636 9988
rect 36578 9948 36636 9976
rect 36578 9945 36590 9948
rect 36532 9939 36590 9945
rect 36630 9936 36636 9948
rect 36688 9936 36694 9988
rect 38120 9976 38148 10007
rect 41046 10004 41052 10056
rect 41104 10044 41110 10056
rect 42530 10047 42588 10053
rect 42530 10044 42542 10047
rect 41104 10016 42542 10044
rect 41104 10004 41110 10016
rect 42530 10013 42542 10016
rect 42576 10013 42588 10047
rect 42530 10007 42588 10013
rect 42702 10004 42708 10056
rect 42760 10044 42766 10056
rect 42797 10047 42855 10053
rect 42797 10044 42809 10047
rect 42760 10016 42809 10044
rect 42760 10004 42766 10016
rect 42797 10013 42809 10016
rect 42843 10013 42855 10047
rect 42797 10007 42855 10013
rect 42812 9976 42840 10007
rect 43162 10004 43168 10056
rect 43220 10044 43226 10056
rect 43530 10053 43536 10056
rect 43257 10047 43315 10053
rect 43257 10044 43269 10047
rect 43220 10016 43269 10044
rect 43220 10004 43226 10016
rect 43257 10013 43269 10016
rect 43303 10013 43315 10047
rect 43524 10044 43536 10053
rect 43491 10016 43536 10044
rect 43257 10007 43315 10013
rect 43524 10007 43536 10016
rect 43530 10004 43536 10007
rect 43588 10004 43594 10056
rect 44634 10044 44640 10056
rect 44468 10016 44640 10044
rect 44468 9976 44496 10016
rect 44634 10004 44640 10016
rect 44692 10004 44698 10056
rect 44910 10004 44916 10056
rect 44968 10044 44974 10056
rect 46106 10044 46112 10056
rect 44968 10016 46112 10044
rect 44968 10004 44974 10016
rect 46106 10004 46112 10016
rect 46164 10004 46170 10056
rect 46293 10047 46351 10053
rect 46293 10013 46305 10047
rect 46339 10044 46351 10047
rect 46768 10044 46796 10152
rect 48774 10140 48780 10152
rect 48832 10140 48838 10192
rect 48222 10112 48228 10124
rect 47688 10084 48228 10112
rect 46934 10044 46940 10056
rect 46339 10016 46796 10044
rect 46895 10016 46940 10044
rect 46339 10013 46351 10016
rect 46293 10007 46351 10013
rect 46934 10004 46940 10016
rect 46992 10004 46998 10056
rect 47121 10047 47179 10053
rect 47121 10013 47133 10047
rect 47167 10044 47179 10047
rect 47302 10044 47308 10056
rect 47167 10016 47308 10044
rect 47167 10013 47179 10016
rect 47121 10007 47179 10013
rect 47302 10004 47308 10016
rect 47360 10004 47366 10056
rect 47486 10004 47492 10056
rect 47544 10044 47550 10056
rect 47688 10053 47716 10084
rect 48222 10072 48228 10084
rect 48280 10072 48286 10124
rect 52454 10112 52460 10124
rect 49804 10084 52460 10112
rect 47673 10047 47731 10053
rect 47673 10044 47685 10047
rect 47544 10016 47685 10044
rect 47544 10004 47550 10016
rect 47673 10013 47685 10016
rect 47719 10013 47731 10047
rect 47673 10007 47731 10013
rect 47780 10016 49648 10044
rect 47780 9976 47808 10016
rect 38120 9948 42472 9976
rect 42812 9948 44496 9976
rect 44560 9948 47808 9976
rect 34974 9908 34980 9920
rect 34256 9880 34980 9908
rect 34149 9871 34207 9877
rect 34974 9868 34980 9880
rect 35032 9868 35038 9920
rect 35805 9911 35863 9917
rect 35805 9877 35817 9911
rect 35851 9908 35863 9911
rect 35894 9908 35900 9920
rect 35851 9880 35900 9908
rect 35851 9877 35863 9880
rect 35805 9871 35863 9877
rect 35894 9868 35900 9880
rect 35952 9868 35958 9920
rect 39390 9908 39396 9920
rect 39351 9880 39396 9908
rect 39390 9868 39396 9880
rect 39448 9868 39454 9920
rect 40957 9911 41015 9917
rect 40957 9877 40969 9911
rect 41003 9908 41015 9911
rect 41782 9908 41788 9920
rect 41003 9880 41788 9908
rect 41003 9877 41015 9880
rect 40957 9871 41015 9877
rect 41782 9868 41788 9880
rect 41840 9868 41846 9920
rect 42444 9908 42472 9948
rect 44560 9908 44588 9948
rect 47854 9936 47860 9988
rect 47912 9976 47918 9988
rect 49142 9976 49148 9988
rect 47912 9948 49148 9976
rect 47912 9936 47918 9948
rect 49142 9936 49148 9948
rect 49200 9936 49206 9988
rect 49510 9976 49516 9988
rect 49568 9985 49574 9988
rect 49480 9948 49516 9976
rect 49510 9936 49516 9948
rect 49568 9939 49580 9985
rect 49620 9976 49648 10016
rect 49694 10004 49700 10056
rect 49752 10044 49758 10056
rect 49804 10053 49832 10084
rect 52454 10072 52460 10084
rect 52512 10072 52518 10124
rect 49789 10047 49847 10053
rect 49789 10044 49801 10047
rect 49752 10016 49801 10044
rect 49752 10004 49758 10016
rect 49789 10013 49801 10016
rect 49835 10013 49847 10047
rect 49789 10007 49847 10013
rect 49970 10004 49976 10056
rect 50028 10044 50034 10056
rect 50617 10047 50675 10053
rect 50617 10044 50629 10047
rect 50028 10016 50629 10044
rect 50028 10004 50034 10016
rect 50617 10013 50629 10016
rect 50663 10013 50675 10047
rect 50617 10007 50675 10013
rect 51077 10047 51135 10053
rect 51077 10013 51089 10047
rect 51123 10044 51135 10047
rect 51166 10044 51172 10056
rect 51123 10016 51172 10044
rect 51123 10013 51135 10016
rect 51077 10007 51135 10013
rect 51166 10004 51172 10016
rect 51224 10004 51230 10056
rect 51442 10004 51448 10056
rect 51500 10044 51506 10056
rect 51813 10047 51871 10053
rect 51813 10044 51825 10047
rect 51500 10016 51825 10044
rect 51500 10004 51506 10016
rect 51813 10013 51825 10016
rect 51859 10013 51871 10047
rect 51994 10044 52000 10056
rect 51955 10016 52000 10044
rect 51813 10007 51871 10013
rect 51994 10004 52000 10016
rect 52052 10004 52058 10056
rect 52564 9976 52592 10220
rect 64230 10208 64236 10220
rect 64288 10208 64294 10260
rect 74810 10248 74816 10260
rect 64340 10220 74816 10248
rect 54018 10180 54024 10192
rect 53979 10152 54024 10180
rect 54018 10140 54024 10152
rect 54076 10140 54082 10192
rect 55585 10183 55643 10189
rect 55585 10149 55597 10183
rect 55631 10180 55643 10183
rect 55950 10180 55956 10192
rect 55631 10152 55956 10180
rect 55631 10149 55643 10152
rect 55585 10143 55643 10149
rect 55950 10140 55956 10152
rect 56008 10140 56014 10192
rect 56226 10180 56232 10192
rect 56187 10152 56232 10180
rect 56226 10140 56232 10152
rect 56284 10140 56290 10192
rect 56704 10152 56916 10180
rect 52638 10072 52644 10124
rect 52696 10112 52702 10124
rect 52696 10084 52741 10112
rect 52696 10072 52702 10084
rect 54386 10072 54392 10124
rect 54444 10112 54450 10124
rect 54481 10115 54539 10121
rect 54481 10112 54493 10115
rect 54444 10084 54493 10112
rect 54444 10072 54450 10084
rect 54481 10081 54493 10084
rect 54527 10081 54539 10115
rect 56704 10112 56732 10152
rect 54481 10075 54539 10081
rect 56152 10084 56732 10112
rect 56888 10112 56916 10152
rect 57054 10140 57060 10192
rect 57112 10180 57118 10192
rect 57606 10180 57612 10192
rect 57112 10152 57612 10180
rect 57112 10140 57118 10152
rect 57606 10140 57612 10152
rect 57664 10140 57670 10192
rect 57882 10180 57888 10192
rect 57843 10152 57888 10180
rect 57882 10140 57888 10152
rect 57940 10140 57946 10192
rect 58710 10140 58716 10192
rect 58768 10180 58774 10192
rect 58989 10183 59047 10189
rect 58989 10180 59001 10183
rect 58768 10152 59001 10180
rect 58768 10140 58774 10152
rect 58989 10149 59001 10152
rect 59035 10149 59047 10183
rect 58989 10143 59047 10149
rect 59814 10140 59820 10192
rect 59872 10180 59878 10192
rect 60001 10183 60059 10189
rect 60001 10180 60013 10183
rect 59872 10152 60013 10180
rect 59872 10140 59878 10152
rect 60001 10149 60013 10152
rect 60047 10149 60059 10183
rect 62022 10180 62028 10192
rect 61983 10152 62028 10180
rect 60001 10143 60059 10149
rect 62022 10140 62028 10152
rect 62080 10140 62086 10192
rect 64340 10180 64368 10220
rect 74810 10208 74816 10220
rect 74868 10208 74874 10260
rect 82633 10251 82691 10257
rect 75012 10220 82308 10248
rect 62132 10152 64368 10180
rect 60642 10112 60648 10124
rect 56888 10084 59860 10112
rect 60603 10084 60648 10112
rect 54665 10047 54723 10053
rect 54665 10044 54677 10047
rect 54220 10016 54677 10044
rect 49620 9948 52592 9976
rect 52908 9979 52966 9985
rect 52908 9945 52920 9979
rect 52954 9976 52966 9979
rect 53190 9976 53196 9988
rect 52954 9948 53196 9976
rect 52954 9945 52966 9948
rect 52908 9939 52966 9945
rect 49568 9936 49574 9939
rect 53190 9936 53196 9948
rect 53248 9936 53254 9988
rect 53282 9936 53288 9988
rect 53340 9976 53346 9988
rect 54220 9976 54248 10016
rect 54665 10013 54677 10016
rect 54711 10013 54723 10047
rect 54665 10007 54723 10013
rect 55030 10004 55036 10056
rect 55088 10044 55094 10056
rect 56045 10047 56103 10053
rect 56045 10044 56057 10047
rect 55088 10016 56057 10044
rect 55088 10004 55094 10016
rect 56045 10013 56057 10016
rect 56091 10013 56103 10047
rect 56045 10007 56103 10013
rect 53340 9948 54248 9976
rect 53340 9936 53346 9948
rect 54570 9936 54576 9988
rect 54628 9976 54634 9988
rect 56152 9976 56180 10084
rect 56686 10004 56692 10056
rect 56744 10044 56750 10056
rect 56781 10047 56839 10053
rect 56781 10044 56793 10047
rect 56744 10016 56793 10044
rect 56744 10004 56750 10016
rect 56781 10013 56793 10016
rect 56827 10044 56839 10047
rect 56870 10044 56876 10056
rect 56827 10016 56876 10044
rect 56827 10013 56839 10016
rect 56781 10007 56839 10013
rect 56870 10004 56876 10016
rect 56928 10004 56934 10056
rect 56965 10047 57023 10053
rect 56965 10013 56977 10047
rect 57011 10013 57023 10047
rect 58802 10044 58808 10056
rect 58763 10016 58808 10044
rect 56965 10007 57023 10013
rect 54628 9948 56180 9976
rect 54628 9936 54634 9948
rect 42444 9880 44588 9908
rect 45554 9868 45560 9920
rect 45612 9908 45618 9920
rect 46753 9911 46811 9917
rect 46753 9908 46765 9911
rect 45612 9880 46765 9908
rect 45612 9868 45618 9880
rect 46753 9877 46765 9880
rect 46799 9877 46811 9911
rect 48406 9908 48412 9920
rect 48367 9880 48412 9908
rect 46753 9871 46811 9877
rect 48406 9868 48412 9880
rect 48464 9868 48470 9920
rect 50614 9868 50620 9920
rect 50672 9908 50678 9920
rect 54386 9908 54392 9920
rect 50672 9880 54392 9908
rect 50672 9868 50678 9880
rect 54386 9868 54392 9880
rect 54444 9868 54450 9920
rect 54846 9908 54852 9920
rect 54807 9880 54852 9908
rect 54846 9868 54852 9880
rect 54904 9868 54910 9920
rect 54938 9868 54944 9920
rect 54996 9908 55002 9920
rect 56980 9908 57008 10007
rect 58802 10004 58808 10016
rect 58860 10004 58866 10056
rect 59832 10053 59860 10084
rect 60642 10072 60648 10084
rect 60700 10072 60706 10124
rect 59817 10047 59875 10053
rect 59817 10013 59829 10047
rect 59863 10013 59875 10047
rect 62132 10044 62160 10152
rect 68830 10140 68836 10192
rect 68888 10180 68894 10192
rect 73706 10180 73712 10192
rect 68888 10152 73712 10180
rect 68888 10140 68894 10152
rect 73706 10140 73712 10152
rect 73764 10140 73770 10192
rect 74718 10140 74724 10192
rect 74776 10180 74782 10192
rect 75012 10180 75040 10220
rect 74776 10152 75040 10180
rect 75089 10183 75147 10189
rect 74776 10140 74782 10152
rect 75089 10149 75101 10183
rect 75135 10180 75147 10183
rect 75822 10180 75828 10192
rect 75135 10152 75828 10180
rect 75135 10149 75147 10152
rect 75089 10143 75147 10149
rect 75822 10140 75828 10152
rect 75880 10140 75886 10192
rect 77297 10183 77355 10189
rect 77297 10149 77309 10183
rect 77343 10180 77355 10183
rect 77343 10152 78352 10180
rect 77343 10149 77355 10152
rect 77297 10143 77355 10149
rect 62390 10072 62396 10124
rect 62448 10112 62454 10124
rect 65242 10112 65248 10124
rect 62448 10084 63264 10112
rect 65203 10084 65248 10112
rect 62448 10072 62454 10084
rect 63034 10044 63040 10056
rect 59817 10007 59875 10013
rect 60844 10016 62160 10044
rect 62408 10016 63040 10044
rect 57698 9976 57704 9988
rect 57659 9948 57704 9976
rect 57698 9936 57704 9948
rect 57756 9936 57762 9988
rect 57790 9936 57796 9988
rect 57848 9976 57854 9988
rect 60844 9976 60872 10016
rect 57848 9948 60872 9976
rect 60912 9979 60970 9985
rect 57848 9936 57854 9948
rect 60912 9945 60924 9979
rect 60958 9945 60970 9979
rect 60912 9939 60970 9945
rect 57054 9908 57060 9920
rect 54996 9880 57060 9908
rect 54996 9868 55002 9880
rect 57054 9868 57060 9880
rect 57112 9868 57118 9920
rect 57149 9911 57207 9917
rect 57149 9877 57161 9911
rect 57195 9908 57207 9911
rect 57514 9908 57520 9920
rect 57195 9880 57520 9908
rect 57195 9877 57207 9880
rect 57149 9871 57207 9877
rect 57514 9868 57520 9880
rect 57572 9868 57578 9920
rect 57606 9868 57612 9920
rect 57664 9908 57670 9920
rect 60458 9908 60464 9920
rect 57664 9880 60464 9908
rect 57664 9868 57670 9880
rect 60458 9868 60464 9880
rect 60516 9868 60522 9920
rect 60642 9868 60648 9920
rect 60700 9908 60706 9920
rect 60936 9908 60964 9939
rect 60700 9880 60964 9908
rect 60700 9868 60706 9880
rect 61010 9868 61016 9920
rect 61068 9908 61074 9920
rect 62408 9908 62436 10016
rect 63034 10004 63040 10016
rect 63092 10004 63098 10056
rect 63236 10053 63264 10084
rect 65242 10072 65248 10084
rect 65300 10072 65306 10124
rect 67174 10112 67180 10124
rect 67135 10084 67180 10112
rect 67174 10072 67180 10084
rect 67232 10072 67238 10124
rect 67284 10084 67588 10112
rect 63221 10047 63279 10053
rect 63221 10013 63233 10047
rect 63267 10013 63279 10047
rect 63221 10007 63279 10013
rect 64690 10004 64696 10056
rect 64748 10044 64754 10056
rect 67284 10044 67312 10084
rect 64748 10016 67312 10044
rect 64748 10004 64754 10016
rect 63144 9948 63908 9976
rect 62485 9911 62543 9917
rect 62485 9908 62497 9911
rect 61068 9880 62497 9908
rect 61068 9868 61074 9880
rect 62485 9877 62497 9880
rect 62531 9877 62543 9911
rect 62485 9871 62543 9877
rect 62574 9868 62580 9920
rect 62632 9908 62638 9920
rect 63144 9908 63172 9948
rect 63402 9908 63408 9920
rect 62632 9880 63172 9908
rect 63363 9880 63408 9908
rect 62632 9868 62638 9880
rect 63402 9868 63408 9880
rect 63460 9868 63466 9920
rect 63880 9917 63908 9948
rect 63954 9936 63960 9988
rect 64012 9976 64018 9988
rect 64978 9979 65036 9985
rect 64978 9976 64990 9979
rect 64012 9948 64990 9976
rect 64012 9936 64018 9948
rect 64978 9945 64990 9948
rect 65024 9945 65036 9979
rect 64978 9939 65036 9945
rect 66714 9936 66720 9988
rect 66772 9976 66778 9988
rect 66910 9979 66968 9985
rect 66910 9976 66922 9979
rect 66772 9948 66922 9976
rect 66772 9936 66778 9948
rect 66910 9945 66922 9948
rect 66956 9945 66968 9979
rect 67560 9976 67588 10084
rect 69014 10072 69020 10124
rect 69072 10112 69078 10124
rect 69474 10112 69480 10124
rect 69072 10084 69480 10112
rect 69072 10072 69078 10084
rect 69474 10072 69480 10084
rect 69532 10112 69538 10124
rect 69532 10084 73844 10112
rect 69532 10072 69538 10084
rect 67652 10018 67864 10046
rect 71222 10044 71228 10056
rect 67652 9976 67680 10018
rect 67560 9948 67680 9976
rect 67836 9976 67864 10018
rect 71183 10016 71228 10044
rect 71222 10004 71228 10016
rect 71280 10004 71286 10056
rect 73709 10047 73767 10053
rect 73709 10013 73721 10047
rect 73755 10013 73767 10047
rect 73816 10044 73844 10084
rect 76285 10047 76343 10053
rect 76285 10044 76297 10047
rect 73816 10016 76297 10044
rect 73709 10007 73767 10013
rect 76285 10013 76297 10016
rect 76331 10013 76343 10047
rect 76285 10007 76343 10013
rect 73430 9976 73436 9988
rect 67836 9948 73436 9976
rect 66910 9939 66968 9945
rect 73430 9936 73436 9948
rect 73488 9936 73494 9988
rect 63865 9911 63923 9917
rect 63865 9877 63877 9911
rect 63911 9877 63923 9911
rect 63865 9871 63923 9877
rect 64414 9868 64420 9920
rect 64472 9908 64478 9920
rect 65797 9911 65855 9917
rect 65797 9908 65809 9911
rect 64472 9880 65809 9908
rect 64472 9868 64478 9880
rect 65797 9877 65809 9880
rect 65843 9877 65855 9911
rect 65797 9871 65855 9877
rect 66070 9868 66076 9920
rect 66128 9908 66134 9920
rect 67726 9908 67732 9920
rect 66128 9880 67732 9908
rect 66128 9868 66134 9880
rect 67726 9868 67732 9880
rect 67784 9868 67790 9920
rect 67818 9868 67824 9920
rect 67876 9908 67882 9920
rect 69569 9911 69627 9917
rect 69569 9908 69581 9911
rect 67876 9880 69581 9908
rect 67876 9868 67882 9880
rect 69569 9877 69581 9880
rect 69615 9908 69627 9911
rect 70026 9908 70032 9920
rect 69615 9880 70032 9908
rect 69615 9877 69627 9880
rect 69569 9871 69627 9877
rect 70026 9868 70032 9880
rect 70084 9908 70090 9920
rect 71774 9908 71780 9920
rect 70084 9880 71780 9908
rect 70084 9868 70090 9880
rect 71774 9868 71780 9880
rect 71832 9868 71838 9920
rect 72602 9908 72608 9920
rect 72563 9880 72608 9908
rect 72602 9868 72608 9880
rect 72660 9868 72666 9920
rect 73154 9908 73160 9920
rect 73115 9880 73160 9908
rect 73154 9868 73160 9880
rect 73212 9908 73218 9920
rect 73724 9908 73752 10007
rect 76374 10004 76380 10056
rect 76432 10044 76438 10056
rect 76650 10044 76656 10056
rect 76432 10016 76656 10044
rect 76432 10004 76438 10016
rect 76650 10004 76656 10016
rect 76708 10004 76714 10056
rect 73976 9979 74034 9985
rect 73976 9945 73988 9979
rect 74022 9976 74034 9979
rect 74718 9976 74724 9988
rect 74022 9948 74724 9976
rect 74022 9945 74034 9948
rect 73976 9939 74034 9945
rect 74718 9936 74724 9948
rect 74776 9936 74782 9988
rect 73212 9880 73752 9908
rect 73212 9868 73218 9880
rect 75178 9868 75184 9920
rect 75236 9908 75242 9920
rect 76101 9911 76159 9917
rect 76101 9908 76113 9911
rect 75236 9880 76113 9908
rect 75236 9868 75242 9880
rect 76101 9877 76113 9880
rect 76147 9877 76159 9911
rect 76101 9871 76159 9877
rect 76558 9868 76564 9920
rect 76616 9908 76622 9920
rect 77404 9908 77432 10152
rect 78324 10053 78352 10152
rect 82280 10112 82308 10220
rect 82633 10217 82645 10251
rect 82679 10248 82691 10251
rect 84102 10248 84108 10260
rect 82679 10220 84108 10248
rect 82679 10217 82691 10220
rect 82633 10211 82691 10217
rect 84102 10208 84108 10220
rect 84160 10208 84166 10260
rect 84562 10208 84568 10260
rect 84620 10248 84626 10260
rect 96801 10251 96859 10257
rect 96801 10248 96813 10251
rect 84620 10220 96813 10248
rect 84620 10208 84626 10220
rect 96801 10217 96813 10220
rect 96847 10217 96859 10251
rect 100754 10248 100760 10260
rect 96801 10211 96859 10217
rect 96908 10220 100616 10248
rect 100715 10220 100760 10248
rect 82722 10140 82728 10192
rect 82780 10180 82786 10192
rect 83090 10180 83096 10192
rect 82780 10152 83096 10180
rect 82780 10140 82786 10152
rect 83090 10140 83096 10152
rect 83148 10140 83154 10192
rect 84746 10140 84752 10192
rect 84804 10180 84810 10192
rect 84841 10183 84899 10189
rect 84841 10180 84853 10183
rect 84804 10152 84853 10180
rect 84804 10140 84810 10152
rect 84841 10149 84853 10152
rect 84887 10149 84899 10183
rect 84841 10143 84899 10149
rect 85577 10183 85635 10189
rect 85577 10149 85589 10183
rect 85623 10180 85635 10183
rect 86402 10180 86408 10192
rect 85623 10152 86408 10180
rect 85623 10149 85635 10152
rect 85577 10143 85635 10149
rect 86402 10140 86408 10152
rect 86460 10180 86466 10192
rect 86770 10180 86776 10192
rect 86460 10152 86776 10180
rect 86460 10140 86466 10152
rect 86770 10140 86776 10152
rect 86828 10140 86834 10192
rect 89714 10140 89720 10192
rect 89772 10180 89778 10192
rect 89772 10152 89817 10180
rect 89772 10140 89778 10152
rect 90542 10140 90548 10192
rect 90600 10180 90606 10192
rect 90821 10183 90879 10189
rect 90821 10180 90833 10183
rect 90600 10152 90833 10180
rect 90600 10140 90606 10152
rect 90821 10149 90833 10152
rect 90867 10149 90879 10183
rect 92842 10180 92848 10192
rect 92803 10152 92848 10180
rect 90821 10143 90879 10149
rect 92842 10140 92848 10152
rect 92900 10140 92906 10192
rect 86954 10112 86960 10124
rect 82280 10084 86960 10112
rect 86954 10072 86960 10084
rect 87012 10072 87018 10124
rect 89530 10072 89536 10124
rect 89588 10112 89594 10124
rect 93210 10112 93216 10124
rect 89588 10084 93216 10112
rect 89588 10072 89594 10084
rect 93210 10072 93216 10084
rect 93268 10072 93274 10124
rect 78309 10047 78367 10053
rect 78309 10013 78321 10047
rect 78355 10044 78367 10047
rect 80701 10047 80759 10053
rect 80701 10044 80713 10047
rect 78355 10016 80713 10044
rect 78355 10013 78367 10016
rect 78309 10007 78367 10013
rect 80701 10013 80713 10016
rect 80747 10044 80759 10047
rect 81250 10044 81256 10056
rect 80747 10016 81256 10044
rect 80747 10013 80759 10016
rect 80701 10007 80759 10013
rect 81250 10004 81256 10016
rect 81308 10004 81314 10056
rect 84205 10047 84263 10053
rect 84205 10013 84217 10047
rect 84251 10044 84263 10047
rect 84562 10044 84568 10056
rect 84251 10016 84568 10044
rect 84251 10013 84263 10016
rect 84205 10007 84263 10013
rect 84562 10004 84568 10016
rect 84620 10004 84626 10056
rect 84746 10004 84752 10056
rect 84804 10044 84810 10056
rect 85393 10047 85451 10053
rect 85393 10044 85405 10047
rect 84804 10016 85405 10044
rect 84804 10004 84810 10016
rect 85393 10013 85405 10016
rect 85439 10044 85451 10047
rect 85482 10044 85488 10056
rect 85439 10016 85488 10044
rect 85439 10013 85451 10016
rect 85393 10007 85451 10013
rect 85482 10004 85488 10016
rect 85540 10004 85546 10056
rect 89257 10047 89315 10053
rect 89257 10044 89269 10047
rect 88352 10016 89269 10044
rect 88352 9988 88380 10016
rect 89257 10013 89269 10016
rect 89303 10013 89315 10047
rect 91646 10044 91652 10056
rect 91559 10016 91652 10044
rect 89257 10007 89315 10013
rect 91646 10004 91652 10016
rect 91704 10044 91710 10056
rect 93578 10044 93584 10056
rect 91704 10016 93584 10044
rect 91704 10004 91710 10016
rect 93578 10004 93584 10016
rect 93636 10004 93642 10056
rect 94225 10047 94283 10053
rect 94225 10044 94237 10047
rect 93872 10016 94237 10044
rect 93872 9988 93900 10016
rect 94225 10013 94237 10016
rect 94271 10044 94283 10047
rect 94777 10047 94835 10053
rect 94777 10044 94789 10047
rect 94271 10016 94789 10044
rect 94271 10013 94283 10016
rect 94225 10007 94283 10013
rect 94777 10013 94789 10016
rect 94823 10044 94835 10047
rect 94866 10044 94872 10056
rect 94823 10016 94872 10044
rect 94823 10013 94835 10016
rect 94777 10007 94835 10013
rect 94866 10004 94872 10016
rect 94924 10004 94930 10056
rect 95044 10047 95102 10053
rect 95044 10013 95056 10047
rect 95090 10044 95102 10047
rect 96908 10044 96936 10220
rect 98822 10180 98828 10192
rect 98783 10152 98828 10180
rect 98822 10140 98828 10152
rect 98880 10140 98886 10192
rect 100588 10180 100616 10220
rect 100754 10208 100760 10220
rect 100812 10208 100818 10260
rect 101309 10251 101367 10257
rect 101309 10248 101321 10251
rect 101232 10220 101321 10248
rect 101122 10180 101128 10192
rect 100588 10152 101128 10180
rect 101122 10140 101128 10152
rect 101180 10140 101186 10192
rect 98362 10112 98368 10124
rect 97000 10084 98368 10112
rect 97000 10053 97028 10084
rect 98362 10072 98368 10084
rect 98420 10072 98426 10124
rect 100205 10115 100263 10121
rect 100205 10081 100217 10115
rect 100251 10112 100263 10115
rect 101232 10112 101260 10220
rect 101309 10217 101321 10220
rect 101355 10248 101367 10251
rect 102226 10248 102232 10260
rect 101355 10220 102232 10248
rect 101355 10217 101367 10220
rect 101309 10211 101367 10217
rect 102226 10208 102232 10220
rect 102284 10208 102290 10260
rect 102870 10208 102876 10260
rect 102928 10248 102934 10260
rect 104342 10248 104348 10260
rect 102928 10220 104204 10248
rect 104303 10220 104348 10248
rect 102928 10208 102934 10220
rect 101858 10180 101864 10192
rect 101819 10152 101864 10180
rect 101858 10140 101864 10152
rect 101916 10140 101922 10192
rect 104176 10180 104204 10220
rect 104342 10208 104348 10220
rect 104400 10208 104406 10260
rect 104526 10208 104532 10260
rect 104584 10248 104590 10260
rect 106826 10248 106832 10260
rect 104584 10220 106832 10248
rect 104584 10208 104590 10220
rect 106826 10208 106832 10220
rect 106884 10208 106890 10260
rect 107105 10251 107163 10257
rect 107105 10217 107117 10251
rect 107151 10248 107163 10251
rect 107562 10248 107568 10260
rect 107151 10220 107568 10248
rect 107151 10217 107163 10220
rect 107105 10211 107163 10217
rect 107562 10208 107568 10220
rect 107620 10208 107626 10260
rect 107657 10251 107715 10257
rect 107657 10217 107669 10251
rect 107703 10248 107715 10251
rect 107746 10248 107752 10260
rect 107703 10220 107752 10248
rect 107703 10217 107715 10220
rect 107657 10211 107715 10217
rect 107746 10208 107752 10220
rect 107804 10208 107810 10260
rect 112530 10248 112536 10260
rect 108040 10220 112392 10248
rect 112491 10220 112536 10248
rect 105906 10180 105912 10192
rect 104176 10152 105912 10180
rect 105906 10140 105912 10152
rect 105964 10140 105970 10192
rect 100251 10084 101260 10112
rect 103241 10115 103299 10121
rect 100251 10081 100263 10084
rect 100205 10075 100263 10081
rect 103241 10081 103253 10115
rect 103287 10112 103299 10115
rect 103422 10112 103428 10124
rect 103287 10084 103428 10112
rect 103287 10081 103299 10084
rect 103241 10075 103299 10081
rect 103422 10072 103428 10084
rect 103480 10072 103486 10124
rect 104066 10072 104072 10124
rect 104124 10112 104130 10124
rect 107470 10112 107476 10124
rect 104124 10084 107476 10112
rect 104124 10072 104130 10084
rect 107470 10072 107476 10084
rect 107528 10072 107534 10124
rect 108040 10112 108068 10220
rect 109773 10183 109831 10189
rect 109773 10149 109785 10183
rect 109819 10149 109831 10183
rect 109773 10143 109831 10149
rect 107580 10084 108068 10112
rect 109788 10112 109816 10143
rect 110690 10140 110696 10192
rect 110748 10180 110754 10192
rect 111242 10180 111248 10192
rect 110748 10152 111248 10180
rect 110748 10140 110754 10152
rect 111242 10140 111248 10152
rect 111300 10140 111306 10192
rect 112364 10180 112392 10220
rect 112530 10208 112536 10220
rect 112588 10208 112594 10260
rect 112640 10220 118464 10248
rect 112640 10180 112668 10220
rect 112364 10152 112668 10180
rect 112990 10140 112996 10192
rect 113048 10180 113054 10192
rect 113048 10152 115704 10180
rect 113048 10140 113054 10152
rect 115566 10112 115572 10124
rect 109788 10084 115572 10112
rect 95090 10016 96936 10044
rect 96985 10047 97043 10053
rect 95090 10013 95102 10016
rect 95044 10007 95102 10013
rect 96985 10013 96997 10047
rect 97031 10013 97043 10047
rect 96985 10007 97043 10013
rect 97074 10004 97080 10056
rect 97132 10044 97138 10056
rect 97813 10047 97871 10053
rect 97132 10016 97177 10044
rect 97132 10004 97138 10016
rect 97813 10013 97825 10047
rect 97859 10013 97871 10047
rect 97813 10007 97871 10013
rect 78576 9979 78634 9985
rect 78576 9945 78588 9979
rect 78622 9976 78634 9979
rect 79594 9976 79600 9988
rect 78622 9948 79600 9976
rect 78622 9945 78634 9948
rect 78576 9939 78634 9945
rect 79594 9936 79600 9948
rect 79652 9936 79658 9988
rect 81520 9979 81578 9985
rect 81520 9945 81532 9979
rect 81566 9976 81578 9979
rect 81894 9976 81900 9988
rect 81566 9948 81900 9976
rect 81566 9945 81578 9948
rect 81520 9939 81578 9945
rect 81894 9936 81900 9948
rect 81952 9936 81958 9988
rect 83016 9948 84148 9976
rect 77846 9908 77852 9920
rect 76616 9880 77432 9908
rect 77807 9880 77852 9908
rect 76616 9868 76622 9880
rect 77846 9868 77852 9880
rect 77904 9868 77910 9920
rect 79689 9911 79747 9917
rect 79689 9877 79701 9911
rect 79735 9908 79747 9911
rect 83016 9908 83044 9948
rect 79735 9880 83044 9908
rect 79735 9877 79747 9880
rect 79689 9871 79747 9877
rect 83090 9868 83096 9920
rect 83148 9908 83154 9920
rect 83148 9880 83193 9908
rect 83148 9868 83154 9880
rect 83458 9868 83464 9920
rect 83516 9908 83522 9920
rect 84013 9911 84071 9917
rect 84013 9908 84025 9911
rect 83516 9880 84025 9908
rect 83516 9868 83522 9880
rect 84013 9877 84025 9880
rect 84059 9877 84071 9911
rect 84120 9908 84148 9948
rect 84838 9936 84844 9988
rect 84896 9976 84902 9988
rect 87325 9979 87383 9985
rect 87325 9976 87337 9979
rect 84896 9948 87337 9976
rect 84896 9936 84902 9948
rect 87325 9945 87337 9948
rect 87371 9976 87383 9979
rect 88334 9976 88340 9988
rect 87371 9948 88340 9976
rect 87371 9945 87383 9948
rect 87325 9939 87383 9945
rect 88334 9936 88340 9948
rect 88392 9936 88398 9988
rect 88990 9979 89048 9985
rect 88990 9976 89002 9979
rect 88444 9948 89002 9976
rect 87690 9908 87696 9920
rect 84120 9880 87696 9908
rect 84013 9871 84071 9877
rect 87690 9868 87696 9880
rect 87748 9868 87754 9920
rect 87874 9908 87880 9920
rect 87835 9880 87880 9908
rect 87874 9868 87880 9880
rect 87932 9868 87938 9920
rect 87966 9868 87972 9920
rect 88024 9908 88030 9920
rect 88444 9908 88472 9948
rect 88990 9945 89002 9948
rect 89036 9945 89048 9979
rect 88990 9939 89048 9945
rect 90818 9936 90824 9988
rect 90876 9976 90882 9988
rect 92201 9979 92259 9985
rect 92201 9976 92213 9979
rect 90876 9948 92213 9976
rect 90876 9936 90882 9948
rect 92201 9945 92213 9948
rect 92247 9976 92259 9979
rect 93854 9976 93860 9988
rect 92247 9948 93860 9976
rect 92247 9945 92259 9948
rect 92201 9939 92259 9945
rect 93854 9936 93860 9948
rect 93912 9936 93918 9988
rect 93946 9936 93952 9988
rect 94004 9985 94010 9988
rect 94004 9976 94016 9985
rect 97828 9976 97856 10007
rect 98270 10004 98276 10056
rect 98328 10044 98334 10056
rect 107580 10044 107608 10084
rect 115566 10072 115572 10084
rect 115624 10072 115630 10124
rect 108390 10044 108396 10056
rect 98328 10016 107608 10044
rect 108351 10016 108396 10044
rect 98328 10004 98334 10016
rect 108390 10004 108396 10016
rect 108448 10044 108454 10056
rect 110233 10047 110291 10053
rect 110233 10044 110245 10047
rect 108448 10016 110245 10044
rect 108448 10004 108454 10016
rect 110233 10013 110245 10016
rect 110279 10013 110291 10047
rect 110233 10007 110291 10013
rect 110414 10004 110420 10056
rect 110472 10044 110478 10056
rect 110598 10044 110604 10056
rect 110472 10016 110604 10044
rect 110472 10004 110478 10016
rect 110598 10004 110604 10016
rect 110656 10044 110662 10056
rect 111337 10047 111395 10053
rect 111337 10044 111349 10047
rect 110656 10016 111349 10044
rect 110656 10004 110662 10016
rect 111337 10013 111349 10016
rect 111383 10044 111395 10047
rect 111518 10044 111524 10056
rect 111383 10016 111524 10044
rect 111383 10013 111395 10016
rect 111337 10007 111395 10013
rect 111518 10004 111524 10016
rect 111576 10004 111582 10056
rect 111610 10004 111616 10056
rect 111668 10044 111674 10056
rect 112898 10044 112904 10056
rect 111668 10016 112904 10044
rect 111668 10004 111674 10016
rect 112898 10004 112904 10016
rect 112956 10004 112962 10056
rect 113542 10004 113548 10056
rect 113600 10044 113606 10056
rect 114373 10047 114431 10053
rect 114373 10044 114385 10047
rect 113600 10016 114385 10044
rect 113600 10004 113606 10016
rect 114373 10013 114385 10016
rect 114419 10013 114431 10047
rect 114373 10007 114431 10013
rect 114557 10047 114615 10053
rect 114557 10013 114569 10047
rect 114603 10044 114615 10047
rect 114738 10044 114744 10056
rect 114603 10016 114744 10044
rect 114603 10013 114615 10016
rect 114557 10007 114615 10013
rect 114738 10004 114744 10016
rect 114796 10004 114802 10056
rect 115676 10053 115704 10152
rect 115842 10072 115848 10124
rect 115900 10112 115906 10124
rect 118436 10112 118464 10220
rect 118510 10208 118516 10260
rect 118568 10248 118574 10260
rect 122558 10248 122564 10260
rect 118568 10220 122564 10248
rect 118568 10208 118574 10220
rect 122558 10208 122564 10220
rect 122616 10208 122622 10260
rect 122926 10208 122932 10260
rect 122984 10248 122990 10260
rect 122984 10220 126100 10248
rect 122984 10208 122990 10220
rect 118697 10183 118755 10189
rect 118697 10149 118709 10183
rect 118743 10180 118755 10183
rect 118786 10180 118792 10192
rect 118743 10152 118792 10180
rect 118743 10149 118755 10152
rect 118697 10143 118755 10149
rect 118786 10140 118792 10152
rect 118844 10140 118850 10192
rect 118970 10140 118976 10192
rect 119028 10180 119034 10192
rect 120537 10183 120595 10189
rect 120537 10180 120549 10183
rect 119028 10152 120549 10180
rect 119028 10140 119034 10152
rect 120537 10149 120549 10152
rect 120583 10180 120595 10183
rect 121457 10183 121515 10189
rect 120583 10152 121224 10180
rect 120583 10149 120595 10152
rect 120537 10143 120595 10149
rect 120718 10112 120724 10124
rect 115900 10084 116348 10112
rect 118436 10084 120724 10112
rect 115900 10072 115906 10084
rect 115661 10047 115719 10053
rect 115661 10013 115673 10047
rect 115707 10013 115719 10047
rect 115661 10007 115719 10013
rect 115934 10004 115940 10056
rect 115992 10044 115998 10056
rect 116320 10053 116348 10084
rect 120718 10072 120724 10084
rect 120776 10072 120782 10124
rect 116121 10047 116179 10053
rect 116121 10044 116133 10047
rect 115992 10016 116133 10044
rect 115992 10004 115998 10016
rect 116121 10013 116133 10016
rect 116167 10013 116179 10047
rect 116121 10007 116179 10013
rect 116305 10047 116363 10053
rect 116305 10013 116317 10047
rect 116351 10013 116363 10047
rect 116305 10007 116363 10013
rect 117222 10004 117228 10056
rect 117280 10044 117286 10056
rect 117317 10047 117375 10053
rect 117317 10044 117329 10047
rect 117280 10016 117329 10044
rect 117280 10004 117286 10016
rect 117317 10013 117329 10016
rect 117363 10013 117375 10047
rect 118602 10044 118608 10056
rect 117317 10007 117375 10013
rect 117424 10016 118608 10044
rect 99466 9976 99472 9988
rect 94004 9948 94049 9976
rect 94148 9948 97856 9976
rect 98012 9948 99472 9976
rect 94004 9939 94016 9948
rect 94004 9936 94010 9939
rect 88024 9880 88472 9908
rect 90361 9911 90419 9917
rect 88024 9868 88030 9880
rect 90361 9877 90373 9911
rect 90407 9908 90419 9911
rect 91094 9908 91100 9920
rect 90407 9880 91100 9908
rect 90407 9877 90419 9880
rect 90361 9871 90419 9877
rect 91094 9868 91100 9880
rect 91152 9868 91158 9920
rect 92382 9868 92388 9920
rect 92440 9908 92446 9920
rect 94148 9908 94176 9948
rect 92440 9880 94176 9908
rect 92440 9868 92446 9880
rect 94866 9868 94872 9920
rect 94924 9908 94930 9920
rect 95694 9908 95700 9920
rect 94924 9880 95700 9908
rect 94924 9868 94930 9880
rect 95694 9868 95700 9880
rect 95752 9868 95758 9920
rect 96154 9908 96160 9920
rect 96115 9880 96160 9908
rect 96154 9868 96160 9880
rect 96212 9868 96218 9920
rect 98012 9917 98040 9948
rect 99466 9936 99472 9948
rect 99524 9936 99530 9988
rect 99960 9979 100018 9985
rect 99960 9945 99972 9979
rect 100006 9976 100018 9979
rect 100754 9976 100760 9988
rect 100006 9948 100760 9976
rect 100006 9945 100018 9948
rect 99960 9939 100018 9945
rect 100754 9936 100760 9948
rect 100812 9936 100818 9988
rect 101122 9936 101128 9988
rect 101180 9976 101186 9988
rect 102870 9976 102876 9988
rect 101180 9948 102876 9976
rect 101180 9936 101186 9948
rect 102870 9936 102876 9948
rect 102928 9936 102934 9988
rect 102996 9979 103054 9985
rect 102996 9945 103008 9979
rect 103042 9976 103054 9979
rect 103422 9976 103428 9988
rect 103042 9948 103428 9976
rect 103042 9945 103054 9948
rect 102996 9939 103054 9945
rect 103422 9936 103428 9948
rect 103480 9936 103486 9988
rect 103716 9948 104940 9976
rect 97997 9911 98055 9917
rect 97997 9877 98009 9911
rect 98043 9877 98055 9911
rect 97997 9871 98055 9877
rect 98086 9868 98092 9920
rect 98144 9908 98150 9920
rect 103716 9908 103744 9948
rect 98144 9880 103744 9908
rect 103793 9911 103851 9917
rect 98144 9868 98150 9880
rect 103793 9877 103805 9911
rect 103839 9908 103851 9911
rect 104526 9908 104532 9920
rect 103839 9880 104532 9908
rect 103839 9877 103851 9880
rect 103793 9871 103851 9877
rect 104526 9868 104532 9880
rect 104584 9868 104590 9920
rect 104802 9908 104808 9920
rect 104763 9880 104808 9908
rect 104802 9868 104808 9880
rect 104860 9868 104866 9920
rect 104912 9908 104940 9948
rect 104986 9936 104992 9988
rect 105044 9976 105050 9988
rect 107746 9976 107752 9988
rect 105044 9948 107752 9976
rect 105044 9936 105050 9948
rect 107746 9936 107752 9948
rect 107804 9936 107810 9988
rect 108666 9985 108672 9988
rect 108660 9939 108672 9985
rect 108724 9976 108730 9988
rect 108724 9948 108760 9976
rect 108666 9936 108672 9939
rect 108724 9936 108730 9948
rect 110322 9936 110328 9988
rect 110380 9976 110386 9988
rect 113910 9976 113916 9988
rect 110380 9948 113916 9976
rect 110380 9936 110386 9948
rect 113910 9936 113916 9948
rect 113968 9936 113974 9988
rect 115842 9936 115848 9988
rect 115900 9976 115906 9988
rect 116026 9976 116032 9988
rect 115900 9948 116032 9976
rect 115900 9936 115906 9948
rect 116026 9936 116032 9948
rect 116084 9936 116090 9988
rect 117424 9976 117452 10016
rect 118602 10004 118608 10016
rect 118660 10004 118666 10056
rect 119154 10044 119160 10056
rect 119115 10016 119160 10044
rect 119154 10004 119160 10016
rect 119212 10044 119218 10056
rect 119893 10047 119951 10053
rect 119893 10044 119905 10047
rect 119212 10016 119905 10044
rect 119212 10004 119218 10016
rect 119893 10013 119905 10016
rect 119939 10013 119951 10047
rect 121086 10044 121092 10056
rect 121047 10016 121092 10044
rect 119893 10007 119951 10013
rect 121086 10004 121092 10016
rect 121144 10004 121150 10056
rect 121196 10044 121224 10152
rect 121457 10149 121469 10183
rect 121503 10180 121515 10183
rect 122282 10180 122288 10192
rect 121503 10152 122288 10180
rect 121503 10149 121515 10152
rect 121457 10143 121515 10149
rect 122282 10140 122288 10152
rect 122340 10140 122346 10192
rect 123205 10183 123263 10189
rect 123205 10149 123217 10183
rect 123251 10180 123263 10183
rect 123386 10180 123392 10192
rect 123251 10152 123392 10180
rect 123251 10149 123263 10152
rect 123205 10143 123263 10149
rect 123386 10140 123392 10152
rect 123444 10180 123450 10192
rect 123754 10180 123760 10192
rect 123444 10152 123760 10180
rect 123444 10140 123450 10152
rect 123754 10140 123760 10152
rect 123812 10140 123818 10192
rect 126072 10180 126100 10220
rect 126146 10208 126152 10260
rect 126204 10248 126210 10260
rect 133690 10248 133696 10260
rect 126204 10220 133696 10248
rect 126204 10208 126210 10220
rect 133690 10208 133696 10220
rect 133748 10208 133754 10260
rect 133782 10208 133788 10260
rect 133840 10248 133846 10260
rect 137373 10251 137431 10257
rect 133840 10220 136956 10248
rect 133840 10208 133846 10220
rect 128170 10180 128176 10192
rect 126072 10152 128176 10180
rect 128170 10140 128176 10152
rect 128228 10140 128234 10192
rect 128354 10140 128360 10192
rect 128412 10180 128418 10192
rect 136928 10180 136956 10220
rect 137373 10217 137385 10251
rect 137419 10248 137431 10251
rect 137738 10248 137744 10260
rect 137419 10220 137744 10248
rect 137419 10217 137431 10220
rect 137373 10211 137431 10217
rect 137738 10208 137744 10220
rect 137796 10208 137802 10260
rect 140314 10248 140320 10260
rect 137848 10220 140320 10248
rect 137848 10180 137876 10220
rect 140314 10208 140320 10220
rect 140372 10208 140378 10260
rect 140498 10208 140504 10260
rect 140556 10248 140562 10260
rect 140556 10220 141372 10248
rect 140556 10208 140562 10220
rect 140866 10180 140872 10192
rect 128412 10152 128457 10180
rect 136928 10152 137876 10180
rect 139412 10152 140872 10180
rect 128412 10140 128418 10152
rect 121914 10072 121920 10124
rect 121972 10112 121978 10124
rect 122374 10112 122380 10124
rect 121972 10084 122380 10112
rect 121972 10072 121978 10084
rect 122374 10072 122380 10084
rect 122432 10072 122438 10124
rect 122742 10072 122748 10124
rect 122800 10112 122806 10124
rect 127713 10115 127771 10121
rect 122800 10084 125272 10112
rect 122800 10072 122806 10084
rect 121259 10047 121317 10053
rect 121259 10044 121271 10047
rect 121196 10016 121271 10044
rect 121259 10013 121271 10016
rect 121305 10013 121317 10047
rect 121259 10007 121317 10013
rect 122558 10004 122564 10056
rect 122616 10044 122622 10056
rect 122653 10047 122711 10053
rect 122653 10044 122665 10047
rect 122616 10016 122665 10044
rect 122616 10004 122622 10016
rect 122653 10013 122665 10016
rect 122699 10013 122711 10047
rect 122653 10007 122711 10013
rect 122834 10004 122840 10056
rect 122892 10044 122898 10056
rect 125137 10047 125195 10053
rect 125137 10044 125149 10047
rect 122892 10016 125149 10044
rect 122892 10004 122898 10016
rect 125137 10013 125149 10016
rect 125183 10013 125195 10047
rect 125244 10044 125272 10084
rect 127713 10081 127725 10115
rect 127759 10112 127771 10115
rect 128078 10112 128084 10124
rect 127759 10084 128084 10112
rect 127759 10081 127771 10084
rect 127713 10075 127771 10081
rect 128078 10072 128084 10084
rect 128136 10072 128142 10124
rect 130194 10072 130200 10124
rect 130252 10112 130258 10124
rect 132773 10115 132831 10121
rect 132773 10112 132785 10115
rect 130252 10084 132785 10112
rect 130252 10072 130258 10084
rect 132773 10081 132785 10084
rect 132819 10081 132831 10115
rect 132773 10075 132831 10081
rect 137554 10072 137560 10124
rect 137612 10112 137618 10124
rect 139412 10112 139440 10152
rect 140866 10140 140872 10152
rect 140924 10140 140930 10192
rect 141344 10180 141372 10220
rect 142154 10208 142160 10260
rect 142212 10248 142218 10260
rect 142212 10220 146616 10248
rect 142212 10208 142218 10220
rect 141344 10152 141556 10180
rect 137612 10084 139440 10112
rect 137612 10072 137618 10084
rect 125244 10016 129688 10044
rect 125137 10007 125195 10013
rect 116412 9948 117452 9976
rect 117584 9979 117642 9985
rect 108206 9908 108212 9920
rect 104912 9880 108212 9908
rect 108206 9868 108212 9880
rect 108264 9868 108270 9920
rect 108758 9868 108764 9920
rect 108816 9908 108822 9920
rect 110690 9908 110696 9920
rect 108816 9880 110696 9908
rect 108816 9868 108822 9880
rect 110690 9868 110696 9880
rect 110748 9868 110754 9920
rect 110874 9908 110880 9920
rect 110835 9880 110880 9908
rect 110874 9868 110880 9880
rect 110932 9868 110938 9920
rect 113082 9908 113088 9920
rect 113043 9880 113088 9908
rect 113082 9868 113088 9880
rect 113140 9868 113146 9920
rect 113542 9868 113548 9920
rect 113600 9908 113606 9920
rect 113637 9911 113695 9917
rect 113637 9908 113649 9911
rect 113600 9880 113649 9908
rect 113600 9868 113606 9880
rect 113637 9877 113649 9880
rect 113683 9877 113695 9911
rect 113637 9871 113695 9877
rect 114094 9868 114100 9920
rect 114152 9908 114158 9920
rect 114189 9911 114247 9917
rect 114189 9908 114201 9911
rect 114152 9880 114201 9908
rect 114152 9868 114158 9880
rect 114189 9877 114201 9880
rect 114235 9877 114247 9911
rect 115474 9908 115480 9920
rect 115435 9880 115480 9908
rect 114189 9871 114247 9877
rect 115474 9868 115480 9880
rect 115532 9868 115538 9920
rect 115566 9868 115572 9920
rect 115624 9908 115630 9920
rect 116412 9908 116440 9948
rect 117584 9945 117596 9979
rect 117630 9976 117642 9979
rect 118326 9976 118332 9988
rect 117630 9948 118332 9976
rect 117630 9945 117642 9948
rect 117584 9939 117642 9945
rect 118326 9936 118332 9948
rect 118384 9936 118390 9988
rect 120442 9976 120448 9988
rect 118666 9948 120448 9976
rect 115624 9880 116440 9908
rect 116489 9911 116547 9917
rect 115624 9868 115630 9880
rect 116489 9877 116501 9911
rect 116535 9908 116547 9911
rect 117406 9908 117412 9920
rect 116535 9880 117412 9908
rect 116535 9877 116547 9880
rect 116489 9871 116547 9877
rect 117406 9868 117412 9880
rect 117464 9868 117470 9920
rect 117958 9868 117964 9920
rect 118016 9908 118022 9920
rect 118666 9908 118694 9948
rect 120442 9936 120448 9948
rect 120500 9936 120506 9988
rect 123570 9936 123576 9988
rect 123628 9976 123634 9988
rect 123849 9979 123907 9985
rect 123849 9976 123861 9979
rect 123628 9948 123861 9976
rect 123628 9936 123634 9948
rect 123849 9945 123861 9948
rect 123895 9976 123907 9979
rect 125404 9979 125462 9985
rect 123895 9948 125364 9976
rect 123895 9945 123907 9948
rect 123849 9939 123907 9945
rect 118016 9880 118694 9908
rect 119341 9911 119399 9917
rect 118016 9868 118022 9880
rect 119341 9877 119353 9911
rect 119387 9908 119399 9911
rect 119982 9908 119988 9920
rect 119387 9880 119988 9908
rect 119387 9877 119399 9880
rect 119341 9871 119399 9877
rect 119982 9868 119988 9880
rect 120040 9868 120046 9920
rect 121546 9868 121552 9920
rect 121604 9908 121610 9920
rect 122469 9911 122527 9917
rect 122469 9908 122481 9911
rect 121604 9880 122481 9908
rect 121604 9868 121610 9880
rect 122469 9877 122481 9880
rect 122515 9877 122527 9911
rect 124398 9908 124404 9920
rect 124359 9880 124404 9908
rect 122469 9871 122527 9877
rect 124398 9868 124404 9880
rect 124456 9868 124462 9920
rect 125336 9908 125364 9948
rect 125404 9945 125416 9979
rect 125450 9976 125462 9979
rect 126977 9979 127035 9985
rect 126977 9976 126989 9979
rect 125450 9948 126989 9976
rect 125450 9945 125462 9948
rect 125404 9939 125462 9945
rect 126977 9945 126989 9948
rect 127023 9976 127035 9979
rect 129660 9976 129688 10016
rect 129734 10004 129740 10056
rect 129792 10044 129798 10056
rect 130010 10044 130016 10056
rect 129792 10016 129837 10044
rect 129971 10016 130016 10044
rect 129792 10004 129798 10016
rect 130010 10004 130016 10016
rect 130068 10004 130074 10056
rect 130473 10047 130531 10053
rect 130473 10013 130485 10047
rect 130519 10044 130531 10047
rect 130562 10044 130568 10056
rect 130519 10016 130568 10044
rect 130519 10013 130531 10016
rect 130473 10007 130531 10013
rect 130562 10004 130568 10016
rect 130620 10004 130626 10056
rect 130749 10047 130807 10053
rect 130749 10013 130761 10047
rect 130795 10044 130807 10047
rect 130930 10044 130936 10056
rect 130795 10016 130936 10044
rect 130795 10013 130807 10016
rect 130749 10007 130807 10013
rect 130930 10004 130936 10016
rect 130988 10004 130994 10056
rect 132678 10004 132684 10056
rect 132736 10044 132742 10056
rect 132957 10047 133015 10053
rect 132957 10044 132969 10047
rect 132736 10016 132969 10044
rect 132736 10004 132742 10016
rect 132957 10013 132969 10016
rect 133003 10013 133015 10047
rect 132957 10007 133015 10013
rect 134150 10004 134156 10056
rect 134208 10044 134214 10056
rect 135438 10044 135444 10056
rect 134208 10016 135444 10044
rect 134208 10004 134214 10016
rect 135438 10004 135444 10016
rect 135496 10004 135502 10056
rect 135530 10004 135536 10056
rect 135588 10044 135594 10056
rect 135993 10047 136051 10053
rect 135588 10016 135633 10044
rect 135588 10004 135594 10016
rect 135993 10013 136005 10047
rect 136039 10013 136051 10047
rect 138845 10047 138903 10053
rect 138845 10044 138857 10047
rect 135993 10007 136051 10013
rect 136652 10016 138857 10044
rect 132129 9979 132187 9985
rect 132129 9976 132141 9979
rect 127023 9948 128354 9976
rect 129660 9948 132141 9976
rect 127023 9945 127035 9948
rect 126977 9939 127035 9945
rect 126422 9908 126428 9920
rect 125336 9880 126428 9908
rect 126422 9868 126428 9880
rect 126480 9868 126486 9920
rect 126517 9911 126575 9917
rect 126517 9877 126529 9911
rect 126563 9908 126575 9911
rect 126790 9908 126796 9920
rect 126563 9880 126796 9908
rect 126563 9877 126575 9880
rect 126517 9871 126575 9877
rect 126790 9868 126796 9880
rect 126848 9868 126854 9920
rect 128326 9908 128354 9948
rect 132129 9945 132141 9948
rect 132175 9976 132187 9979
rect 132770 9976 132776 9988
rect 132175 9948 132776 9976
rect 132175 9945 132187 9948
rect 132129 9939 132187 9945
rect 132770 9936 132776 9948
rect 132828 9936 132834 9988
rect 134058 9976 134064 9988
rect 133248 9948 134064 9976
rect 133248 9908 133276 9948
rect 134058 9936 134064 9948
rect 134116 9936 134122 9988
rect 135288 9979 135346 9985
rect 135288 9945 135300 9979
rect 135334 9976 135346 9979
rect 135622 9976 135628 9988
rect 135334 9948 135628 9976
rect 135334 9945 135346 9948
rect 135288 9939 135346 9945
rect 135622 9936 135628 9948
rect 135680 9936 135686 9988
rect 133506 9908 133512 9920
rect 128326 9880 133276 9908
rect 133467 9880 133512 9908
rect 133506 9868 133512 9880
rect 133564 9868 133570 9920
rect 133966 9868 133972 9920
rect 134024 9908 134030 9920
rect 134153 9911 134211 9917
rect 134153 9908 134165 9911
rect 134024 9880 134165 9908
rect 134024 9868 134030 9880
rect 134153 9877 134165 9880
rect 134199 9877 134211 9911
rect 134153 9871 134211 9877
rect 134702 9868 134708 9920
rect 134760 9908 134766 9920
rect 136008 9908 136036 10007
rect 136266 9985 136272 9988
rect 136260 9976 136272 9985
rect 136179 9948 136272 9976
rect 136260 9939 136272 9948
rect 136324 9976 136330 9988
rect 136652 9976 136680 10016
rect 138845 10013 138857 10016
rect 138891 10044 138903 10047
rect 140038 10044 140044 10056
rect 138891 10016 140044 10044
rect 138891 10013 138903 10016
rect 138845 10007 138903 10013
rect 140038 10004 140044 10016
rect 140096 10004 140102 10056
rect 140593 10047 140651 10053
rect 140593 10013 140605 10047
rect 140639 10044 140651 10047
rect 141528 10044 141556 10152
rect 144362 10140 144368 10192
rect 144420 10180 144426 10192
rect 144914 10180 144920 10192
rect 144420 10152 144920 10180
rect 144420 10140 144426 10152
rect 144914 10140 144920 10152
rect 144972 10140 144978 10192
rect 146588 10180 146616 10220
rect 146662 10208 146668 10260
rect 146720 10248 146726 10260
rect 147030 10248 147036 10260
rect 146720 10220 147036 10248
rect 146720 10208 146726 10220
rect 147030 10208 147036 10220
rect 147088 10208 147094 10260
rect 147766 10248 147772 10260
rect 147140 10220 147772 10248
rect 147140 10180 147168 10220
rect 147766 10208 147772 10220
rect 147824 10208 147830 10260
rect 147858 10208 147864 10260
rect 147916 10248 147922 10260
rect 157337 10251 157395 10257
rect 157337 10248 157349 10251
rect 147916 10220 157349 10248
rect 147916 10208 147922 10220
rect 157337 10217 157349 10220
rect 157383 10217 157395 10251
rect 157337 10211 157395 10217
rect 146588 10152 147168 10180
rect 147306 10140 147312 10192
rect 147364 10180 147370 10192
rect 148229 10183 148287 10189
rect 148229 10180 148241 10183
rect 147364 10152 148241 10180
rect 147364 10140 147370 10152
rect 148229 10149 148241 10152
rect 148275 10149 148287 10183
rect 150250 10180 150256 10192
rect 148229 10143 148287 10149
rect 149716 10152 150256 10180
rect 145190 10112 145196 10124
rect 145151 10084 145196 10112
rect 145190 10072 145196 10084
rect 145248 10072 145254 10124
rect 146202 10072 146208 10124
rect 146260 10112 146266 10124
rect 148594 10112 148600 10124
rect 146260 10084 148600 10112
rect 146260 10072 146266 10084
rect 148594 10072 148600 10084
rect 148652 10072 148658 10124
rect 149606 10112 149612 10124
rect 149567 10084 149612 10112
rect 149606 10072 149612 10084
rect 149664 10072 149670 10124
rect 142525 10047 142583 10053
rect 142525 10044 142537 10047
rect 140639 10016 141464 10044
rect 141528 10016 142537 10044
rect 140639 10013 140651 10016
rect 140593 10007 140651 10013
rect 136324 9948 136680 9976
rect 136266 9936 136272 9939
rect 136324 9936 136330 9948
rect 136726 9936 136732 9988
rect 136784 9976 136790 9988
rect 138109 9979 138167 9985
rect 138109 9976 138121 9979
rect 136784 9948 138121 9976
rect 136784 9936 136790 9948
rect 138109 9945 138121 9948
rect 138155 9976 138167 9979
rect 139305 9979 139363 9985
rect 139305 9976 139317 9979
rect 138155 9948 139317 9976
rect 138155 9945 138167 9948
rect 138109 9939 138167 9945
rect 139305 9945 139317 9948
rect 139351 9945 139363 9979
rect 139305 9939 139363 9945
rect 139762 9936 139768 9988
rect 139820 9976 139826 9988
rect 139820 9948 140452 9976
rect 139820 9936 139826 9948
rect 136450 9908 136456 9920
rect 134760 9880 136456 9908
rect 134760 9868 134766 9880
rect 136450 9868 136456 9880
rect 136508 9868 136514 9920
rect 138198 9908 138204 9920
rect 138111 9880 138204 9908
rect 138198 9868 138204 9880
rect 138256 9908 138262 9920
rect 138658 9908 138664 9920
rect 138256 9880 138664 9908
rect 138256 9868 138262 9880
rect 138658 9868 138664 9880
rect 138716 9908 138722 9920
rect 139854 9908 139860 9920
rect 138716 9880 139860 9908
rect 138716 9868 138722 9880
rect 139854 9868 139860 9880
rect 139912 9868 139918 9920
rect 139949 9911 140007 9917
rect 139949 9877 139961 9911
rect 139995 9908 140007 9911
rect 140314 9908 140320 9920
rect 139995 9880 140320 9908
rect 139995 9877 140007 9880
rect 139949 9871 140007 9877
rect 140314 9868 140320 9880
rect 140372 9868 140378 9920
rect 140424 9917 140452 9948
rect 140774 9936 140780 9988
rect 140832 9976 140838 9988
rect 141436 9976 141464 10016
rect 142525 10013 142537 10016
rect 142571 10044 142583 10047
rect 142890 10044 142896 10056
rect 142571 10016 142896 10044
rect 142571 10013 142583 10016
rect 142525 10007 142583 10013
rect 142890 10004 142896 10016
rect 142948 10044 142954 10056
rect 143353 10047 143411 10053
rect 143353 10044 143365 10047
rect 142948 10016 143365 10044
rect 142948 10004 142954 10016
rect 143353 10013 143365 10016
rect 143399 10044 143411 10047
rect 143442 10044 143448 10056
rect 143399 10016 143448 10044
rect 143399 10013 143411 10016
rect 143353 10007 143411 10013
rect 143442 10004 143448 10016
rect 143500 10004 143506 10056
rect 144914 10044 144920 10056
rect 143552 10016 144920 10044
rect 142154 9976 142160 9988
rect 140832 9948 141280 9976
rect 141436 9948 142160 9976
rect 140832 9936 140838 9948
rect 140409 9911 140467 9917
rect 140409 9877 140421 9911
rect 140455 9877 140467 9911
rect 141142 9908 141148 9920
rect 141103 9880 141148 9908
rect 140409 9871 140467 9877
rect 141142 9868 141148 9880
rect 141200 9868 141206 9920
rect 141252 9908 141280 9948
rect 142154 9936 142160 9948
rect 142212 9936 142218 9988
rect 142280 9979 142338 9985
rect 142280 9945 142292 9979
rect 142326 9976 142338 9979
rect 143552 9976 143580 10016
rect 144914 10004 144920 10016
rect 144972 10004 144978 10056
rect 145460 10047 145518 10053
rect 145460 10013 145472 10047
rect 145506 10044 145518 10047
rect 146018 10044 146024 10056
rect 145506 10016 146024 10044
rect 145506 10013 145518 10016
rect 145460 10007 145518 10013
rect 146018 10004 146024 10016
rect 146076 10004 146082 10056
rect 147030 10004 147036 10056
rect 147088 10044 147094 10056
rect 147214 10044 147220 10056
rect 147088 10016 147220 10044
rect 147088 10004 147094 10016
rect 147214 10004 147220 10016
rect 147272 10044 147278 10056
rect 147585 10047 147643 10053
rect 147585 10044 147597 10047
rect 147272 10016 147597 10044
rect 147272 10004 147278 10016
rect 147585 10013 147597 10016
rect 147631 10013 147643 10047
rect 148042 10044 148048 10056
rect 147585 10007 147643 10013
rect 147692 10016 148048 10044
rect 142326 9948 143580 9976
rect 143620 9979 143678 9985
rect 142326 9945 142338 9948
rect 142280 9939 142338 9945
rect 143620 9945 143632 9979
rect 143666 9976 143678 9979
rect 144638 9976 144644 9988
rect 143666 9948 144644 9976
rect 143666 9945 143678 9948
rect 143620 9939 143678 9945
rect 144638 9936 144644 9948
rect 144696 9936 144702 9988
rect 146110 9936 146116 9988
rect 146168 9976 146174 9988
rect 147692 9976 147720 10016
rect 148042 10004 148048 10016
rect 148100 10004 148106 10056
rect 149330 10044 149336 10056
rect 149388 10053 149394 10056
rect 149300 10016 149336 10044
rect 149330 10004 149336 10016
rect 149388 10007 149400 10053
rect 149388 10004 149394 10007
rect 149716 9976 149744 10152
rect 150250 10140 150256 10152
rect 150308 10140 150314 10192
rect 153654 10180 153660 10192
rect 151924 10152 153660 10180
rect 150066 10072 150072 10124
rect 150124 10112 150130 10124
rect 150434 10112 150440 10124
rect 150124 10084 150440 10112
rect 150124 10072 150130 10084
rect 150434 10072 150440 10084
rect 150492 10072 150498 10124
rect 151924 10121 151952 10152
rect 153654 10140 153660 10152
rect 153712 10140 153718 10192
rect 153838 10180 153844 10192
rect 153799 10152 153844 10180
rect 153838 10140 153844 10152
rect 153896 10140 153902 10192
rect 156230 10180 156236 10192
rect 155236 10152 156236 10180
rect 151909 10115 151967 10121
rect 151372 10084 151584 10112
rect 151372 10044 151400 10084
rect 146168 9948 147720 9976
rect 147784 9948 149744 9976
rect 149900 10016 151400 10044
rect 151449 10047 151507 10053
rect 146168 9936 146174 9948
rect 144086 9908 144092 9920
rect 141252 9880 144092 9908
rect 144086 9868 144092 9880
rect 144144 9868 144150 9920
rect 144270 9868 144276 9920
rect 144328 9908 144334 9920
rect 144730 9908 144736 9920
rect 144328 9880 144736 9908
rect 144328 9868 144334 9880
rect 144730 9868 144736 9880
rect 144788 9868 144794 9920
rect 144822 9868 144828 9920
rect 144880 9908 144886 9920
rect 145466 9908 145472 9920
rect 144880 9880 145472 9908
rect 144880 9868 144886 9880
rect 145466 9868 145472 9880
rect 145524 9868 145530 9920
rect 146573 9911 146631 9917
rect 146573 9877 146585 9911
rect 146619 9908 146631 9911
rect 147784 9908 147812 9948
rect 146619 9880 147812 9908
rect 146619 9877 146631 9880
rect 146573 9871 146631 9877
rect 147858 9868 147864 9920
rect 147916 9908 147922 9920
rect 149900 9908 149928 10016
rect 151449 10013 151461 10047
rect 151495 10013 151507 10047
rect 151556 10044 151584 10084
rect 151909 10081 151921 10115
rect 151955 10081 151967 10115
rect 153930 10112 153936 10124
rect 151909 10075 151967 10081
rect 152016 10084 153936 10112
rect 152016 10044 152044 10084
rect 153930 10072 153936 10084
rect 153988 10072 153994 10124
rect 155236 10112 155264 10152
rect 156230 10140 156236 10152
rect 156288 10140 156294 10192
rect 155144 10084 155264 10112
rect 151556 10016 152044 10044
rect 152093 10047 152151 10053
rect 151449 10007 151507 10013
rect 152093 10013 152105 10047
rect 152139 10013 152151 10047
rect 152093 10007 152151 10013
rect 152277 10047 152335 10053
rect 152277 10013 152289 10047
rect 152323 10044 152335 10047
rect 154666 10044 154672 10056
rect 152323 10016 154672 10044
rect 152323 10013 152335 10016
rect 152277 10007 152335 10013
rect 150250 9936 150256 9988
rect 150308 9976 150314 9988
rect 151182 9979 151240 9985
rect 151182 9976 151194 9979
rect 150308 9948 151194 9976
rect 150308 9936 150314 9948
rect 151182 9945 151194 9948
rect 151228 9976 151240 9979
rect 151354 9976 151360 9988
rect 151228 9948 151360 9976
rect 151228 9945 151240 9948
rect 151182 9939 151240 9945
rect 151354 9936 151360 9948
rect 151412 9936 151418 9988
rect 151464 9976 151492 10007
rect 151998 9976 152004 9988
rect 151464 9948 152004 9976
rect 151998 9936 152004 9948
rect 152056 9936 152062 9988
rect 150066 9908 150072 9920
rect 147916 9880 149928 9908
rect 150027 9880 150072 9908
rect 147916 9868 147922 9880
rect 150066 9868 150072 9880
rect 150124 9868 150130 9920
rect 150710 9868 150716 9920
rect 150768 9908 150774 9920
rect 150894 9908 150900 9920
rect 150768 9880 150900 9908
rect 150768 9868 150774 9880
rect 150894 9868 150900 9880
rect 150952 9868 150958 9920
rect 151446 9868 151452 9920
rect 151504 9908 151510 9920
rect 152108 9908 152136 10007
rect 154666 10004 154672 10016
rect 154724 10004 154730 10056
rect 154965 10047 155023 10053
rect 154965 10044 154977 10047
rect 154776 10016 154977 10044
rect 154776 9976 154804 10016
rect 154965 10013 154977 10016
rect 155011 10044 155023 10047
rect 155144 10044 155172 10084
rect 155402 10072 155408 10124
rect 155460 10112 155466 10124
rect 155681 10115 155739 10121
rect 155681 10112 155693 10115
rect 155460 10084 155693 10112
rect 155460 10072 155466 10084
rect 155681 10081 155693 10084
rect 155727 10081 155739 10115
rect 155681 10075 155739 10081
rect 156049 10115 156107 10121
rect 156049 10081 156061 10115
rect 156095 10112 156107 10115
rect 157702 10112 157708 10124
rect 156095 10084 157708 10112
rect 156095 10081 156107 10084
rect 156049 10075 156107 10081
rect 157702 10072 157708 10084
rect 157760 10072 157766 10124
rect 155011 10016 155172 10044
rect 155221 10047 155279 10053
rect 155011 10013 155023 10016
rect 154965 10007 155023 10013
rect 155221 10013 155233 10047
rect 155267 10044 155279 10047
rect 155267 10016 155356 10044
rect 155267 10013 155279 10016
rect 155221 10007 155279 10013
rect 152200 9948 154804 9976
rect 152200 9920 152228 9948
rect 151504 9880 152136 9908
rect 151504 9868 151510 9880
rect 152182 9868 152188 9920
rect 152240 9868 152246 9920
rect 152274 9868 152280 9920
rect 152332 9908 152338 9920
rect 152737 9911 152795 9917
rect 152737 9908 152749 9911
rect 152332 9880 152749 9908
rect 152332 9868 152338 9880
rect 152737 9877 152749 9880
rect 152783 9877 152795 9911
rect 152737 9871 152795 9877
rect 154022 9868 154028 9920
rect 154080 9908 154086 9920
rect 155328 9908 155356 10016
rect 155770 10004 155776 10056
rect 155828 10044 155834 10056
rect 155865 10047 155923 10053
rect 155865 10044 155877 10047
rect 155828 10016 155877 10044
rect 155828 10004 155834 10016
rect 155865 10013 155877 10016
rect 155911 10013 155923 10047
rect 155865 10007 155923 10013
rect 155954 10004 155960 10056
rect 156012 10044 156018 10056
rect 156598 10044 156604 10056
rect 156012 10016 156604 10044
rect 156012 10004 156018 10016
rect 156598 10004 156604 10016
rect 156656 10004 156662 10056
rect 156693 10047 156751 10053
rect 156693 10013 156705 10047
rect 156739 10013 156751 10047
rect 157518 10044 157524 10056
rect 157479 10016 157524 10044
rect 156693 10007 156751 10013
rect 154080 9880 155356 9908
rect 154080 9868 154086 9880
rect 155402 9868 155408 9920
rect 155460 9908 155466 9920
rect 156708 9908 156736 10007
rect 157518 10004 157524 10016
rect 157576 10004 157582 10056
rect 155460 9880 156736 9908
rect 156877 9911 156935 9917
rect 155460 9868 155466 9880
rect 156877 9877 156889 9911
rect 156923 9908 156935 9911
rect 157886 9908 157892 9920
rect 156923 9880 157892 9908
rect 156923 9877 156935 9880
rect 156877 9871 156935 9877
rect 157886 9868 157892 9880
rect 157944 9868 157950 9920
rect 1104 9818 159043 9840
rect 1104 9766 40394 9818
rect 40446 9766 40458 9818
rect 40510 9766 40522 9818
rect 40574 9766 40586 9818
rect 40638 9766 40650 9818
rect 40702 9766 79839 9818
rect 79891 9766 79903 9818
rect 79955 9766 79967 9818
rect 80019 9766 80031 9818
rect 80083 9766 80095 9818
rect 80147 9766 119284 9818
rect 119336 9766 119348 9818
rect 119400 9766 119412 9818
rect 119464 9766 119476 9818
rect 119528 9766 119540 9818
rect 119592 9766 158729 9818
rect 158781 9766 158793 9818
rect 158845 9766 158857 9818
rect 158909 9766 158921 9818
rect 158973 9766 158985 9818
rect 159037 9766 159043 9818
rect 1104 9744 159043 9766
rect 1578 9704 1584 9716
rect 1539 9676 1584 9704
rect 1578 9664 1584 9676
rect 1636 9664 1642 9716
rect 5718 9704 5724 9716
rect 5679 9676 5724 9704
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 29086 9704 29092 9716
rect 5828 9676 29092 9704
rect 5166 9596 5172 9648
rect 5224 9636 5230 9648
rect 5828 9636 5856 9676
rect 29086 9664 29092 9676
rect 29144 9664 29150 9716
rect 29454 9664 29460 9716
rect 29512 9704 29518 9716
rect 31294 9704 31300 9716
rect 29512 9676 31300 9704
rect 29512 9664 29518 9676
rect 5224 9608 5856 9636
rect 5224 9596 5230 9608
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 10100 9608 11989 9636
rect 10100 9596 10106 9608
rect 11977 9605 11989 9608
rect 12023 9636 12035 9639
rect 13446 9636 13452 9648
rect 12023 9608 13452 9636
rect 12023 9605 12035 9608
rect 11977 9599 12035 9605
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 14274 9636 14280 9648
rect 13556 9608 14280 9636
rect 3786 9568 3792 9580
rect 3747 9540 3792 9568
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4056 9571 4114 9577
rect 4056 9537 4068 9571
rect 4102 9568 4114 9571
rect 5718 9568 5724 9580
rect 4102 9540 5724 9568
rect 4102 9537 4114 9540
rect 4056 9531 4114 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 13556 9577 13584 9608
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 15378 9636 15384 9648
rect 15339 9608 15384 9636
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 17770 9636 17776 9648
rect 16684 9608 17776 9636
rect 16684 9580 16712 9608
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 19334 9636 19340 9648
rect 19247 9608 19340 9636
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12400 9540 12541 9568
rect 12400 9528 12406 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 13808 9571 13866 9577
rect 13808 9537 13820 9571
rect 13854 9568 13866 9571
rect 14090 9568 14096 9580
rect 13854 9540 14096 9568
rect 13854 9537 13866 9540
rect 13808 9531 13866 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 15562 9568 15568 9580
rect 14240 9540 14964 9568
rect 15523 9540 15568 9568
rect 14240 9528 14246 9540
rect 14936 9441 14964 9540
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 15746 9568 15752 9580
rect 15707 9540 15752 9568
rect 15746 9528 15752 9540
rect 15804 9568 15810 9580
rect 16666 9568 16672 9580
rect 15804 9540 16672 9568
rect 15804 9528 15810 9540
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17218 9568 17224 9580
rect 17179 9540 17224 9568
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 19260 9577 19288 9608
rect 19334 9596 19340 9608
rect 19392 9636 19398 9648
rect 20530 9636 20536 9648
rect 19392 9608 20536 9636
rect 19392 9596 19398 9608
rect 20530 9596 20536 9608
rect 20588 9636 20594 9648
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 20588 9608 21097 9636
rect 20588 9596 20594 9608
rect 21085 9605 21097 9608
rect 21131 9605 21143 9639
rect 21085 9599 21143 9605
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 28362 9639 28420 9645
rect 28362 9636 28374 9639
rect 23440 9608 28374 9636
rect 23440 9596 23446 9608
rect 28362 9605 28374 9608
rect 28408 9605 28420 9639
rect 28362 9599 28420 9605
rect 28626 9596 28632 9648
rect 28684 9636 28690 9648
rect 30650 9636 30656 9648
rect 28684 9608 30656 9636
rect 28684 9596 28690 9608
rect 30650 9596 30656 9608
rect 30708 9596 30714 9648
rect 30944 9645 30972 9676
rect 31294 9664 31300 9676
rect 31352 9664 31358 9716
rect 31662 9704 31668 9716
rect 31623 9676 31668 9704
rect 31662 9664 31668 9676
rect 31720 9664 31726 9716
rect 35805 9707 35863 9713
rect 35805 9673 35817 9707
rect 35851 9704 35863 9707
rect 35894 9704 35900 9716
rect 35851 9676 35900 9704
rect 35851 9673 35863 9676
rect 35805 9667 35863 9673
rect 30929 9639 30987 9645
rect 30929 9605 30941 9639
rect 30975 9605 30987 9639
rect 32030 9636 32036 9648
rect 30929 9599 30987 9605
rect 31496 9608 32036 9636
rect 18989 9571 19047 9577
rect 18989 9537 19001 9571
rect 19035 9568 19047 9571
rect 19245 9571 19303 9577
rect 19035 9540 19196 9568
rect 19035 9537 19047 9540
rect 18989 9531 19047 9537
rect 15010 9460 15016 9512
rect 15068 9500 15074 9512
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 15068 9472 16221 9500
rect 15068 9460 15074 9472
rect 16209 9469 16221 9472
rect 16255 9500 16267 9503
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16255 9472 17049 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 17037 9469 17049 9472
rect 17083 9469 17095 9503
rect 19168 9500 19196 9540
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 19484 9540 19717 9568
rect 19484 9528 19490 9540
rect 19705 9537 19717 9540
rect 19751 9537 19763 9571
rect 19886 9568 19892 9580
rect 19847 9540 19892 9568
rect 19705 9531 19763 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 26073 9571 26131 9577
rect 26073 9537 26085 9571
rect 26119 9568 26131 9571
rect 26878 9568 26884 9580
rect 26119 9540 26884 9568
rect 26119 9537 26131 9540
rect 26073 9531 26131 9537
rect 26878 9528 26884 9540
rect 26936 9528 26942 9580
rect 29356 9571 29414 9577
rect 29356 9537 29368 9571
rect 29402 9568 29414 9571
rect 30742 9568 30748 9580
rect 29402 9540 30748 9568
rect 29402 9537 29414 9540
rect 29356 9531 29414 9537
rect 30742 9528 30748 9540
rect 30800 9528 30806 9580
rect 31496 9577 31524 9608
rect 32030 9596 32036 9608
rect 32088 9596 32094 9648
rect 34238 9636 34244 9648
rect 32692 9608 34244 9636
rect 32692 9577 32720 9608
rect 34238 9596 34244 9608
rect 34296 9636 34302 9648
rect 35820 9636 35848 9667
rect 35894 9664 35900 9676
rect 35952 9704 35958 9716
rect 36722 9704 36728 9716
rect 35952 9676 36728 9704
rect 35952 9664 35958 9676
rect 36722 9664 36728 9676
rect 36780 9704 36786 9716
rect 36817 9707 36875 9713
rect 36817 9704 36829 9707
rect 36780 9676 36829 9704
rect 36780 9664 36786 9676
rect 36817 9673 36829 9676
rect 36863 9704 36875 9707
rect 38654 9704 38660 9716
rect 36863 9676 38660 9704
rect 36863 9673 36875 9676
rect 36817 9667 36875 9673
rect 38654 9664 38660 9676
rect 38712 9664 38718 9716
rect 42812 9676 43576 9704
rect 34296 9608 35848 9636
rect 34296 9596 34302 9608
rect 38562 9596 38568 9648
rect 38620 9596 38626 9648
rect 38672 9636 38700 9664
rect 39390 9636 39396 9648
rect 38672 9608 39396 9636
rect 31481 9571 31539 9577
rect 31481 9537 31493 9571
rect 31527 9537 31539 9571
rect 32677 9571 32735 9577
rect 32677 9568 32689 9571
rect 31481 9531 31539 9537
rect 31726 9540 32689 9568
rect 19518 9500 19524 9512
rect 19168 9472 19524 9500
rect 17037 9463 17095 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 20070 9500 20076 9512
rect 20031 9472 20076 9500
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 26326 9500 26332 9512
rect 26287 9472 26332 9500
rect 26326 9460 26332 9472
rect 26384 9460 26390 9512
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9469 28687 9503
rect 29086 9500 29092 9512
rect 29047 9472 29092 9500
rect 28629 9463 28687 9469
rect 14921 9435 14979 9441
rect 14921 9401 14933 9435
rect 14967 9432 14979 9435
rect 19794 9432 19800 9444
rect 14967 9404 18000 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 8018 9364 8024 9376
rect 5215 9336 8024 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 12713 9367 12771 9373
rect 12713 9333 12725 9367
rect 12759 9364 12771 9367
rect 14458 9364 14464 9376
rect 12759 9336 14464 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 17552 9336 17877 9364
rect 17552 9324 17558 9336
rect 17865 9333 17877 9336
rect 17911 9333 17923 9367
rect 17972 9364 18000 9404
rect 19260 9404 19800 9432
rect 19260 9364 19288 9404
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 27062 9392 27068 9444
rect 27120 9432 27126 9444
rect 27249 9435 27307 9441
rect 27249 9432 27261 9435
rect 27120 9404 27261 9432
rect 27120 9392 27126 9404
rect 27249 9401 27261 9404
rect 27295 9401 27307 9435
rect 27249 9395 27307 9401
rect 17972 9336 19288 9364
rect 17865 9327 17923 9333
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 20625 9367 20683 9373
rect 20625 9364 20637 9367
rect 19944 9336 20637 9364
rect 19944 9324 19950 9336
rect 20625 9333 20637 9336
rect 20671 9364 20683 9367
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 20671 9336 24961 9364
rect 20671 9333 20683 9336
rect 20625 9327 20683 9333
rect 24949 9333 24961 9336
rect 24995 9364 25007 9367
rect 26510 9364 26516 9376
rect 24995 9336 26516 9364
rect 24995 9333 25007 9336
rect 24949 9327 25007 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 27706 9324 27712 9376
rect 27764 9364 27770 9376
rect 28644 9364 28672 9463
rect 29086 9460 29092 9472
rect 29144 9460 29150 9512
rect 31018 9460 31024 9512
rect 31076 9500 31082 9512
rect 31726 9500 31754 9540
rect 32677 9537 32689 9540
rect 32723 9537 32735 9571
rect 32677 9531 32735 9537
rect 32944 9571 33002 9577
rect 32944 9537 32956 9571
rect 32990 9568 33002 9571
rect 33318 9568 33324 9580
rect 32990 9540 33324 9568
rect 32990 9537 33002 9540
rect 32944 9531 33002 9537
rect 33318 9528 33324 9540
rect 33376 9528 33382 9580
rect 34514 9568 34520 9580
rect 34475 9540 34520 9568
rect 34514 9528 34520 9540
rect 34572 9528 34578 9580
rect 38580 9568 38608 9596
rect 38948 9577 38976 9608
rect 39390 9596 39396 9608
rect 39448 9636 39454 9648
rect 39577 9639 39635 9645
rect 39577 9636 39589 9639
rect 39448 9608 39589 9636
rect 39448 9596 39454 9608
rect 39577 9605 39589 9608
rect 39623 9605 39635 9639
rect 40218 9636 40224 9648
rect 40179 9608 40224 9636
rect 39577 9599 39635 9605
rect 34624 9540 38608 9568
rect 38677 9571 38735 9577
rect 31076 9472 31754 9500
rect 31076 9460 31082 9472
rect 33870 9460 33876 9512
rect 33928 9500 33934 9512
rect 34624 9500 34652 9540
rect 38677 9537 38689 9571
rect 38723 9568 38735 9571
rect 38933 9571 38991 9577
rect 38723 9540 38884 9568
rect 38723 9537 38735 9540
rect 38677 9531 38735 9537
rect 33928 9472 34652 9500
rect 38856 9500 38884 9540
rect 38933 9537 38945 9571
rect 38979 9537 38991 9571
rect 39592 9568 39620 9599
rect 40218 9596 40224 9608
rect 40276 9596 40282 9648
rect 40954 9645 40960 9648
rect 40948 9636 40960 9645
rect 40915 9608 40960 9636
rect 40948 9599 40960 9608
rect 40954 9596 40960 9599
rect 41012 9596 41018 9648
rect 42812 9636 42840 9676
rect 41386 9608 42840 9636
rect 40681 9571 40739 9577
rect 40681 9568 40693 9571
rect 39592 9540 40693 9568
rect 38933 9531 38991 9537
rect 40681 9537 40693 9540
rect 40727 9537 40739 9571
rect 41386 9568 41414 9608
rect 42886 9596 42892 9648
rect 42944 9636 42950 9648
rect 43410 9639 43468 9645
rect 43410 9636 43422 9639
rect 42944 9608 43422 9636
rect 42944 9596 42950 9608
rect 43410 9605 43422 9608
rect 43456 9605 43468 9639
rect 43548 9636 43576 9676
rect 45186 9664 45192 9716
rect 45244 9704 45250 9716
rect 47118 9704 47124 9716
rect 45244 9676 47124 9704
rect 45244 9664 45250 9676
rect 47118 9664 47124 9676
rect 47176 9664 47182 9716
rect 47213 9707 47271 9713
rect 47213 9673 47225 9707
rect 47259 9704 47271 9707
rect 47762 9704 47768 9716
rect 47259 9676 47768 9704
rect 47259 9673 47271 9676
rect 47213 9667 47271 9673
rect 47762 9664 47768 9676
rect 47820 9664 47826 9716
rect 48222 9664 48228 9716
rect 48280 9664 48286 9716
rect 49878 9664 49884 9716
rect 49936 9704 49942 9716
rect 54202 9704 54208 9716
rect 49936 9676 54208 9704
rect 49936 9664 49942 9676
rect 54202 9664 54208 9676
rect 54260 9664 54266 9716
rect 55953 9707 56011 9713
rect 55953 9704 55965 9707
rect 54404 9676 55965 9704
rect 48130 9636 48136 9648
rect 43548 9608 48136 9636
rect 43410 9599 43468 9605
rect 48130 9596 48136 9608
rect 48188 9596 48194 9648
rect 48240 9636 48268 9664
rect 49329 9639 49387 9645
rect 49329 9636 49341 9639
rect 48240 9608 49341 9636
rect 49329 9605 49341 9608
rect 49375 9636 49387 9639
rect 49694 9636 49700 9648
rect 49375 9608 49700 9636
rect 49375 9605 49387 9608
rect 49329 9599 49387 9605
rect 49694 9596 49700 9608
rect 49752 9596 49758 9648
rect 50614 9636 50620 9648
rect 50356 9608 50620 9636
rect 40681 9531 40739 9537
rect 40788 9540 41414 9568
rect 40034 9500 40040 9512
rect 38856 9472 40040 9500
rect 33928 9460 33934 9472
rect 40034 9460 40040 9472
rect 40092 9460 40098 9512
rect 40788 9500 40816 9540
rect 41506 9528 41512 9580
rect 41564 9568 41570 9580
rect 41782 9568 41788 9580
rect 41564 9540 41788 9568
rect 41564 9528 41570 9540
rect 41782 9528 41788 9540
rect 41840 9528 41846 9580
rect 43070 9528 43076 9580
rect 43128 9568 43134 9580
rect 45005 9571 45063 9577
rect 45005 9568 45017 9571
rect 43128 9540 45017 9568
rect 43128 9528 43134 9540
rect 45005 9537 45017 9540
rect 45051 9537 45063 9571
rect 45005 9531 45063 9537
rect 46750 9528 46756 9580
rect 46808 9568 46814 9580
rect 46845 9571 46903 9577
rect 46845 9568 46857 9571
rect 46808 9540 46857 9568
rect 46808 9528 46814 9540
rect 46845 9537 46857 9540
rect 46891 9537 46903 9571
rect 47026 9568 47032 9580
rect 46987 9540 47032 9568
rect 46845 9531 46903 9537
rect 47026 9528 47032 9540
rect 47084 9528 47090 9580
rect 47670 9528 47676 9580
rect 47728 9568 47734 9580
rect 48225 9571 48283 9577
rect 48225 9568 48237 9571
rect 47728 9540 48237 9568
rect 47728 9528 47734 9540
rect 48225 9537 48237 9540
rect 48271 9537 48283 9571
rect 48225 9531 48283 9537
rect 48409 9571 48467 9577
rect 48409 9537 48421 9571
rect 48455 9568 48467 9571
rect 48590 9568 48596 9580
rect 48455 9540 48596 9568
rect 48455 9537 48467 9540
rect 48409 9531 48467 9537
rect 48590 9528 48596 9540
rect 48648 9528 48654 9580
rect 48866 9528 48872 9580
rect 48924 9568 48930 9580
rect 49145 9571 49203 9577
rect 49145 9568 49157 9571
rect 48924 9540 49157 9568
rect 48924 9528 48930 9540
rect 49145 9537 49157 9540
rect 49191 9537 49203 9571
rect 49145 9531 49203 9537
rect 49786 9528 49792 9580
rect 49844 9568 49850 9580
rect 50249 9571 50307 9577
rect 50249 9568 50261 9571
rect 49844 9540 50261 9568
rect 49844 9528 49850 9540
rect 50249 9537 50261 9540
rect 50295 9537 50307 9571
rect 50249 9531 50307 9537
rect 43162 9500 43168 9512
rect 40144 9472 40816 9500
rect 43123 9472 43168 9500
rect 30469 9435 30527 9441
rect 30469 9401 30481 9435
rect 30515 9432 30527 9435
rect 37550 9432 37556 9444
rect 30515 9404 31754 9432
rect 37511 9404 37556 9432
rect 30515 9401 30527 9404
rect 30469 9395 30527 9401
rect 30006 9364 30012 9376
rect 27764 9336 30012 9364
rect 27764 9324 27770 9336
rect 30006 9324 30012 9336
rect 30064 9324 30070 9376
rect 31726 9364 31754 9404
rect 37550 9392 37556 9404
rect 37608 9392 37614 9444
rect 33042 9364 33048 9376
rect 31726 9336 33048 9364
rect 33042 9324 33048 9336
rect 33100 9324 33106 9376
rect 33870 9324 33876 9376
rect 33928 9364 33934 9376
rect 34057 9367 34115 9373
rect 34057 9364 34069 9367
rect 33928 9336 34069 9364
rect 33928 9324 33934 9336
rect 34057 9333 34069 9336
rect 34103 9333 34115 9367
rect 37568 9364 37596 9392
rect 38562 9364 38568 9376
rect 37568 9336 38568 9364
rect 34057 9327 34115 9333
rect 38562 9324 38568 9336
rect 38620 9324 38626 9376
rect 38746 9324 38752 9376
rect 38804 9364 38810 9376
rect 40144 9364 40172 9472
rect 43162 9460 43168 9472
rect 43220 9460 43226 9512
rect 50356 9500 50384 9608
rect 50614 9596 50620 9608
rect 50672 9636 50678 9648
rect 50798 9636 50804 9648
rect 50672 9608 50804 9636
rect 50672 9596 50678 9608
rect 50798 9596 50804 9608
rect 50856 9596 50862 9648
rect 51442 9596 51448 9648
rect 51500 9636 51506 9648
rect 51500 9608 53788 9636
rect 51500 9596 51506 9608
rect 50516 9571 50574 9577
rect 50516 9537 50528 9571
rect 50562 9568 50574 9571
rect 52917 9571 52975 9577
rect 50562 9540 52868 9568
rect 50562 9537 50574 9540
rect 50516 9531 50574 9537
rect 44560 9472 50384 9500
rect 52840 9500 52868 9540
rect 52917 9537 52929 9571
rect 52963 9568 52975 9571
rect 53006 9568 53012 9580
rect 52963 9540 53012 9568
rect 52963 9537 52975 9540
rect 52917 9531 52975 9537
rect 53006 9528 53012 9540
rect 53064 9528 53070 9580
rect 53184 9571 53242 9577
rect 53184 9537 53196 9571
rect 53230 9568 53242 9571
rect 53466 9568 53472 9580
rect 53230 9540 53472 9568
rect 53230 9537 53242 9540
rect 53184 9531 53242 9537
rect 53466 9528 53472 9540
rect 53524 9528 53530 9580
rect 53760 9568 53788 9608
rect 53834 9596 53840 9648
rect 53892 9636 53898 9648
rect 54404 9636 54432 9676
rect 55953 9673 55965 9676
rect 55999 9673 56011 9707
rect 55953 9667 56011 9673
rect 56060 9676 56548 9704
rect 53892 9608 54432 9636
rect 53892 9596 53898 9608
rect 54478 9596 54484 9648
rect 54536 9636 54542 9648
rect 56060 9636 56088 9676
rect 54536 9608 56088 9636
rect 56520 9636 56548 9676
rect 56594 9664 56600 9716
rect 56652 9704 56658 9716
rect 56781 9707 56839 9713
rect 56781 9704 56793 9707
rect 56652 9676 56793 9704
rect 56652 9664 56658 9676
rect 56781 9673 56793 9676
rect 56827 9673 56839 9707
rect 56781 9667 56839 9673
rect 57054 9664 57060 9716
rect 57112 9704 57118 9716
rect 61194 9704 61200 9716
rect 57112 9676 61200 9704
rect 57112 9664 57118 9676
rect 61194 9664 61200 9676
rect 61252 9664 61258 9716
rect 63034 9664 63040 9716
rect 63092 9704 63098 9716
rect 64966 9704 64972 9716
rect 63092 9676 64972 9704
rect 63092 9664 63098 9676
rect 64966 9664 64972 9676
rect 65024 9664 65030 9716
rect 65242 9664 65248 9716
rect 65300 9704 65306 9716
rect 65521 9707 65579 9713
rect 65521 9704 65533 9707
rect 65300 9676 65533 9704
rect 65300 9664 65306 9676
rect 65521 9673 65533 9676
rect 65567 9673 65579 9707
rect 72602 9704 72608 9716
rect 65521 9667 65579 9673
rect 65628 9676 72608 9704
rect 56520 9608 56640 9636
rect 54536 9596 54542 9608
rect 54294 9568 54300 9580
rect 53760 9540 54300 9568
rect 54294 9528 54300 9540
rect 54352 9528 54358 9580
rect 55125 9571 55183 9577
rect 55125 9537 55137 9571
rect 55171 9568 55183 9571
rect 55490 9568 55496 9580
rect 55171 9540 55496 9568
rect 55171 9537 55183 9540
rect 55125 9531 55183 9537
rect 55490 9528 55496 9540
rect 55548 9528 55554 9580
rect 56137 9571 56195 9577
rect 56137 9537 56149 9571
rect 56183 9566 56195 9571
rect 56226 9566 56232 9580
rect 56183 9538 56232 9566
rect 56183 9537 56195 9538
rect 56137 9531 56195 9537
rect 56226 9528 56232 9538
rect 56284 9528 56290 9580
rect 56612 9577 56640 9608
rect 57146 9596 57152 9648
rect 57204 9636 57210 9648
rect 58066 9636 58072 9648
rect 57204 9608 58072 9636
rect 57204 9596 57210 9608
rect 58066 9596 58072 9608
rect 58124 9596 58130 9648
rect 58176 9608 62068 9636
rect 56597 9571 56655 9577
rect 56597 9537 56609 9571
rect 56643 9537 56655 9571
rect 57514 9568 57520 9580
rect 57475 9540 57520 9568
rect 56597 9531 56655 9537
rect 57514 9528 57520 9540
rect 57572 9528 57578 9580
rect 57698 9528 57704 9580
rect 57756 9568 57762 9580
rect 58176 9568 58204 9608
rect 57756 9540 58204 9568
rect 58253 9571 58311 9577
rect 57756 9528 57762 9540
rect 58253 9537 58265 9571
rect 58299 9537 58311 9571
rect 58253 9531 58311 9537
rect 56686 9500 56692 9512
rect 52840 9472 52960 9500
rect 41874 9392 41880 9444
rect 41932 9432 41938 9444
rect 42061 9435 42119 9441
rect 42061 9432 42073 9435
rect 41932 9404 42073 9432
rect 41932 9392 41938 9404
rect 42061 9401 42073 9404
rect 42107 9401 42119 9435
rect 42061 9395 42119 9401
rect 38804 9336 40172 9364
rect 38804 9324 38810 9336
rect 40218 9324 40224 9376
rect 40276 9364 40282 9376
rect 41966 9364 41972 9376
rect 40276 9336 41972 9364
rect 40276 9324 40282 9336
rect 41966 9324 41972 9336
rect 42024 9324 42030 9376
rect 42705 9367 42763 9373
rect 42705 9333 42717 9367
rect 42751 9364 42763 9367
rect 43070 9364 43076 9376
rect 42751 9336 43076 9364
rect 42751 9333 42763 9336
rect 42705 9327 42763 9333
rect 43070 9324 43076 9336
rect 43128 9364 43134 9376
rect 43898 9364 43904 9376
rect 43128 9336 43904 9364
rect 43128 9324 43134 9336
rect 43898 9324 43904 9336
rect 43956 9324 43962 9376
rect 44560 9373 44588 9472
rect 44726 9392 44732 9444
rect 44784 9432 44790 9444
rect 44784 9404 48820 9432
rect 44784 9392 44790 9404
rect 44545 9367 44603 9373
rect 44545 9333 44557 9367
rect 44591 9333 44603 9367
rect 45186 9364 45192 9376
rect 45147 9336 45192 9364
rect 44545 9327 44603 9333
rect 45186 9324 45192 9336
rect 45244 9324 45250 9376
rect 45738 9364 45744 9376
rect 45699 9336 45744 9364
rect 45738 9324 45744 9336
rect 45796 9324 45802 9376
rect 46290 9324 46296 9376
rect 46348 9364 46354 9376
rect 46348 9336 46393 9364
rect 46348 9324 46354 9336
rect 46750 9324 46756 9376
rect 46808 9364 46814 9376
rect 47302 9364 47308 9376
rect 46808 9336 47308 9364
rect 46808 9324 46814 9336
rect 47302 9324 47308 9336
rect 47360 9324 47366 9376
rect 48593 9367 48651 9373
rect 48593 9333 48605 9367
rect 48639 9364 48651 9367
rect 48682 9364 48688 9376
rect 48639 9336 48688 9364
rect 48639 9333 48651 9336
rect 48593 9327 48651 9333
rect 48682 9324 48688 9336
rect 48740 9324 48746 9376
rect 48792 9364 48820 9404
rect 49234 9392 49240 9444
rect 49292 9432 49298 9444
rect 49510 9432 49516 9444
rect 49292 9404 49516 9432
rect 49292 9392 49298 9404
rect 49510 9392 49516 9404
rect 49568 9392 49574 9444
rect 51629 9435 51687 9441
rect 51629 9401 51641 9435
rect 51675 9432 51687 9435
rect 52822 9432 52828 9444
rect 51675 9404 52828 9432
rect 51675 9401 51687 9404
rect 51629 9395 51687 9401
rect 52822 9392 52828 9404
rect 52880 9392 52886 9444
rect 51166 9364 51172 9376
rect 48792 9336 51172 9364
rect 51166 9324 51172 9336
rect 51224 9324 51230 9376
rect 52178 9324 52184 9376
rect 52236 9364 52242 9376
rect 52273 9367 52331 9373
rect 52273 9364 52285 9367
rect 52236 9336 52285 9364
rect 52236 9324 52242 9336
rect 52273 9333 52285 9336
rect 52319 9333 52331 9367
rect 52932 9364 52960 9472
rect 55324 9472 56692 9500
rect 55324 9441 55352 9472
rect 56686 9460 56692 9472
rect 56744 9460 56750 9512
rect 56870 9460 56876 9512
rect 56928 9500 56934 9512
rect 58268 9500 58296 9531
rect 59998 9528 60004 9580
rect 60056 9568 60062 9580
rect 60470 9571 60528 9577
rect 60470 9568 60482 9571
rect 60056 9540 60482 9568
rect 60056 9528 60062 9540
rect 60470 9537 60482 9540
rect 60516 9537 60528 9571
rect 60470 9531 60528 9537
rect 60734 9528 60740 9580
rect 60792 9568 60798 9580
rect 62040 9568 62068 9608
rect 62114 9596 62120 9648
rect 62172 9636 62178 9648
rect 62209 9639 62267 9645
rect 62209 9636 62221 9639
rect 62172 9608 62221 9636
rect 62172 9596 62178 9608
rect 62209 9605 62221 9608
rect 62255 9636 62267 9639
rect 65260 9636 65288 9664
rect 62255 9608 65288 9636
rect 62255 9605 62267 9608
rect 62209 9599 62267 9605
rect 63494 9568 63500 9580
rect 60792 9540 60837 9568
rect 62040 9540 63500 9568
rect 60792 9528 60798 9540
rect 63494 9528 63500 9540
rect 63552 9528 63558 9580
rect 63589 9571 63647 9577
rect 63589 9537 63601 9571
rect 63635 9568 63647 9571
rect 64693 9571 64751 9577
rect 64693 9568 64705 9571
rect 63635 9540 64705 9568
rect 63635 9537 63647 9540
rect 63589 9531 63647 9537
rect 64693 9537 64705 9540
rect 64739 9537 64751 9571
rect 64874 9568 64880 9580
rect 64835 9540 64880 9568
rect 64693 9531 64751 9537
rect 64874 9528 64880 9540
rect 64932 9528 64938 9580
rect 64966 9528 64972 9580
rect 65024 9568 65030 9580
rect 65024 9540 65069 9568
rect 65024 9528 65030 9540
rect 56928 9472 58296 9500
rect 56928 9460 56934 9472
rect 63678 9460 63684 9512
rect 63736 9500 63742 9512
rect 65628 9500 65656 9676
rect 72602 9664 72608 9676
rect 72660 9664 72666 9716
rect 73706 9664 73712 9716
rect 73764 9704 73770 9716
rect 82722 9704 82728 9716
rect 73764 9676 82728 9704
rect 73764 9664 73770 9676
rect 82722 9664 82728 9676
rect 82780 9664 82786 9716
rect 88334 9704 88340 9716
rect 85040 9676 85436 9704
rect 88295 9676 88340 9704
rect 66717 9639 66775 9645
rect 66717 9605 66729 9639
rect 66763 9636 66775 9639
rect 66898 9636 66904 9648
rect 66763 9608 66904 9636
rect 66763 9605 66775 9608
rect 66717 9599 66775 9605
rect 66898 9596 66904 9608
rect 66956 9596 66962 9648
rect 71774 9596 71780 9648
rect 71832 9636 71838 9648
rect 72881 9639 72939 9645
rect 72881 9636 72893 9639
rect 71832 9608 72893 9636
rect 71832 9596 71838 9608
rect 72881 9605 72893 9608
rect 72927 9605 72939 9639
rect 72881 9599 72939 9605
rect 67450 9528 67456 9580
rect 67508 9568 67514 9580
rect 67637 9571 67695 9577
rect 67637 9568 67649 9571
rect 67508 9540 67649 9568
rect 67508 9528 67514 9540
rect 67637 9537 67649 9540
rect 67683 9537 67695 9571
rect 67637 9531 67695 9537
rect 63736 9472 65656 9500
rect 72896 9500 72924 9599
rect 73430 9596 73436 9648
rect 73488 9636 73494 9648
rect 74718 9636 74724 9648
rect 73488 9608 73844 9636
rect 74679 9608 74724 9636
rect 73488 9596 73494 9608
rect 73706 9568 73712 9580
rect 73667 9540 73712 9568
rect 73706 9528 73712 9540
rect 73764 9528 73770 9580
rect 73816 9568 73844 9608
rect 74718 9596 74724 9608
rect 74776 9596 74782 9648
rect 75914 9596 75920 9648
rect 75972 9636 75978 9648
rect 75972 9608 76420 9636
rect 75972 9596 75978 9608
rect 76294 9571 76352 9577
rect 76294 9568 76306 9571
rect 73816 9540 76306 9568
rect 76294 9537 76306 9540
rect 76340 9537 76352 9571
rect 76392 9568 76420 9608
rect 76650 9596 76656 9648
rect 76708 9636 76714 9648
rect 77665 9639 77723 9645
rect 77665 9636 77677 9639
rect 76708 9608 77677 9636
rect 76708 9596 76714 9608
rect 77665 9605 77677 9608
rect 77711 9605 77723 9639
rect 77665 9599 77723 9605
rect 77021 9571 77079 9577
rect 77021 9568 77033 9571
rect 76392 9540 76512 9568
rect 76294 9531 76352 9537
rect 73893 9503 73951 9509
rect 73893 9500 73905 9503
rect 72896 9472 73905 9500
rect 63736 9460 63742 9472
rect 73893 9469 73905 9472
rect 73939 9469 73951 9503
rect 73893 9463 73951 9469
rect 74442 9460 74448 9512
rect 74500 9500 74506 9512
rect 76484 9500 76512 9540
rect 76668 9540 77033 9568
rect 76558 9500 76564 9512
rect 74500 9472 75592 9500
rect 76471 9472 76564 9500
rect 74500 9460 74506 9472
rect 55309 9435 55367 9441
rect 55309 9401 55321 9435
rect 55355 9401 55367 9435
rect 56594 9432 56600 9444
rect 55309 9395 55367 9401
rect 55508 9404 56600 9432
rect 54202 9364 54208 9376
rect 52932 9336 54208 9364
rect 52273 9327 52331 9333
rect 54202 9324 54208 9336
rect 54260 9324 54266 9376
rect 54297 9367 54355 9373
rect 54297 9333 54309 9367
rect 54343 9364 54355 9367
rect 55508 9364 55536 9404
rect 56594 9392 56600 9404
rect 56652 9392 56658 9444
rect 58434 9432 58440 9444
rect 58395 9404 58440 9432
rect 58434 9392 58440 9404
rect 58492 9392 58498 9444
rect 66254 9392 66260 9444
rect 66312 9432 66318 9444
rect 75181 9435 75239 9441
rect 75181 9432 75193 9435
rect 66312 9404 75193 9432
rect 66312 9392 66318 9404
rect 75181 9401 75193 9404
rect 75227 9401 75239 9435
rect 75181 9395 75239 9401
rect 54343 9336 55536 9364
rect 54343 9333 54355 9336
rect 54297 9327 54355 9333
rect 56410 9324 56416 9376
rect 56468 9364 56474 9376
rect 57333 9367 57391 9373
rect 57333 9364 57345 9367
rect 56468 9336 57345 9364
rect 56468 9324 56474 9336
rect 57333 9333 57345 9336
rect 57379 9333 57391 9367
rect 57333 9327 57391 9333
rect 58066 9324 58072 9376
rect 58124 9364 58130 9376
rect 59357 9367 59415 9373
rect 59357 9364 59369 9367
rect 58124 9336 59369 9364
rect 58124 9324 58130 9336
rect 59357 9333 59369 9336
rect 59403 9333 59415 9367
rect 61654 9364 61660 9376
rect 61615 9336 61660 9364
rect 59357 9327 59415 9333
rect 61654 9324 61660 9336
rect 61712 9324 61718 9376
rect 63770 9364 63776 9376
rect 63731 9336 63776 9364
rect 63770 9324 63776 9336
rect 63828 9324 63834 9376
rect 65794 9324 65800 9376
rect 65852 9364 65858 9376
rect 66073 9367 66131 9373
rect 66073 9364 66085 9367
rect 65852 9336 66085 9364
rect 65852 9324 65858 9336
rect 66073 9333 66085 9336
rect 66119 9333 66131 9367
rect 66073 9327 66131 9333
rect 66714 9324 66720 9376
rect 66772 9364 66778 9376
rect 67453 9367 67511 9373
rect 67453 9364 67465 9367
rect 66772 9336 67465 9364
rect 66772 9324 66778 9336
rect 67453 9333 67465 9336
rect 67499 9333 67511 9367
rect 73522 9364 73528 9376
rect 73483 9336 73528 9364
rect 67453 9327 67511 9333
rect 73522 9324 73528 9336
rect 73580 9324 73586 9376
rect 75564 9364 75592 9472
rect 76558 9460 76564 9472
rect 76616 9460 76622 9512
rect 76668 9364 76696 9540
rect 77021 9537 77033 9540
rect 77067 9537 77079 9571
rect 77021 9531 77079 9537
rect 77680 9500 77708 9599
rect 79870 9596 79876 9648
rect 79928 9636 79934 9648
rect 84838 9636 84844 9648
rect 79928 9608 84844 9636
rect 79928 9596 79934 9608
rect 84838 9596 84844 9608
rect 84896 9596 84902 9648
rect 84942 9639 85000 9645
rect 84942 9605 84954 9639
rect 84988 9636 85000 9639
rect 85040 9636 85068 9676
rect 84988 9608 85068 9636
rect 84988 9605 85000 9608
rect 84942 9599 85000 9605
rect 85114 9596 85120 9648
rect 85172 9636 85178 9648
rect 85408 9636 85436 9676
rect 88334 9664 88340 9676
rect 88392 9664 88398 9716
rect 89070 9664 89076 9716
rect 89128 9704 89134 9716
rect 95418 9704 95424 9716
rect 89128 9676 89576 9704
rect 89128 9664 89134 9676
rect 85761 9639 85819 9645
rect 85761 9636 85773 9639
rect 85172 9608 85344 9636
rect 85408 9608 85773 9636
rect 85172 9596 85178 9608
rect 79686 9528 79692 9580
rect 79744 9568 79750 9580
rect 83185 9571 83243 9577
rect 83185 9568 83197 9571
rect 79744 9540 83197 9568
rect 79744 9528 79750 9540
rect 83185 9537 83197 9540
rect 83231 9568 83243 9571
rect 85209 9571 85267 9577
rect 85209 9568 85221 9571
rect 83231 9540 85221 9568
rect 83231 9537 83243 9540
rect 83185 9531 83243 9537
rect 85209 9537 85221 9540
rect 85255 9537 85267 9571
rect 85209 9531 85267 9537
rect 82538 9500 82544 9512
rect 77680 9472 82544 9500
rect 82538 9460 82544 9472
rect 82596 9460 82602 9512
rect 82998 9460 83004 9512
rect 83056 9500 83062 9512
rect 85316 9500 85344 9608
rect 85761 9605 85773 9608
rect 85807 9636 85819 9639
rect 89548 9636 89576 9676
rect 89732 9676 92152 9704
rect 89732 9636 89760 9676
rect 85807 9608 89484 9636
rect 89548 9608 89760 9636
rect 85807 9605 85819 9608
rect 85761 9599 85819 9605
rect 85390 9528 85396 9580
rect 85448 9568 85454 9580
rect 88242 9568 88248 9580
rect 85448 9540 88248 9568
rect 85448 9528 85454 9540
rect 88242 9528 88248 9540
rect 88300 9528 88306 9580
rect 88334 9528 88340 9580
rect 88392 9568 88398 9580
rect 89073 9571 89131 9577
rect 89073 9568 89085 9571
rect 88392 9540 89085 9568
rect 88392 9528 88398 9540
rect 89073 9537 89085 9540
rect 89119 9537 89131 9571
rect 89329 9571 89387 9577
rect 89329 9568 89341 9571
rect 89073 9531 89131 9537
rect 89180 9540 89341 9568
rect 89180 9500 89208 9540
rect 89329 9537 89341 9540
rect 89375 9537 89387 9571
rect 89456 9568 89484 9608
rect 90450 9596 90456 9648
rect 90508 9636 90514 9648
rect 92026 9639 92084 9645
rect 92026 9636 92038 9639
rect 90508 9608 92038 9636
rect 90508 9596 90514 9608
rect 92026 9605 92038 9608
rect 92072 9605 92084 9639
rect 92124 9636 92152 9676
rect 93504 9676 93992 9704
rect 93504 9636 93532 9676
rect 92124 9608 93532 9636
rect 93581 9639 93639 9645
rect 92026 9599 92084 9605
rect 93581 9605 93593 9639
rect 93627 9636 93639 9639
rect 93854 9636 93860 9648
rect 93627 9608 93860 9636
rect 93627 9605 93639 9608
rect 93581 9599 93639 9605
rect 93854 9596 93860 9608
rect 93912 9596 93918 9648
rect 93964 9636 93992 9676
rect 94792 9676 95424 9704
rect 94792 9636 94820 9676
rect 95418 9664 95424 9676
rect 95476 9664 95482 9716
rect 96341 9707 96399 9713
rect 96341 9704 96353 9707
rect 95620 9676 96353 9704
rect 93964 9608 94820 9636
rect 95522 9639 95580 9645
rect 95522 9605 95534 9639
rect 95568 9636 95580 9639
rect 95620 9636 95648 9676
rect 96341 9673 96353 9676
rect 96387 9704 96399 9707
rect 98086 9704 98092 9716
rect 96387 9676 98092 9704
rect 96387 9673 96399 9676
rect 96341 9667 96399 9673
rect 98086 9664 98092 9676
rect 98144 9664 98150 9716
rect 98564 9676 98868 9704
rect 95568 9608 95648 9636
rect 95568 9605 95580 9608
rect 95522 9599 95580 9605
rect 95694 9596 95700 9648
rect 95752 9636 95758 9648
rect 98564 9636 98592 9676
rect 98730 9636 98736 9648
rect 95752 9608 95832 9636
rect 95752 9596 95758 9608
rect 95804 9577 95832 9608
rect 95896 9608 98592 9636
rect 98691 9608 98736 9636
rect 95789 9571 95847 9577
rect 89456 9540 95731 9568
rect 89329 9531 89387 9537
rect 83056 9472 84240 9500
rect 85316 9472 89208 9500
rect 83056 9460 83062 9472
rect 77205 9435 77263 9441
rect 77205 9401 77217 9435
rect 77251 9432 77263 9435
rect 77294 9432 77300 9444
rect 77251 9404 77300 9432
rect 77251 9401 77263 9404
rect 77205 9395 77263 9401
rect 77294 9392 77300 9404
rect 77352 9392 77358 9444
rect 78674 9392 78680 9444
rect 78732 9432 78738 9444
rect 79962 9432 79968 9444
rect 78732 9404 79968 9432
rect 78732 9392 78738 9404
rect 79962 9392 79968 9404
rect 80020 9392 80026 9444
rect 82262 9392 82268 9444
rect 82320 9432 82326 9444
rect 83829 9435 83887 9441
rect 83829 9432 83841 9435
rect 82320 9404 83841 9432
rect 82320 9392 82326 9404
rect 83829 9401 83841 9404
rect 83875 9401 83887 9435
rect 84212 9432 84240 9472
rect 90082 9460 90088 9512
rect 90140 9500 90146 9512
rect 92290 9500 92296 9512
rect 90140 9472 91048 9500
rect 92251 9472 92296 9500
rect 90140 9460 90146 9472
rect 84212 9404 84332 9432
rect 83829 9395 83887 9401
rect 84304 9376 84332 9404
rect 85206 9392 85212 9444
rect 85264 9432 85270 9444
rect 89070 9432 89076 9444
rect 85264 9404 89076 9432
rect 85264 9392 85270 9404
rect 89070 9392 89076 9404
rect 89128 9392 89134 9444
rect 90913 9435 90971 9441
rect 90913 9432 90925 9435
rect 90284 9404 90925 9432
rect 75564 9336 76696 9364
rect 79594 9324 79600 9376
rect 79652 9364 79658 9376
rect 79873 9367 79931 9373
rect 79873 9364 79885 9367
rect 79652 9336 79885 9364
rect 79652 9324 79658 9336
rect 79873 9333 79885 9336
rect 79919 9364 79931 9367
rect 81434 9364 81440 9376
rect 79919 9336 81440 9364
rect 79919 9333 79931 9336
rect 79873 9327 79931 9333
rect 81434 9324 81440 9336
rect 81492 9324 81498 9376
rect 82630 9324 82636 9376
rect 82688 9364 82694 9376
rect 84194 9364 84200 9376
rect 82688 9336 84200 9364
rect 82688 9324 82694 9336
rect 84194 9324 84200 9336
rect 84252 9324 84258 9376
rect 84286 9324 84292 9376
rect 84344 9324 84350 9376
rect 84470 9324 84476 9376
rect 84528 9364 84534 9376
rect 90284 9364 90312 9404
rect 90913 9401 90925 9404
rect 90959 9401 90971 9435
rect 90913 9395 90971 9401
rect 90450 9364 90456 9376
rect 84528 9336 90312 9364
rect 90411 9336 90456 9364
rect 84528 9324 84534 9336
rect 90450 9324 90456 9336
rect 90508 9324 90514 9376
rect 91020 9364 91048 9472
rect 92290 9460 92296 9472
rect 92348 9500 92354 9512
rect 92934 9500 92940 9512
rect 92348 9472 92940 9500
rect 92348 9460 92354 9472
rect 92934 9460 92940 9472
rect 92992 9460 92998 9512
rect 95703 9500 95731 9540
rect 95789 9537 95801 9571
rect 95835 9537 95847 9571
rect 95789 9531 95847 9537
rect 95896 9500 95924 9608
rect 98730 9596 98736 9608
rect 98788 9596 98794 9648
rect 98840 9636 98868 9676
rect 98914 9664 98920 9716
rect 98972 9704 98978 9716
rect 113542 9704 113548 9716
rect 98972 9676 113548 9704
rect 98972 9664 98978 9676
rect 113542 9664 113548 9676
rect 113600 9664 113606 9716
rect 113726 9664 113732 9716
rect 113784 9704 113790 9716
rect 113784 9676 117268 9704
rect 113784 9664 113790 9676
rect 108022 9636 108028 9648
rect 98840 9608 108028 9636
rect 108022 9596 108028 9608
rect 108080 9596 108086 9648
rect 108500 9608 113588 9636
rect 98549 9571 98607 9577
rect 98549 9568 98561 9571
rect 95703 9472 95924 9500
rect 97276 9540 98561 9568
rect 92842 9364 92848 9376
rect 91020 9336 92848 9364
rect 92842 9324 92848 9336
rect 92900 9324 92906 9376
rect 93854 9324 93860 9376
rect 93912 9364 93918 9376
rect 94409 9367 94467 9373
rect 94409 9364 94421 9367
rect 93912 9336 94421 9364
rect 93912 9324 93918 9336
rect 94409 9333 94421 9336
rect 94455 9333 94467 9367
rect 94409 9327 94467 9333
rect 94498 9324 94504 9376
rect 94556 9364 94562 9376
rect 97276 9364 97304 9540
rect 98549 9537 98561 9540
rect 98595 9537 98607 9571
rect 99374 9568 99380 9580
rect 98549 9531 98607 9537
rect 98840 9540 99380 9568
rect 98365 9503 98423 9509
rect 98365 9469 98377 9503
rect 98411 9500 98423 9503
rect 98840 9500 98868 9540
rect 99374 9528 99380 9540
rect 99432 9528 99438 9580
rect 99552 9571 99610 9577
rect 99552 9537 99564 9571
rect 99598 9568 99610 9571
rect 104250 9568 104256 9580
rect 99598 9540 104256 9568
rect 99598 9537 99610 9540
rect 99552 9531 99610 9537
rect 104250 9528 104256 9540
rect 104308 9528 104314 9580
rect 104434 9568 104440 9580
rect 104395 9540 104440 9568
rect 104434 9528 104440 9540
rect 104492 9528 104498 9580
rect 104618 9568 104624 9580
rect 104579 9540 104624 9568
rect 104618 9528 104624 9540
rect 104676 9528 104682 9580
rect 105630 9568 105636 9580
rect 105591 9540 105636 9568
rect 105630 9528 105636 9540
rect 105688 9528 105694 9580
rect 105814 9528 105820 9580
rect 105872 9568 105878 9580
rect 107838 9568 107844 9580
rect 105872 9540 107844 9568
rect 105872 9528 105878 9540
rect 107838 9528 107844 9540
rect 107896 9528 107902 9580
rect 108393 9572 108451 9577
rect 108500 9572 108528 9608
rect 108393 9571 108528 9572
rect 108393 9537 108405 9571
rect 108439 9544 108528 9571
rect 108439 9537 108451 9544
rect 108393 9531 108451 9537
rect 110782 9528 110788 9580
rect 110840 9568 110846 9580
rect 111521 9571 111579 9577
rect 111521 9568 111533 9571
rect 110840 9540 111533 9568
rect 110840 9528 110846 9540
rect 111521 9537 111533 9540
rect 111567 9537 111579 9571
rect 113453 9571 113511 9577
rect 113453 9568 113465 9571
rect 111521 9531 111579 9537
rect 112732 9540 113465 9568
rect 98411 9472 98868 9500
rect 99285 9503 99343 9509
rect 98411 9469 98423 9472
rect 98365 9463 98423 9469
rect 99285 9469 99297 9503
rect 99331 9469 99343 9503
rect 99285 9463 99343 9469
rect 97350 9392 97356 9444
rect 97408 9432 97414 9444
rect 99300 9432 99328 9463
rect 107654 9460 107660 9512
rect 107712 9500 107718 9512
rect 112732 9509 112760 9540
rect 113453 9537 113465 9540
rect 113499 9537 113511 9571
rect 113560 9568 113588 9608
rect 113818 9596 113824 9648
rect 113876 9636 113882 9648
rect 116302 9636 116308 9648
rect 113876 9608 116308 9636
rect 113876 9596 113882 9608
rect 116302 9596 116308 9608
rect 116360 9596 116366 9648
rect 116578 9596 116584 9648
rect 116636 9645 116642 9648
rect 116636 9636 116648 9645
rect 117240 9636 117268 9676
rect 117314 9664 117320 9716
rect 117372 9704 117378 9716
rect 117409 9707 117467 9713
rect 117409 9704 117421 9707
rect 117372 9676 117421 9704
rect 117372 9664 117378 9676
rect 117409 9673 117421 9676
rect 117455 9673 117467 9707
rect 117409 9667 117467 9673
rect 117424 9636 117452 9667
rect 120994 9664 121000 9716
rect 121052 9704 121058 9716
rect 132589 9707 132647 9713
rect 121052 9676 132540 9704
rect 121052 9664 121058 9676
rect 130286 9636 130292 9648
rect 116636 9608 116681 9636
rect 117240 9608 117360 9636
rect 117424 9608 130292 9636
rect 116636 9599 116648 9608
rect 116636 9596 116642 9599
rect 117332 9568 117360 9608
rect 117958 9568 117964 9580
rect 113560 9540 117268 9568
rect 117332 9540 117964 9568
rect 113453 9531 113511 9537
rect 112717 9503 112775 9509
rect 112717 9500 112729 9503
rect 107712 9472 112729 9500
rect 107712 9460 107718 9472
rect 112717 9469 112729 9472
rect 112763 9469 112775 9503
rect 113266 9500 113272 9512
rect 113227 9472 113272 9500
rect 112717 9463 112775 9469
rect 113266 9460 113272 9472
rect 113324 9460 113330 9512
rect 113818 9500 113824 9512
rect 113376 9472 113824 9500
rect 101214 9432 101220 9444
rect 97408 9404 99328 9432
rect 97408 9392 97414 9404
rect 97813 9367 97871 9373
rect 97813 9364 97825 9367
rect 94556 9336 97825 9364
rect 94556 9324 94562 9336
rect 97813 9333 97825 9336
rect 97859 9333 97871 9367
rect 99300 9364 99328 9404
rect 100588 9404 101220 9432
rect 100588 9364 100616 9404
rect 101214 9392 101220 9404
rect 101272 9432 101278 9444
rect 108390 9432 108396 9444
rect 101272 9404 108396 9432
rect 101272 9392 101278 9404
rect 108390 9392 108396 9404
rect 108448 9392 108454 9444
rect 108577 9435 108635 9441
rect 108577 9401 108589 9435
rect 108623 9432 108635 9435
rect 108666 9432 108672 9444
rect 108623 9404 108672 9432
rect 108623 9401 108635 9404
rect 108577 9395 108635 9401
rect 108666 9392 108672 9404
rect 108724 9392 108730 9444
rect 113376 9432 113404 9472
rect 113818 9460 113824 9472
rect 113876 9460 113882 9512
rect 114738 9500 114744 9512
rect 114699 9472 114744 9500
rect 114738 9460 114744 9472
rect 114796 9460 114802 9512
rect 115382 9460 115388 9512
rect 115440 9500 115446 9512
rect 115842 9500 115848 9512
rect 115440 9472 115848 9500
rect 115440 9460 115446 9472
rect 115842 9460 115848 9472
rect 115900 9460 115906 9512
rect 116857 9503 116915 9509
rect 116857 9469 116869 9503
rect 116903 9500 116915 9503
rect 117130 9500 117136 9512
rect 116903 9472 117136 9500
rect 116903 9469 116915 9472
rect 116857 9463 116915 9469
rect 117130 9460 117136 9472
rect 117188 9460 117194 9512
rect 108776 9404 113404 9432
rect 113637 9435 113695 9441
rect 99300 9336 100616 9364
rect 100665 9367 100723 9373
rect 97813 9327 97871 9333
rect 100665 9333 100677 9367
rect 100711 9364 100723 9367
rect 103238 9364 103244 9376
rect 100711 9336 103244 9364
rect 100711 9333 100723 9336
rect 100665 9327 100723 9333
rect 103238 9324 103244 9336
rect 103296 9324 103302 9376
rect 103422 9364 103428 9376
rect 103383 9336 103428 9364
rect 103422 9324 103428 9336
rect 103480 9324 103486 9376
rect 104805 9367 104863 9373
rect 104805 9333 104817 9367
rect 104851 9364 104863 9367
rect 105354 9364 105360 9376
rect 104851 9336 105360 9364
rect 104851 9333 104863 9336
rect 104805 9327 104863 9333
rect 105354 9324 105360 9336
rect 105412 9324 105418 9376
rect 105446 9324 105452 9376
rect 105504 9364 105510 9376
rect 107194 9364 107200 9376
rect 105504 9336 105549 9364
rect 107155 9336 107200 9364
rect 105504 9324 105510 9336
rect 107194 9324 107200 9336
rect 107252 9324 107258 9376
rect 107286 9324 107292 9376
rect 107344 9364 107350 9376
rect 108776 9364 108804 9404
rect 113637 9401 113649 9435
rect 113683 9432 113695 9435
rect 117240 9432 117268 9540
rect 117958 9528 117964 9540
rect 118016 9528 118022 9580
rect 120997 9571 121055 9577
rect 120997 9537 121009 9571
rect 121043 9568 121055 9571
rect 121086 9568 121092 9580
rect 121043 9540 121092 9568
rect 121043 9537 121055 9540
rect 120997 9531 121055 9537
rect 121086 9528 121092 9540
rect 121144 9528 121150 9580
rect 121825 9571 121883 9577
rect 121825 9537 121837 9571
rect 121871 9568 121883 9571
rect 121914 9568 121920 9580
rect 121871 9540 121920 9568
rect 121871 9537 121883 9540
rect 121825 9531 121883 9537
rect 121914 9528 121920 9540
rect 121972 9528 121978 9580
rect 122092 9571 122150 9577
rect 122092 9537 122104 9571
rect 122138 9568 122150 9571
rect 123665 9571 123723 9577
rect 123665 9568 123677 9571
rect 122138 9540 123677 9568
rect 122138 9537 122150 9540
rect 122092 9531 122150 9537
rect 123665 9537 123677 9540
rect 123711 9537 123723 9571
rect 124398 9568 124404 9580
rect 124359 9540 124404 9568
rect 123665 9531 123723 9537
rect 118329 9503 118387 9509
rect 118329 9469 118341 9503
rect 118375 9500 118387 9503
rect 121730 9500 121736 9512
rect 118375 9472 121736 9500
rect 118375 9469 118387 9472
rect 118329 9463 118387 9469
rect 121730 9460 121736 9472
rect 121788 9460 121794 9512
rect 123680 9500 123708 9531
rect 124398 9528 124404 9540
rect 124456 9528 124462 9580
rect 125505 9571 125563 9577
rect 125505 9537 125517 9571
rect 125551 9568 125563 9571
rect 127894 9568 127900 9580
rect 125551 9540 127900 9568
rect 125551 9537 125563 9540
rect 125505 9531 125563 9537
rect 127894 9528 127900 9540
rect 127952 9528 127958 9580
rect 129660 9577 129688 9608
rect 130286 9596 130292 9608
rect 130344 9596 130350 9648
rect 130930 9596 130936 9648
rect 130988 9636 130994 9648
rect 132512 9636 132540 9676
rect 132589 9673 132601 9707
rect 132635 9704 132647 9707
rect 133782 9704 133788 9716
rect 132635 9676 133788 9704
rect 132635 9673 132647 9676
rect 132589 9667 132647 9673
rect 133782 9664 133788 9676
rect 133840 9664 133846 9716
rect 133892 9676 136864 9704
rect 133892 9636 133920 9676
rect 136836 9645 136864 9676
rect 136910 9664 136916 9716
rect 136968 9704 136974 9716
rect 143534 9704 143540 9716
rect 136968 9676 138888 9704
rect 136968 9664 136974 9676
rect 130988 9608 132264 9636
rect 132512 9608 133920 9636
rect 136821 9639 136879 9645
rect 130988 9596 130994 9608
rect 131224 9577 131252 9608
rect 129389 9571 129447 9577
rect 129389 9537 129401 9571
rect 129435 9568 129447 9571
rect 129645 9571 129703 9577
rect 129435 9540 129596 9568
rect 129435 9537 129447 9540
rect 129389 9531 129447 9537
rect 125686 9500 125692 9512
rect 123680 9472 125456 9500
rect 125647 9472 125692 9500
rect 123205 9435 123263 9441
rect 113683 9404 115612 9432
rect 117240 9404 121868 9432
rect 113683 9401 113695 9404
rect 113637 9395 113695 9401
rect 110046 9364 110052 9376
rect 107344 9336 108804 9364
rect 110007 9336 110052 9364
rect 107344 9324 107350 9336
rect 110046 9324 110052 9336
rect 110104 9324 110110 9376
rect 110782 9324 110788 9376
rect 110840 9364 110846 9376
rect 110966 9364 110972 9376
rect 110840 9336 110972 9364
rect 110840 9324 110846 9336
rect 110966 9324 110972 9336
rect 111024 9324 111030 9376
rect 111242 9324 111248 9376
rect 111300 9364 111306 9376
rect 111337 9367 111395 9373
rect 111337 9364 111349 9367
rect 111300 9336 111349 9364
rect 111300 9324 111306 9336
rect 111337 9333 111349 9336
rect 111383 9333 111395 9367
rect 111337 9327 111395 9333
rect 114002 9324 114008 9376
rect 114060 9364 114066 9376
rect 114097 9367 114155 9373
rect 114097 9364 114109 9367
rect 114060 9336 114109 9364
rect 114060 9324 114066 9336
rect 114097 9333 114109 9336
rect 114143 9364 114155 9367
rect 114186 9364 114192 9376
rect 114143 9336 114192 9364
rect 114143 9333 114155 9336
rect 114097 9327 114155 9333
rect 114186 9324 114192 9336
rect 114244 9324 114250 9376
rect 115382 9324 115388 9376
rect 115440 9364 115446 9376
rect 115477 9367 115535 9373
rect 115477 9364 115489 9367
rect 115440 9336 115489 9364
rect 115440 9324 115446 9336
rect 115477 9333 115489 9336
rect 115523 9333 115535 9367
rect 115584 9364 115612 9404
rect 117498 9364 117504 9376
rect 115584 9336 117504 9364
rect 115477 9327 115535 9333
rect 117498 9324 117504 9336
rect 117556 9324 117562 9376
rect 118326 9324 118332 9376
rect 118384 9364 118390 9376
rect 118789 9367 118847 9373
rect 118789 9364 118801 9367
rect 118384 9336 118801 9364
rect 118384 9324 118390 9336
rect 118789 9333 118801 9336
rect 118835 9333 118847 9367
rect 118789 9327 118847 9333
rect 119798 9324 119804 9376
rect 119856 9364 119862 9376
rect 119893 9367 119951 9373
rect 119893 9364 119905 9367
rect 119856 9336 119905 9364
rect 119856 9324 119862 9336
rect 119893 9333 119905 9336
rect 119939 9333 119951 9367
rect 119893 9327 119951 9333
rect 119982 9324 119988 9376
rect 120040 9364 120046 9376
rect 121362 9364 121368 9376
rect 120040 9336 121368 9364
rect 120040 9324 120046 9336
rect 121362 9324 121368 9336
rect 121420 9324 121426 9376
rect 121840 9364 121868 9404
rect 123205 9401 123217 9435
rect 123251 9432 123263 9435
rect 123294 9432 123300 9444
rect 123251 9404 123300 9432
rect 123251 9401 123263 9404
rect 123205 9395 123263 9401
rect 123294 9392 123300 9404
rect 123352 9392 123358 9444
rect 125321 9435 125379 9441
rect 125321 9432 125333 9435
rect 123404 9404 125333 9432
rect 123404 9364 123432 9404
rect 125321 9401 125333 9404
rect 125367 9401 125379 9435
rect 125428 9432 125456 9472
rect 125686 9460 125692 9472
rect 125744 9460 125750 9512
rect 125962 9460 125968 9512
rect 126020 9500 126026 9512
rect 127526 9500 127532 9512
rect 126020 9472 127532 9500
rect 126020 9460 126026 9472
rect 127526 9460 127532 9472
rect 127584 9460 127590 9512
rect 129568 9500 129596 9540
rect 129645 9537 129657 9571
rect 129691 9537 129703 9571
rect 129645 9531 129703 9537
rect 131209 9571 131267 9577
rect 131209 9537 131221 9571
rect 131255 9537 131267 9571
rect 131465 9571 131523 9577
rect 131465 9568 131477 9571
rect 131209 9531 131267 9537
rect 131316 9540 131477 9568
rect 130194 9500 130200 9512
rect 129568 9472 130200 9500
rect 130194 9460 130200 9472
rect 130252 9460 130258 9512
rect 130286 9460 130292 9512
rect 130344 9500 130350 9512
rect 131316 9500 131344 9540
rect 131465 9537 131477 9540
rect 131511 9537 131523 9571
rect 131465 9531 131523 9537
rect 130344 9472 131344 9500
rect 132236 9500 132264 9608
rect 136821 9605 136833 9639
rect 136867 9636 136879 9639
rect 137554 9636 137560 9648
rect 136867 9608 137560 9636
rect 136867 9605 136879 9608
rect 136821 9599 136879 9605
rect 137554 9596 137560 9608
rect 137612 9596 137618 9648
rect 138860 9636 138888 9676
rect 143368 9676 143540 9704
rect 139486 9636 139492 9648
rect 137664 9608 138327 9636
rect 138860 9608 139492 9636
rect 132586 9528 132592 9580
rect 132644 9568 132650 9580
rect 133506 9568 133512 9580
rect 132644 9540 133512 9568
rect 132644 9528 132650 9540
rect 133506 9528 133512 9540
rect 133564 9568 133570 9580
rect 133673 9571 133731 9577
rect 133673 9568 133685 9571
rect 133564 9540 133685 9568
rect 133564 9528 133570 9540
rect 133673 9537 133685 9540
rect 133719 9537 133731 9571
rect 133673 9531 133731 9537
rect 134058 9528 134064 9580
rect 134116 9568 134122 9580
rect 134978 9568 134984 9580
rect 134116 9540 134984 9568
rect 134116 9528 134122 9540
rect 134978 9528 134984 9540
rect 135036 9568 135042 9580
rect 137462 9568 137468 9580
rect 135036 9540 137468 9568
rect 135036 9528 135042 9540
rect 137462 9528 137468 9540
rect 137520 9528 137526 9580
rect 133138 9500 133144 9512
rect 132236 9472 133144 9500
rect 130344 9460 130350 9472
rect 133138 9460 133144 9472
rect 133196 9500 133202 9512
rect 133417 9503 133475 9509
rect 133417 9500 133429 9503
rect 133196 9472 133429 9500
rect 133196 9460 133202 9472
rect 133417 9469 133429 9472
rect 133463 9469 133475 9503
rect 137664 9500 137692 9608
rect 138181 9571 138239 9577
rect 138181 9568 138193 9571
rect 133417 9463 133475 9469
rect 134444 9472 137692 9500
rect 137756 9540 138193 9568
rect 127713 9435 127771 9441
rect 127713 9432 127725 9435
rect 125428 9404 127725 9432
rect 125321 9395 125379 9401
rect 127713 9401 127725 9404
rect 127759 9432 127771 9435
rect 127759 9404 128768 9432
rect 127759 9401 127771 9404
rect 127713 9395 127771 9401
rect 121840 9336 123432 9364
rect 123846 9324 123852 9376
rect 123904 9364 123910 9376
rect 125594 9364 125600 9376
rect 123904 9336 125600 9364
rect 123904 9324 123910 9336
rect 125594 9324 125600 9336
rect 125652 9364 125658 9376
rect 126146 9364 126152 9376
rect 125652 9336 126152 9364
rect 125652 9324 125658 9336
rect 126146 9324 126152 9336
rect 126204 9324 126210 9376
rect 126238 9324 126244 9376
rect 126296 9364 126302 9376
rect 126701 9367 126759 9373
rect 126701 9364 126713 9367
rect 126296 9336 126713 9364
rect 126296 9324 126302 9336
rect 126701 9333 126713 9336
rect 126747 9333 126759 9367
rect 126701 9327 126759 9333
rect 127066 9324 127072 9376
rect 127124 9364 127130 9376
rect 128262 9364 128268 9376
rect 127124 9336 128268 9364
rect 127124 9324 127130 9336
rect 128262 9324 128268 9336
rect 128320 9324 128326 9376
rect 128740 9364 128768 9404
rect 129642 9392 129648 9444
rect 129700 9432 129706 9444
rect 131114 9432 131120 9444
rect 129700 9404 131120 9432
rect 129700 9392 129706 9404
rect 131114 9392 131120 9404
rect 131172 9392 131178 9444
rect 132218 9392 132224 9444
rect 132276 9432 132282 9444
rect 132276 9404 132632 9432
rect 132276 9392 132282 9404
rect 132494 9364 132500 9376
rect 128740 9336 132500 9364
rect 132494 9324 132500 9336
rect 132552 9324 132558 9376
rect 132604 9364 132632 9404
rect 134444 9364 134472 9472
rect 135530 9392 135536 9444
rect 135588 9432 135594 9444
rect 135717 9435 135775 9441
rect 135717 9432 135729 9435
rect 135588 9404 135729 9432
rect 135588 9392 135594 9404
rect 135717 9401 135729 9404
rect 135763 9432 135775 9435
rect 136361 9435 136419 9441
rect 136361 9432 136373 9435
rect 135763 9404 136373 9432
rect 135763 9401 135775 9404
rect 135717 9395 135775 9401
rect 136361 9401 136373 9404
rect 136407 9432 136419 9435
rect 136910 9432 136916 9444
rect 136407 9404 136916 9432
rect 136407 9401 136419 9404
rect 136361 9395 136419 9401
rect 136910 9392 136916 9404
rect 136968 9392 136974 9444
rect 134794 9364 134800 9376
rect 132604 9336 134472 9364
rect 134755 9336 134800 9364
rect 134794 9324 134800 9336
rect 134852 9324 134858 9376
rect 137370 9364 137376 9376
rect 137331 9336 137376 9364
rect 137370 9324 137376 9336
rect 137428 9364 137434 9376
rect 137756 9364 137784 9540
rect 138181 9537 138193 9540
rect 138227 9537 138239 9571
rect 138299 9568 138327 9608
rect 139486 9596 139492 9608
rect 139544 9596 139550 9648
rect 140590 9596 140596 9648
rect 140648 9636 140654 9648
rect 143368 9636 143396 9676
rect 143534 9664 143540 9676
rect 143592 9664 143598 9716
rect 143902 9664 143908 9716
rect 143960 9704 143966 9716
rect 147398 9704 147404 9716
rect 143960 9676 147404 9704
rect 143960 9664 143966 9676
rect 147398 9664 147404 9676
rect 147456 9664 147462 9716
rect 147950 9664 147956 9716
rect 148008 9704 148014 9716
rect 149514 9704 149520 9716
rect 148008 9676 149520 9704
rect 148008 9664 148014 9676
rect 149514 9664 149520 9676
rect 149572 9664 149578 9716
rect 149793 9707 149851 9713
rect 149793 9673 149805 9707
rect 149839 9704 149851 9707
rect 150986 9704 150992 9716
rect 149839 9676 150992 9704
rect 149839 9673 149851 9676
rect 149793 9667 149851 9673
rect 150986 9664 150992 9676
rect 151044 9664 151050 9716
rect 151262 9704 151268 9716
rect 151223 9676 151268 9704
rect 151262 9664 151268 9676
rect 151320 9664 151326 9716
rect 151722 9664 151728 9716
rect 151780 9704 151786 9716
rect 158070 9704 158076 9716
rect 151780 9676 158076 9704
rect 151780 9664 151786 9676
rect 158070 9664 158076 9676
rect 158128 9664 158134 9716
rect 158254 9704 158260 9716
rect 158215 9676 158260 9704
rect 158254 9664 158260 9676
rect 158312 9664 158318 9716
rect 140648 9608 143396 9636
rect 143460 9608 145144 9636
rect 140648 9596 140654 9608
rect 140038 9568 140044 9580
rect 138299 9540 140044 9568
rect 138181 9531 138239 9537
rect 140038 9528 140044 9540
rect 140096 9528 140102 9580
rect 141160 9577 141188 9608
rect 143460 9580 143488 9608
rect 140961 9571 141019 9577
rect 140961 9537 140973 9571
rect 141007 9537 141019 9571
rect 140961 9531 141019 9537
rect 141145 9571 141203 9577
rect 141145 9537 141157 9571
rect 141191 9537 141203 9571
rect 141145 9531 141203 9537
rect 143005 9571 143063 9577
rect 143005 9537 143017 9571
rect 143051 9568 143063 9571
rect 143261 9571 143319 9577
rect 143051 9540 143212 9568
rect 143051 9537 143063 9540
rect 143005 9531 143063 9537
rect 137925 9503 137983 9509
rect 137925 9469 137937 9503
rect 137971 9469 137983 9503
rect 137925 9463 137983 9469
rect 137428 9336 137784 9364
rect 137428 9324 137434 9336
rect 137830 9324 137836 9376
rect 137888 9364 137894 9376
rect 137940 9364 137968 9463
rect 138934 9460 138940 9512
rect 138992 9500 138998 9512
rect 138992 9472 139440 9500
rect 138992 9460 138998 9472
rect 139302 9432 139308 9444
rect 139263 9404 139308 9432
rect 139302 9392 139308 9404
rect 139360 9392 139366 9444
rect 139412 9432 139440 9472
rect 139486 9460 139492 9512
rect 139544 9500 139550 9512
rect 140976 9500 141004 9531
rect 141694 9500 141700 9512
rect 139544 9472 141700 9500
rect 139544 9460 139550 9472
rect 141694 9460 141700 9472
rect 141752 9460 141758 9512
rect 143184 9500 143212 9540
rect 143261 9537 143273 9571
rect 143307 9568 143319 9571
rect 143442 9568 143448 9580
rect 143307 9540 143448 9568
rect 143307 9537 143319 9540
rect 143261 9531 143319 9537
rect 143442 9528 143448 9540
rect 143500 9528 143506 9580
rect 143534 9528 143540 9580
rect 143592 9568 143598 9580
rect 144362 9568 144368 9580
rect 143592 9540 144368 9568
rect 143592 9528 143598 9540
rect 144362 9528 144368 9540
rect 144420 9528 144426 9580
rect 144845 9571 144903 9577
rect 144845 9537 144857 9571
rect 144891 9568 144903 9571
rect 145006 9568 145012 9580
rect 144891 9540 145012 9568
rect 144891 9537 144903 9540
rect 144845 9531 144903 9537
rect 145006 9528 145012 9540
rect 145064 9528 145070 9580
rect 145116 9509 145144 9608
rect 145466 9596 145472 9648
rect 145524 9636 145530 9648
rect 149146 9636 149152 9648
rect 145524 9608 149152 9636
rect 145524 9596 145530 9608
rect 149146 9596 149152 9608
rect 149204 9596 149210 9648
rect 153930 9636 153936 9648
rect 153891 9608 153936 9636
rect 153930 9596 153936 9608
rect 153988 9596 153994 9648
rect 154040 9608 155080 9636
rect 146869 9571 146927 9577
rect 146869 9537 146881 9571
rect 146915 9568 146927 9571
rect 147306 9568 147312 9580
rect 146915 9540 147312 9568
rect 146915 9537 146927 9540
rect 146869 9531 146927 9537
rect 147306 9528 147312 9540
rect 147364 9528 147370 9580
rect 147841 9571 147899 9577
rect 147841 9537 147853 9571
rect 147887 9568 147899 9571
rect 147887 9540 149284 9568
rect 147887 9537 147899 9540
rect 147841 9531 147899 9537
rect 145101 9503 145159 9509
rect 143184 9472 144132 9500
rect 139412 9404 141924 9432
rect 139854 9364 139860 9376
rect 137888 9336 139860 9364
rect 137888 9324 137894 9336
rect 139854 9324 139860 9336
rect 139912 9324 139918 9376
rect 140774 9364 140780 9376
rect 140735 9336 140780 9364
rect 140774 9324 140780 9336
rect 140832 9324 140838 9376
rect 141896 9373 141924 9404
rect 141881 9367 141939 9373
rect 141881 9333 141893 9367
rect 141927 9364 141939 9367
rect 142154 9364 142160 9376
rect 141927 9336 142160 9364
rect 141927 9333 141939 9336
rect 141881 9327 141939 9333
rect 142154 9324 142160 9336
rect 142212 9324 142218 9376
rect 143718 9364 143724 9376
rect 143679 9336 143724 9364
rect 143718 9324 143724 9336
rect 143776 9324 143782 9376
rect 144104 9364 144132 9472
rect 145101 9469 145113 9503
rect 145147 9500 145159 9503
rect 145190 9500 145196 9512
rect 145147 9472 145196 9500
rect 145147 9469 145159 9472
rect 145101 9463 145159 9469
rect 145190 9460 145196 9472
rect 145248 9500 145254 9512
rect 145650 9500 145656 9512
rect 145248 9472 145656 9500
rect 145248 9460 145254 9472
rect 145650 9460 145656 9472
rect 145708 9460 145714 9512
rect 147122 9500 147128 9512
rect 147083 9472 147128 9500
rect 147122 9460 147128 9472
rect 147180 9500 147186 9512
rect 147585 9503 147643 9509
rect 147585 9500 147597 9503
rect 147180 9472 147597 9500
rect 147180 9460 147186 9472
rect 147585 9469 147597 9472
rect 147631 9469 147643 9503
rect 149256 9500 149284 9540
rect 149330 9528 149336 9580
rect 149388 9568 149394 9580
rect 149425 9571 149483 9577
rect 149425 9568 149437 9571
rect 149388 9540 149437 9568
rect 149388 9528 149394 9540
rect 149425 9537 149437 9540
rect 149471 9537 149483 9571
rect 149425 9531 149483 9537
rect 149514 9528 149520 9580
rect 149572 9568 149578 9580
rect 149609 9571 149667 9577
rect 149609 9568 149621 9571
rect 149572 9540 149621 9568
rect 149572 9528 149578 9540
rect 149609 9537 149621 9540
rect 149655 9537 149667 9571
rect 149609 9531 149667 9537
rect 149716 9540 149928 9568
rect 149716 9500 149744 9540
rect 149256 9472 149744 9500
rect 149900 9500 149928 9540
rect 150986 9528 150992 9580
rect 151044 9568 151050 9580
rect 152090 9568 152096 9580
rect 151044 9540 152096 9568
rect 151044 9528 151050 9540
rect 152090 9528 152096 9540
rect 152148 9528 152154 9580
rect 152389 9574 152447 9577
rect 152389 9571 152504 9574
rect 152389 9537 152401 9571
rect 152435 9568 152504 9571
rect 152550 9568 152556 9580
rect 152435 9546 152556 9568
rect 152435 9537 152447 9546
rect 152476 9540 152556 9546
rect 152389 9531 152447 9537
rect 152550 9528 152556 9540
rect 152608 9528 152614 9580
rect 153286 9568 153292 9580
rect 153247 9540 153292 9568
rect 153286 9528 153292 9540
rect 153344 9528 153350 9580
rect 153654 9528 153660 9580
rect 153712 9568 153718 9580
rect 154040 9568 154068 9608
rect 155052 9580 155080 9608
rect 155310 9596 155316 9648
rect 155368 9636 155374 9648
rect 158272 9636 158300 9664
rect 155368 9608 158300 9636
rect 155368 9596 155374 9608
rect 153712 9540 154068 9568
rect 154131 9569 154189 9575
rect 153712 9528 153718 9540
rect 154131 9535 154143 9569
rect 154177 9535 154189 9569
rect 154131 9529 154189 9535
rect 151446 9500 151452 9512
rect 149900 9472 151452 9500
rect 147585 9463 147643 9469
rect 151446 9460 151452 9472
rect 151504 9460 151510 9512
rect 152642 9460 152648 9512
rect 152700 9500 152706 9512
rect 152700 9472 152793 9500
rect 152700 9460 152706 9472
rect 153010 9460 153016 9512
rect 153068 9500 153074 9512
rect 153470 9500 153476 9512
rect 153068 9472 153476 9500
rect 153068 9460 153074 9472
rect 153470 9460 153476 9472
rect 153528 9460 153534 9512
rect 149146 9392 149152 9444
rect 149204 9432 149210 9444
rect 149204 9404 149652 9432
rect 149204 9392 149210 9404
rect 145558 9364 145564 9376
rect 144104 9336 145564 9364
rect 145558 9324 145564 9336
rect 145616 9324 145622 9376
rect 145742 9364 145748 9376
rect 145703 9336 145748 9364
rect 145742 9324 145748 9336
rect 145800 9364 145806 9376
rect 148870 9364 148876 9376
rect 145800 9336 148876 9364
rect 145800 9324 145806 9336
rect 148870 9324 148876 9336
rect 148928 9324 148934 9376
rect 148965 9367 149023 9373
rect 148965 9333 148977 9367
rect 149011 9364 149023 9367
rect 149514 9364 149520 9376
rect 149011 9336 149520 9364
rect 149011 9333 149023 9336
rect 148965 9327 149023 9333
rect 149514 9324 149520 9336
rect 149572 9324 149578 9376
rect 149624 9364 149652 9404
rect 150526 9392 150532 9444
rect 150584 9432 150590 9444
rect 151630 9432 151636 9444
rect 150584 9404 151636 9432
rect 150584 9392 150590 9404
rect 151630 9392 151636 9404
rect 151688 9392 151694 9444
rect 152660 9432 152688 9460
rect 154132 9444 154160 9529
rect 154666 9528 154672 9580
rect 154724 9568 154730 9580
rect 154945 9571 155003 9577
rect 154945 9568 154957 9571
rect 154724 9540 154957 9568
rect 154724 9528 154730 9540
rect 154945 9537 154957 9540
rect 154991 9537 155003 9571
rect 154945 9531 155003 9537
rect 155034 9528 155040 9580
rect 155092 9568 155098 9580
rect 155092 9540 155185 9568
rect 155092 9528 155098 9540
rect 156138 9528 156144 9580
rect 156196 9568 156202 9580
rect 156196 9540 156241 9568
rect 156196 9528 156202 9540
rect 156322 9528 156328 9580
rect 156380 9568 156386 9580
rect 156969 9571 157027 9577
rect 156969 9568 156981 9571
rect 156380 9540 156981 9568
rect 156380 9528 156386 9540
rect 156969 9537 156981 9540
rect 157015 9537 157027 9571
rect 157794 9568 157800 9580
rect 157755 9540 157800 9568
rect 156969 9531 157027 9537
rect 157794 9528 157800 9540
rect 157852 9528 157858 9580
rect 154298 9460 154304 9512
rect 154356 9500 154362 9512
rect 154356 9472 154401 9500
rect 154356 9460 154362 9472
rect 154758 9460 154764 9512
rect 154816 9500 154822 9512
rect 155494 9500 155500 9512
rect 154816 9472 155500 9500
rect 154816 9460 154822 9472
rect 155494 9460 155500 9472
rect 155552 9460 155558 9512
rect 155862 9460 155868 9512
rect 155920 9500 155926 9512
rect 155957 9503 156015 9509
rect 155957 9500 155969 9503
rect 155920 9472 155969 9500
rect 155920 9460 155926 9472
rect 155957 9469 155969 9472
rect 156003 9469 156015 9503
rect 155957 9463 156015 9469
rect 156785 9503 156843 9509
rect 156785 9469 156797 9503
rect 156831 9469 156843 9503
rect 156785 9463 156843 9469
rect 154022 9432 154028 9444
rect 152660 9404 154028 9432
rect 154022 9392 154028 9404
rect 154080 9392 154086 9444
rect 154114 9392 154120 9444
rect 154172 9392 154178 9444
rect 152274 9364 152280 9376
rect 149624 9336 152280 9364
rect 152274 9324 152280 9336
rect 152332 9324 152338 9376
rect 153102 9364 153108 9376
rect 153063 9336 153108 9364
rect 153102 9324 153108 9336
rect 153160 9324 153166 9376
rect 153838 9324 153844 9376
rect 153896 9364 153902 9376
rect 154761 9367 154819 9373
rect 154761 9364 154773 9367
rect 153896 9336 154773 9364
rect 153896 9324 153902 9336
rect 154761 9333 154773 9336
rect 154807 9333 154819 9367
rect 155880 9364 155908 9460
rect 156800 9432 156828 9463
rect 156966 9432 156972 9444
rect 156800 9404 156972 9432
rect 156966 9392 156972 9404
rect 157024 9392 157030 9444
rect 157978 9432 157984 9444
rect 157306 9404 157984 9432
rect 156230 9364 156236 9376
rect 155880 9336 156236 9364
rect 154761 9327 154819 9333
rect 156230 9324 156236 9336
rect 156288 9324 156294 9376
rect 156325 9367 156383 9373
rect 156325 9333 156337 9367
rect 156371 9364 156383 9367
rect 157058 9364 157064 9376
rect 156371 9336 157064 9364
rect 156371 9333 156383 9336
rect 156325 9327 156383 9333
rect 157058 9324 157064 9336
rect 157116 9324 157122 9376
rect 157153 9367 157211 9373
rect 157153 9333 157165 9367
rect 157199 9364 157211 9367
rect 157306 9364 157334 9404
rect 157978 9392 157984 9404
rect 158036 9392 158042 9444
rect 157199 9336 157334 9364
rect 157199 9333 157211 9336
rect 157153 9327 157211 9333
rect 157518 9324 157524 9376
rect 157576 9364 157582 9376
rect 157613 9367 157671 9373
rect 157613 9364 157625 9367
rect 157576 9336 157625 9364
rect 157576 9324 157582 9336
rect 157613 9333 157625 9336
rect 157659 9333 157671 9367
rect 157613 9327 157671 9333
rect 1104 9274 158884 9296
rect 1104 9222 20672 9274
rect 20724 9222 20736 9274
rect 20788 9222 20800 9274
rect 20852 9222 20864 9274
rect 20916 9222 20928 9274
rect 20980 9222 60117 9274
rect 60169 9222 60181 9274
rect 60233 9222 60245 9274
rect 60297 9222 60309 9274
rect 60361 9222 60373 9274
rect 60425 9222 99562 9274
rect 99614 9222 99626 9274
rect 99678 9222 99690 9274
rect 99742 9222 99754 9274
rect 99806 9222 99818 9274
rect 99870 9222 139007 9274
rect 139059 9222 139071 9274
rect 139123 9222 139135 9274
rect 139187 9222 139199 9274
rect 139251 9222 139263 9274
rect 139315 9222 158884 9274
rect 1104 9200 158884 9222
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 11054 9160 11060 9172
rect 4019 9132 11060 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 11054 9120 11060 9132
rect 11112 9160 11118 9172
rect 13725 9163 13783 9169
rect 11112 9132 13400 9160
rect 11112 9120 11118 9132
rect 10686 9092 10692 9104
rect 10647 9064 10692 9092
rect 10686 9052 10692 9064
rect 10744 9092 10750 9104
rect 10744 9064 11284 9092
rect 10744 9052 10750 9064
rect 11256 9033 11284 9064
rect 11241 9027 11299 9033
rect 11241 8993 11253 9027
rect 11287 8993 11299 9027
rect 11241 8987 11299 8993
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 5810 8956 5816 8968
rect 5399 8928 5816 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 11422 8956 11428 8968
rect 11383 8928 11428 8956
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8956 12403 8959
rect 12434 8956 12440 8968
rect 12391 8928 12440 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 5108 8891 5166 8897
rect 5108 8857 5120 8891
rect 5154 8888 5166 8891
rect 5258 8888 5264 8900
rect 5154 8860 5264 8888
rect 5154 8857 5166 8860
rect 5108 8851 5166 8857
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 12590 8891 12648 8897
rect 12590 8888 12602 8891
rect 12406 8860 12602 8888
rect 12406 8832 12434 8860
rect 12590 8857 12602 8860
rect 12636 8857 12648 8891
rect 13372 8888 13400 9132
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 17678 9160 17684 9172
rect 13771 9132 17684 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 19444 9132 21373 9160
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18598 9092 18604 9104
rect 17828 9064 18604 9092
rect 17828 9052 17834 9064
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 19444 9036 19472 9132
rect 21361 9129 21373 9132
rect 21407 9160 21419 9163
rect 26326 9160 26332 9172
rect 21407 9132 26332 9160
rect 21407 9129 21419 9132
rect 21361 9123 21419 9129
rect 26326 9120 26332 9132
rect 26384 9160 26390 9172
rect 26421 9163 26479 9169
rect 26421 9160 26433 9163
rect 26384 9132 26433 9160
rect 26384 9120 26390 9132
rect 26421 9129 26433 9132
rect 26467 9129 26479 9163
rect 26421 9123 26479 9129
rect 26510 9120 26516 9172
rect 26568 9160 26574 9172
rect 26568 9132 38148 9160
rect 26568 9120 26574 9132
rect 29181 9095 29239 9101
rect 29181 9061 29193 9095
rect 29227 9092 29239 9095
rect 29730 9092 29736 9104
rect 29227 9064 29736 9092
rect 29227 9061 29239 9064
rect 29181 9055 29239 9061
rect 29730 9052 29736 9064
rect 29788 9052 29794 9104
rect 33137 9095 33195 9101
rect 33137 9061 33149 9095
rect 33183 9092 33195 9095
rect 38120 9092 38148 9132
rect 38654 9120 38660 9172
rect 38712 9160 38718 9172
rect 39390 9160 39396 9172
rect 38712 9132 39396 9160
rect 38712 9120 38718 9132
rect 39390 9120 39396 9132
rect 39448 9160 39454 9172
rect 43901 9163 43959 9169
rect 39448 9132 41828 9160
rect 39448 9120 39454 9132
rect 40218 9092 40224 9104
rect 33183 9064 35756 9092
rect 38120 9064 40224 9092
rect 33183 9061 33195 9064
rect 33137 9055 33195 9061
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 14274 9024 14280 9036
rect 13504 8996 14280 9024
rect 13504 8984 13510 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 15102 9024 15108 9036
rect 15063 8996 15108 9024
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 16942 9024 16948 9036
rect 16903 8996 16948 9024
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 19426 9024 19432 9036
rect 17736 8996 18000 9024
rect 19339 8996 19432 9024
rect 17736 8984 17742 8996
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8956 14519 8959
rect 16758 8956 16764 8968
rect 14507 8928 16764 8956
rect 14507 8925 14519 8928
rect 14461 8919 14519 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8925 17187 8959
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 17129 8919 17187 8925
rect 15372 8891 15430 8897
rect 13372 8860 15332 8888
rect 12590 8851 12648 8857
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 12158 8820 12164 8832
rect 11655 8792 12164 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12342 8780 12348 8832
rect 12400 8792 12434 8832
rect 12400 8780 12406 8792
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 14424 8792 14657 8820
rect 14424 8780 14430 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 15304 8820 15332 8860
rect 15372 8857 15384 8891
rect 15418 8888 15430 8891
rect 15654 8888 15660 8900
rect 15418 8860 15660 8888
rect 15418 8857 15430 8860
rect 15372 8851 15430 8857
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 17144 8888 17172 8919
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 17972 8965 18000 8996
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 27614 9024 27620 9036
rect 22066 8996 27620 9024
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 21174 8956 21180 8968
rect 18187 8928 21180 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 17586 8888 17592 8900
rect 17144 8860 17592 8888
rect 17586 8848 17592 8860
rect 17644 8888 17650 8900
rect 17644 8860 18736 8888
rect 17644 8848 17650 8860
rect 18708 8832 18736 8860
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19674 8891 19732 8897
rect 19674 8888 19686 8891
rect 19392 8860 19686 8888
rect 19392 8848 19398 8860
rect 19674 8857 19686 8860
rect 19720 8857 19732 8891
rect 22066 8888 22094 8996
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 27706 8984 27712 9036
rect 27764 9024 27770 9036
rect 27801 9027 27859 9033
rect 27801 9024 27813 9027
rect 27764 8996 27813 9024
rect 27764 8984 27770 8996
rect 27801 8993 27813 8996
rect 27847 8993 27859 9027
rect 27801 8987 27859 8993
rect 31662 8984 31668 9036
rect 31720 9024 31726 9036
rect 31757 9027 31815 9033
rect 31757 9024 31769 9027
rect 31720 8996 31769 9024
rect 31720 8984 31726 8996
rect 31757 8993 31769 8996
rect 31803 8993 31815 9027
rect 31757 8987 31815 8993
rect 33226 8984 33232 9036
rect 33284 9024 33290 9036
rect 33594 9024 33600 9036
rect 33284 8996 33600 9024
rect 33284 8984 33290 8996
rect 33594 8984 33600 8996
rect 33652 9024 33658 9036
rect 33965 9027 34023 9033
rect 33965 9024 33977 9027
rect 33652 8996 33977 9024
rect 33652 8984 33658 8996
rect 33965 8993 33977 8996
rect 34011 8993 34023 9027
rect 33965 8987 34023 8993
rect 27154 8956 27160 8968
rect 27115 8928 27160 8956
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 27264 8928 27936 8956
rect 19674 8851 19732 8857
rect 19812 8860 22094 8888
rect 16114 8820 16120 8832
rect 15304 8792 16120 8820
rect 14645 8783 14703 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17313 8823 17371 8829
rect 17313 8789 17325 8823
rect 17359 8820 17371 8823
rect 18046 8820 18052 8832
rect 17359 8792 18052 8820
rect 17359 8789 17371 8792
rect 17313 8783 17371 8789
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18690 8780 18696 8832
rect 18748 8820 18754 8832
rect 19812 8820 19840 8860
rect 18748 8792 19840 8820
rect 20809 8823 20867 8829
rect 18748 8780 18754 8792
rect 20809 8789 20821 8823
rect 20855 8820 20867 8823
rect 20990 8820 20996 8832
rect 20855 8792 20996 8820
rect 20855 8789 20867 8792
rect 20809 8783 20867 8789
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 26050 8780 26056 8832
rect 26108 8820 26114 8832
rect 27264 8820 27292 8928
rect 27908 8888 27936 8928
rect 29086 8916 29092 8968
rect 29144 8956 29150 8968
rect 29733 8959 29791 8965
rect 29733 8956 29745 8959
rect 29144 8928 29745 8956
rect 29144 8916 29150 8928
rect 29733 8925 29745 8928
rect 29779 8925 29791 8959
rect 29733 8919 29791 8925
rect 30466 8916 30472 8968
rect 30524 8956 30530 8968
rect 32858 8956 32864 8968
rect 30524 8928 32864 8956
rect 30524 8916 30530 8928
rect 32858 8916 32864 8928
rect 32916 8916 32922 8968
rect 32950 8916 32956 8968
rect 33008 8956 33014 8968
rect 33781 8959 33839 8965
rect 33781 8956 33793 8959
rect 33008 8928 33793 8956
rect 33008 8916 33014 8928
rect 33781 8925 33793 8928
rect 33827 8925 33839 8959
rect 35728 8956 35756 9064
rect 40218 9052 40224 9064
rect 40276 9052 40282 9104
rect 36722 9024 36728 9036
rect 36683 8996 36728 9024
rect 36722 8984 36728 8996
rect 36780 9024 36786 9036
rect 41800 9033 41828 9132
rect 43901 9129 43913 9163
rect 43947 9160 43959 9163
rect 44726 9160 44732 9172
rect 43947 9132 44732 9160
rect 43947 9129 43959 9132
rect 43901 9123 43959 9129
rect 44726 9120 44732 9132
rect 44784 9120 44790 9172
rect 45462 9120 45468 9172
rect 45520 9160 45526 9172
rect 48685 9163 48743 9169
rect 45520 9132 48636 9160
rect 45520 9120 45526 9132
rect 47026 9052 47032 9104
rect 47084 9092 47090 9104
rect 47213 9095 47271 9101
rect 47213 9092 47225 9095
rect 47084 9064 47225 9092
rect 47084 9052 47090 9064
rect 47213 9061 47225 9064
rect 47259 9092 47271 9095
rect 48314 9092 48320 9104
rect 47259 9064 48320 9092
rect 47259 9061 47271 9064
rect 47213 9055 47271 9061
rect 48314 9052 48320 9064
rect 48372 9052 48378 9104
rect 48608 9092 48636 9132
rect 48685 9129 48697 9163
rect 48731 9160 48743 9163
rect 49602 9160 49608 9172
rect 48731 9132 49608 9160
rect 48731 9129 48743 9132
rect 48685 9123 48743 9129
rect 49602 9120 49608 9132
rect 49660 9120 49666 9172
rect 49694 9120 49700 9172
rect 49752 9160 49758 9172
rect 53374 9160 53380 9172
rect 49752 9132 53236 9160
rect 53335 9132 53380 9160
rect 49752 9120 49758 9132
rect 49418 9092 49424 9104
rect 48608 9064 49424 9092
rect 49418 9052 49424 9064
rect 49476 9052 49482 9104
rect 49510 9052 49516 9104
rect 49568 9092 49574 9104
rect 49789 9095 49847 9101
rect 49789 9092 49801 9095
rect 49568 9064 49801 9092
rect 49568 9052 49574 9064
rect 49789 9061 49801 9064
rect 49835 9061 49847 9095
rect 49789 9055 49847 9061
rect 49878 9052 49884 9104
rect 49936 9092 49942 9104
rect 53208 9092 53236 9132
rect 53374 9120 53380 9132
rect 53432 9120 53438 9172
rect 55677 9163 55735 9169
rect 55677 9160 55689 9163
rect 53760 9132 55689 9160
rect 53760 9092 53788 9132
rect 55677 9129 55689 9132
rect 55723 9129 55735 9163
rect 55677 9123 55735 9129
rect 49936 9064 50752 9092
rect 53208 9064 53788 9092
rect 49936 9052 49942 9064
rect 37185 9027 37243 9033
rect 37185 9024 37197 9027
rect 36780 8996 37197 9024
rect 36780 8984 36786 8996
rect 37185 8993 37197 8996
rect 37231 8993 37243 9027
rect 37185 8987 37243 8993
rect 41785 9027 41843 9033
rect 41785 8993 41797 9027
rect 41831 9024 41843 9027
rect 45554 9024 45560 9036
rect 41831 8996 42656 9024
rect 41831 8993 41843 8996
rect 41785 8987 41843 8993
rect 41046 8956 41052 8968
rect 35728 8928 41052 8956
rect 33781 8919 33839 8925
rect 41046 8916 41052 8928
rect 41104 8916 41110 8968
rect 41690 8916 41696 8968
rect 41748 8956 41754 8968
rect 42521 8959 42579 8965
rect 42521 8956 42533 8959
rect 41748 8928 42533 8956
rect 41748 8916 41754 8928
rect 42521 8925 42533 8928
rect 42567 8925 42579 8959
rect 42628 8956 42656 8996
rect 45204 8996 45560 9024
rect 43162 8956 43168 8968
rect 42628 8928 43168 8956
rect 42521 8919 42579 8925
rect 43162 8916 43168 8928
rect 43220 8956 43226 8968
rect 43990 8956 43996 8968
rect 43220 8928 43996 8956
rect 43220 8916 43226 8928
rect 43990 8916 43996 8928
rect 44048 8916 44054 8968
rect 45204 8965 45232 8996
rect 45554 8984 45560 8996
rect 45612 8984 45618 9036
rect 47670 8984 47676 9036
rect 47728 9024 47734 9036
rect 50338 9024 50344 9036
rect 47728 8996 50344 9024
rect 47728 8984 47734 8996
rect 50338 8984 50344 8996
rect 50396 8984 50402 9036
rect 50724 9033 50752 9064
rect 54202 9052 54208 9104
rect 54260 9092 54266 9104
rect 55692 9092 55720 9123
rect 55858 9120 55864 9172
rect 55916 9160 55922 9172
rect 56870 9160 56876 9172
rect 55916 9132 56876 9160
rect 55916 9120 55922 9132
rect 56870 9120 56876 9132
rect 56928 9120 56934 9172
rect 56962 9120 56968 9172
rect 57020 9160 57026 9172
rect 57057 9163 57115 9169
rect 57057 9160 57069 9163
rect 57020 9132 57069 9160
rect 57020 9120 57026 9132
rect 57057 9129 57069 9132
rect 57103 9129 57115 9163
rect 57057 9123 57115 9129
rect 59814 9120 59820 9172
rect 59872 9160 59878 9172
rect 64509 9163 64567 9169
rect 64509 9160 64521 9163
rect 59872 9132 64521 9160
rect 59872 9120 59878 9132
rect 64509 9129 64521 9132
rect 64555 9160 64567 9163
rect 64874 9160 64880 9172
rect 64555 9132 64880 9160
rect 64555 9129 64567 9132
rect 64509 9123 64567 9129
rect 64874 9120 64880 9132
rect 64932 9120 64938 9172
rect 64966 9120 64972 9172
rect 65024 9160 65030 9172
rect 65153 9163 65211 9169
rect 65153 9160 65165 9163
rect 65024 9132 65165 9160
rect 65024 9120 65030 9132
rect 65153 9129 65165 9132
rect 65199 9129 65211 9163
rect 67177 9163 67235 9169
rect 65153 9123 65211 9129
rect 65812 9132 66852 9160
rect 57698 9092 57704 9104
rect 54260 9064 55628 9092
rect 55692 9064 57704 9092
rect 54260 9052 54266 9064
rect 50709 9027 50767 9033
rect 50709 8993 50721 9027
rect 50755 8993 50767 9027
rect 50709 8987 50767 8993
rect 54018 8984 54024 9036
rect 54076 9024 54082 9036
rect 55600 9024 55628 9064
rect 57698 9052 57704 9064
rect 57756 9052 57762 9104
rect 59081 9095 59139 9101
rect 59081 9061 59093 9095
rect 59127 9092 59139 9095
rect 60642 9092 60648 9104
rect 59127 9064 60648 9092
rect 59127 9061 59139 9064
rect 59081 9055 59139 9061
rect 60642 9052 60648 9064
rect 60700 9052 60706 9104
rect 63494 9052 63500 9104
rect 63552 9092 63558 9104
rect 65812 9092 65840 9132
rect 63552 9064 65840 9092
rect 63552 9052 63558 9064
rect 62114 9024 62120 9036
rect 54076 8996 54524 9024
rect 55600 8996 57836 9024
rect 62075 8996 62120 9024
rect 54076 8984 54082 8996
rect 45189 8959 45247 8965
rect 45189 8925 45201 8959
rect 45235 8925 45247 8959
rect 45189 8919 45247 8925
rect 45370 8916 45376 8968
rect 45428 8956 45434 8968
rect 45833 8959 45891 8965
rect 45833 8956 45845 8959
rect 45428 8928 45845 8956
rect 45428 8916 45434 8928
rect 45833 8925 45845 8928
rect 45879 8956 45891 8959
rect 46658 8956 46664 8968
rect 45879 8928 46664 8956
rect 45879 8925 45891 8928
rect 45833 8919 45891 8925
rect 46658 8916 46664 8928
rect 46716 8916 46722 8968
rect 48406 8916 48412 8968
rect 48464 8956 48470 8968
rect 53374 8956 53380 8968
rect 48464 8928 53380 8956
rect 48464 8916 48470 8928
rect 53374 8916 53380 8928
rect 53432 8916 53438 8968
rect 53561 8959 53619 8965
rect 53561 8925 53573 8959
rect 53607 8956 53619 8959
rect 53834 8956 53840 8968
rect 53607 8928 53840 8956
rect 53607 8925 53619 8928
rect 53561 8919 53619 8925
rect 53834 8916 53840 8928
rect 53892 8956 53898 8968
rect 54110 8956 54116 8968
rect 53892 8928 54116 8956
rect 53892 8916 53898 8928
rect 54110 8916 54116 8928
rect 54168 8916 54174 8968
rect 54294 8956 54300 8968
rect 54255 8928 54300 8956
rect 54294 8916 54300 8928
rect 54352 8916 54358 8968
rect 54496 8965 54524 8996
rect 57808 8968 57836 8996
rect 62114 8984 62120 8996
rect 62172 8984 62178 9036
rect 54481 8959 54539 8965
rect 54481 8925 54493 8959
rect 54527 8925 54539 8959
rect 54481 8919 54539 8925
rect 55398 8916 55404 8968
rect 55456 8956 55462 8968
rect 56229 8959 56287 8965
rect 56229 8956 56241 8959
rect 55456 8928 56241 8956
rect 55456 8916 55462 8928
rect 56229 8925 56241 8928
rect 56275 8925 56287 8959
rect 56229 8919 56287 8925
rect 57241 8959 57299 8965
rect 57241 8925 57253 8959
rect 57287 8925 57299 8959
rect 57698 8956 57704 8968
rect 57659 8928 57704 8956
rect 57241 8919 57299 8925
rect 28046 8891 28104 8897
rect 28046 8888 28058 8891
rect 27908 8860 28058 8888
rect 28046 8857 28058 8860
rect 28092 8857 28104 8891
rect 29978 8891 30036 8897
rect 29978 8888 29990 8891
rect 28046 8851 28104 8857
rect 28653 8860 29990 8888
rect 26108 8792 27292 8820
rect 27341 8823 27399 8829
rect 26108 8780 26114 8792
rect 27341 8789 27353 8823
rect 27387 8820 27399 8823
rect 28653 8820 28681 8860
rect 29978 8857 29990 8860
rect 30024 8857 30036 8891
rect 29978 8851 30036 8857
rect 32024 8891 32082 8897
rect 32024 8857 32036 8891
rect 32070 8888 32082 8891
rect 32398 8888 32404 8900
rect 32070 8860 32404 8888
rect 32070 8857 32082 8860
rect 32024 8851 32082 8857
rect 32398 8848 32404 8860
rect 32456 8848 32462 8900
rect 33686 8888 33692 8900
rect 33428 8860 33692 8888
rect 27387 8792 28681 8820
rect 31113 8823 31171 8829
rect 27387 8789 27399 8792
rect 27341 8783 27399 8789
rect 31113 8789 31125 8823
rect 31159 8820 31171 8823
rect 33428 8820 33456 8860
rect 33686 8848 33692 8860
rect 33744 8848 33750 8900
rect 36480 8891 36538 8897
rect 36480 8857 36492 8891
rect 36526 8888 36538 8891
rect 37274 8888 37280 8900
rect 36526 8860 37280 8888
rect 36526 8857 36538 8860
rect 36480 8851 36538 8857
rect 37274 8848 37280 8860
rect 37332 8848 37338 8900
rect 37452 8891 37510 8897
rect 37452 8857 37464 8891
rect 37498 8888 37510 8891
rect 40954 8888 40960 8900
rect 37498 8860 40960 8888
rect 37498 8857 37510 8860
rect 37452 8851 37510 8857
rect 40954 8848 40960 8860
rect 41012 8848 41018 8900
rect 41506 8888 41512 8900
rect 41564 8897 41570 8900
rect 41476 8860 41512 8888
rect 41506 8848 41512 8860
rect 41564 8851 41576 8897
rect 41564 8848 41570 8851
rect 41874 8848 41880 8900
rect 41932 8888 41938 8900
rect 42766 8891 42824 8897
rect 42766 8888 42778 8891
rect 41932 8860 42778 8888
rect 41932 8848 41938 8860
rect 42766 8857 42778 8860
rect 42812 8857 42824 8891
rect 45462 8888 45468 8900
rect 42766 8851 42824 8857
rect 45296 8860 45468 8888
rect 33594 8820 33600 8832
rect 31159 8792 33456 8820
rect 33555 8792 33600 8820
rect 31159 8789 31171 8792
rect 31113 8783 31171 8789
rect 33594 8780 33600 8792
rect 33652 8780 33658 8832
rect 34146 8780 34152 8832
rect 34204 8820 34210 8832
rect 35345 8823 35403 8829
rect 35345 8820 35357 8823
rect 34204 8792 35357 8820
rect 34204 8780 34210 8792
rect 35345 8789 35357 8792
rect 35391 8820 35403 8823
rect 38010 8820 38016 8832
rect 35391 8792 38016 8820
rect 35391 8789 35403 8792
rect 35345 8783 35403 8789
rect 38010 8780 38016 8792
rect 38068 8780 38074 8832
rect 38565 8823 38623 8829
rect 38565 8789 38577 8823
rect 38611 8820 38623 8823
rect 39758 8820 39764 8832
rect 38611 8792 39764 8820
rect 38611 8789 38623 8792
rect 38565 8783 38623 8789
rect 39758 8780 39764 8792
rect 39816 8780 39822 8832
rect 40034 8780 40040 8832
rect 40092 8820 40098 8832
rect 40405 8823 40463 8829
rect 40405 8820 40417 8823
rect 40092 8792 40417 8820
rect 40092 8780 40098 8792
rect 40405 8789 40417 8792
rect 40451 8789 40463 8823
rect 40405 8783 40463 8789
rect 41046 8780 41052 8832
rect 41104 8820 41110 8832
rect 44174 8820 44180 8832
rect 41104 8792 44180 8820
rect 41104 8780 41110 8792
rect 44174 8780 44180 8792
rect 44232 8780 44238 8832
rect 44637 8823 44695 8829
rect 44637 8789 44649 8823
rect 44683 8820 44695 8823
rect 45296 8820 45324 8860
rect 45462 8848 45468 8860
rect 45520 8848 45526 8900
rect 45554 8848 45560 8900
rect 45612 8888 45618 8900
rect 46078 8891 46136 8897
rect 46078 8888 46090 8891
rect 45612 8860 46090 8888
rect 45612 8848 45618 8860
rect 46078 8857 46090 8860
rect 46124 8857 46136 8891
rect 50954 8891 51012 8897
rect 50954 8888 50966 8891
rect 46078 8851 46136 8857
rect 48056 8860 50966 8888
rect 44683 8792 45324 8820
rect 45373 8823 45431 8829
rect 44683 8789 44695 8792
rect 44637 8783 44695 8789
rect 45373 8789 45385 8823
rect 45419 8820 45431 8823
rect 46382 8820 46388 8832
rect 45419 8792 46388 8820
rect 45419 8789 45431 8792
rect 45373 8783 45431 8789
rect 46382 8780 46388 8792
rect 46440 8780 46446 8832
rect 47210 8780 47216 8832
rect 47268 8820 47274 8832
rect 48056 8829 48084 8860
rect 50954 8857 50966 8860
rect 51000 8857 51012 8891
rect 57256 8888 57284 8919
rect 57698 8916 57704 8928
rect 57756 8916 57762 8968
rect 57790 8916 57796 8968
rect 57848 8916 57854 8968
rect 57974 8965 57980 8968
rect 57968 8919 57980 8965
rect 58032 8956 58038 8968
rect 58032 8928 58068 8956
rect 57974 8916 57980 8919
rect 58032 8916 58038 8928
rect 61654 8916 61660 8968
rect 61712 8956 61718 8968
rect 61712 8928 62804 8956
rect 61712 8916 61718 8928
rect 58158 8888 58164 8900
rect 50954 8851 51012 8857
rect 51046 8860 56548 8888
rect 57256 8860 58164 8888
rect 48041 8823 48099 8829
rect 48041 8820 48053 8823
rect 47268 8792 48053 8820
rect 47268 8780 47274 8792
rect 48041 8789 48053 8792
rect 48087 8789 48099 8823
rect 49234 8820 49240 8832
rect 49195 8792 49240 8820
rect 48041 8783 48099 8789
rect 49234 8780 49240 8792
rect 49292 8820 49298 8832
rect 49970 8820 49976 8832
rect 49292 8792 49976 8820
rect 49292 8780 49298 8792
rect 49970 8780 49976 8792
rect 50028 8780 50034 8832
rect 50062 8780 50068 8832
rect 50120 8820 50126 8832
rect 50798 8820 50804 8832
rect 50120 8792 50804 8820
rect 50120 8780 50126 8792
rect 50798 8780 50804 8792
rect 50856 8820 50862 8832
rect 51046 8820 51074 8860
rect 50856 8792 51074 8820
rect 52089 8823 52147 8829
rect 50856 8780 50862 8792
rect 52089 8789 52101 8823
rect 52135 8820 52147 8823
rect 52730 8820 52736 8832
rect 52135 8792 52736 8820
rect 52135 8789 52147 8792
rect 52089 8783 52147 8789
rect 52730 8780 52736 8792
rect 52788 8780 52794 8832
rect 52825 8823 52883 8829
rect 52825 8789 52837 8823
rect 52871 8820 52883 8823
rect 53466 8820 53472 8832
rect 52871 8792 53472 8820
rect 52871 8789 52883 8792
rect 52825 8783 52883 8789
rect 53466 8780 53472 8792
rect 53524 8820 53530 8832
rect 54570 8820 54576 8832
rect 53524 8792 54576 8820
rect 53524 8780 53530 8792
rect 54570 8780 54576 8792
rect 54628 8780 54634 8832
rect 54665 8823 54723 8829
rect 54665 8789 54677 8823
rect 54711 8820 54723 8823
rect 54938 8820 54944 8832
rect 54711 8792 54944 8820
rect 54711 8789 54723 8792
rect 54665 8783 54723 8789
rect 54938 8780 54944 8792
rect 54996 8780 55002 8832
rect 56410 8820 56416 8832
rect 56371 8792 56416 8820
rect 56410 8780 56416 8792
rect 56468 8780 56474 8832
rect 56520 8820 56548 8860
rect 58158 8848 58164 8860
rect 58216 8848 58222 8900
rect 60826 8888 60832 8900
rect 60739 8860 60832 8888
rect 60826 8848 60832 8860
rect 60884 8888 60890 8900
rect 61746 8888 61752 8900
rect 60884 8860 61752 8888
rect 60884 8848 60890 8860
rect 61746 8848 61752 8860
rect 61804 8848 61810 8900
rect 62384 8891 62442 8897
rect 62384 8857 62396 8891
rect 62430 8888 62442 8891
rect 62666 8888 62672 8900
rect 62430 8860 62672 8888
rect 62430 8857 62442 8860
rect 62384 8851 62442 8857
rect 62666 8848 62672 8860
rect 62724 8848 62730 8900
rect 62776 8888 62804 8928
rect 65242 8916 65248 8968
rect 65300 8956 65306 8968
rect 65794 8956 65800 8968
rect 65300 8928 65800 8956
rect 65300 8916 65306 8928
rect 65794 8916 65800 8928
rect 65852 8916 65858 8968
rect 65886 8916 65892 8968
rect 65944 8956 65950 8968
rect 66053 8959 66111 8965
rect 66053 8956 66065 8959
rect 65944 8928 66065 8956
rect 65944 8916 65950 8928
rect 66053 8925 66065 8928
rect 66099 8925 66111 8959
rect 66824 8956 66852 9132
rect 67177 9129 67189 9163
rect 67223 9160 67235 9163
rect 69014 9160 69020 9172
rect 67223 9132 69020 9160
rect 67223 9129 67235 9132
rect 67177 9123 67235 9129
rect 69014 9120 69020 9132
rect 69072 9120 69078 9172
rect 74445 9163 74503 9169
rect 74445 9129 74457 9163
rect 74491 9160 74503 9163
rect 75914 9160 75920 9172
rect 74491 9132 75920 9160
rect 74491 9129 74503 9132
rect 74445 9123 74503 9129
rect 75914 9120 75920 9132
rect 75972 9120 75978 9172
rect 82630 9160 82636 9172
rect 76024 9132 82636 9160
rect 69750 9052 69756 9104
rect 69808 9092 69814 9104
rect 76024 9092 76052 9132
rect 82630 9120 82636 9132
rect 82688 9120 82694 9172
rect 82722 9120 82728 9172
rect 82780 9160 82786 9172
rect 87785 9163 87843 9169
rect 82780 9132 87368 9160
rect 82780 9120 82786 9132
rect 69808 9064 76052 9092
rect 69808 9052 69814 9064
rect 83918 9052 83924 9104
rect 83976 9092 83982 9104
rect 85390 9092 85396 9104
rect 83976 9064 85396 9092
rect 83976 9052 83982 9064
rect 85390 9052 85396 9064
rect 85448 9052 85454 9104
rect 87340 9092 87368 9132
rect 87785 9129 87797 9163
rect 87831 9160 87843 9163
rect 88150 9160 88156 9172
rect 87831 9132 88156 9160
rect 87831 9129 87843 9132
rect 87785 9123 87843 9129
rect 88150 9120 88156 9132
rect 88208 9120 88214 9172
rect 88334 9120 88340 9172
rect 88392 9160 88398 9172
rect 88797 9163 88855 9169
rect 88797 9160 88809 9163
rect 88392 9132 88809 9160
rect 88392 9120 88398 9132
rect 88797 9129 88809 9132
rect 88843 9160 88855 9163
rect 90818 9160 90824 9172
rect 88843 9132 90824 9160
rect 88843 9129 88855 9132
rect 88797 9123 88855 9129
rect 90818 9120 90824 9132
rect 90876 9120 90882 9172
rect 90910 9120 90916 9172
rect 90968 9160 90974 9172
rect 101030 9160 101036 9172
rect 90968 9132 101036 9160
rect 90968 9120 90974 9132
rect 101030 9120 101036 9132
rect 101088 9120 101094 9172
rect 101214 9160 101220 9172
rect 101175 9132 101220 9160
rect 101214 9120 101220 9132
rect 101272 9120 101278 9172
rect 103238 9120 103244 9172
rect 103296 9160 103302 9172
rect 114462 9160 114468 9172
rect 103296 9132 114468 9160
rect 103296 9120 103302 9132
rect 114462 9120 114468 9132
rect 114520 9120 114526 9172
rect 114922 9160 114928 9172
rect 114883 9132 114928 9160
rect 114922 9120 114928 9132
rect 114980 9120 114986 9172
rect 115477 9163 115535 9169
rect 115477 9129 115489 9163
rect 115523 9160 115535 9163
rect 115566 9160 115572 9172
rect 115523 9132 115572 9160
rect 115523 9129 115535 9132
rect 115477 9123 115535 9129
rect 115566 9120 115572 9132
rect 115624 9120 115630 9172
rect 115842 9120 115848 9172
rect 115900 9160 115906 9172
rect 117961 9163 118019 9169
rect 117961 9160 117973 9163
rect 115900 9132 117973 9160
rect 115900 9120 115906 9132
rect 117961 9129 117973 9132
rect 118007 9129 118019 9163
rect 117961 9123 118019 9129
rect 118326 9120 118332 9172
rect 118384 9160 118390 9172
rect 128262 9160 128268 9172
rect 118384 9132 128268 9160
rect 118384 9120 118390 9132
rect 128262 9120 128268 9132
rect 128320 9120 128326 9172
rect 130930 9160 130936 9172
rect 129200 9132 130936 9160
rect 89622 9092 89628 9104
rect 87340 9064 89628 9092
rect 89622 9052 89628 9064
rect 89680 9052 89686 9104
rect 71130 8984 71136 9036
rect 71188 9024 71194 9036
rect 71188 8996 75316 9024
rect 71188 8984 71194 8996
rect 68097 8959 68155 8965
rect 68097 8956 68109 8959
rect 66824 8928 68109 8956
rect 66053 8919 66111 8925
rect 68097 8925 68109 8928
rect 68143 8956 68155 8959
rect 68833 8959 68891 8965
rect 68833 8956 68845 8959
rect 68143 8928 68845 8956
rect 68143 8925 68155 8928
rect 68097 8919 68155 8925
rect 68833 8925 68845 8928
rect 68879 8925 68891 8959
rect 68833 8919 68891 8925
rect 75089 8959 75147 8965
rect 75089 8925 75101 8959
rect 75135 8956 75147 8959
rect 75178 8956 75184 8968
rect 75135 8928 75184 8956
rect 75135 8925 75147 8928
rect 75089 8919 75147 8925
rect 75178 8916 75184 8928
rect 75236 8916 75242 8968
rect 69842 8888 69848 8900
rect 62776 8860 69848 8888
rect 69842 8848 69848 8860
rect 69900 8848 69906 8900
rect 71682 8848 71688 8900
rect 71740 8888 71746 8900
rect 75288 8888 75316 8996
rect 75454 8984 75460 9036
rect 75512 9024 75518 9036
rect 79686 9024 79692 9036
rect 75512 8996 79692 9024
rect 75512 8984 75518 8996
rect 79686 8984 79692 8996
rect 79744 8984 79750 9036
rect 84470 9024 84476 9036
rect 79888 8996 84476 9024
rect 75362 8916 75368 8968
rect 75420 8956 75426 8968
rect 76285 8959 76343 8965
rect 76285 8956 76297 8959
rect 75420 8928 76297 8956
rect 75420 8916 75426 8928
rect 76285 8925 76297 8928
rect 76331 8925 76343 8959
rect 76285 8919 76343 8925
rect 76469 8959 76527 8965
rect 76469 8925 76481 8959
rect 76515 8956 76527 8959
rect 76650 8956 76656 8968
rect 76515 8928 76656 8956
rect 76515 8925 76527 8928
rect 76469 8919 76527 8925
rect 76650 8916 76656 8928
rect 76708 8956 76714 8968
rect 76929 8959 76987 8965
rect 76929 8956 76941 8959
rect 76708 8928 76941 8956
rect 76708 8916 76714 8928
rect 76929 8925 76941 8928
rect 76975 8925 76987 8959
rect 76929 8919 76987 8925
rect 79888 8888 79916 8996
rect 84470 8984 84476 8996
rect 84528 8984 84534 9036
rect 90836 9033 90864 9120
rect 94777 9095 94835 9101
rect 94777 9061 94789 9095
rect 94823 9061 94835 9095
rect 94777 9055 94835 9061
rect 90821 9027 90879 9033
rect 84672 8996 86540 9024
rect 80330 8916 80336 8968
rect 80388 8956 80394 8968
rect 84672 8956 84700 8996
rect 86402 8956 86408 8968
rect 80388 8928 84700 8956
rect 86363 8928 86408 8956
rect 80388 8916 80394 8928
rect 86402 8916 86408 8928
rect 86460 8916 86466 8968
rect 86512 8956 86540 8996
rect 90821 8993 90833 9027
rect 90867 8993 90879 9027
rect 92934 9024 92940 9036
rect 92895 8996 92940 9024
rect 90821 8987 90879 8993
rect 92934 8984 92940 8996
rect 92992 9024 92998 9036
rect 93397 9027 93455 9033
rect 93397 9024 93409 9027
rect 92992 8996 93409 9024
rect 92992 8984 92998 8996
rect 93397 8993 93409 8996
rect 93443 8993 93455 9027
rect 93397 8987 93455 8993
rect 89714 8956 89720 8968
rect 86512 8928 89720 8956
rect 89714 8916 89720 8928
rect 89772 8916 89778 8968
rect 90554 8959 90612 8965
rect 90554 8958 90566 8959
rect 90468 8930 90566 8958
rect 90468 8900 90496 8930
rect 90554 8925 90566 8930
rect 90600 8925 90612 8959
rect 90554 8919 90612 8925
rect 90910 8916 90916 8968
rect 90968 8956 90974 8968
rect 94792 8956 94820 9055
rect 95234 9052 95240 9104
rect 95292 9092 95298 9104
rect 96709 9095 96767 9101
rect 96709 9092 96721 9095
rect 95292 9064 96721 9092
rect 95292 9052 95298 9064
rect 96709 9061 96721 9064
rect 96755 9061 96767 9095
rect 96709 9055 96767 9061
rect 98086 9052 98092 9104
rect 98144 9092 98150 9104
rect 98549 9095 98607 9101
rect 98549 9092 98561 9095
rect 98144 9064 98561 9092
rect 98144 9052 98150 9064
rect 98549 9061 98561 9064
rect 98595 9092 98607 9095
rect 99374 9092 99380 9104
rect 98595 9064 99380 9092
rect 98595 9061 98607 9064
rect 98549 9055 98607 9061
rect 99374 9052 99380 9064
rect 99432 9092 99438 9104
rect 99742 9092 99748 9104
rect 99432 9064 99748 9092
rect 99432 9052 99438 9064
rect 99742 9052 99748 9064
rect 99800 9052 99806 9104
rect 95510 8984 95516 9036
rect 95568 9024 95574 9036
rect 96065 9027 96123 9033
rect 96065 9024 96077 9027
rect 95568 8996 96077 9024
rect 95568 8984 95574 8996
rect 96065 8993 96077 8996
rect 96111 8993 96123 9027
rect 96065 8987 96123 8993
rect 100757 9027 100815 9033
rect 100757 8993 100769 9027
rect 100803 9024 100815 9027
rect 101232 9024 101260 9120
rect 104434 9052 104440 9104
rect 104492 9092 104498 9104
rect 104897 9095 104955 9101
rect 104897 9092 104909 9095
rect 104492 9064 104909 9092
rect 104492 9052 104498 9064
rect 104897 9061 104909 9064
rect 104943 9061 104955 9095
rect 104897 9055 104955 9061
rect 107470 9052 107476 9104
rect 107528 9092 107534 9104
rect 120718 9092 120724 9104
rect 107528 9064 120724 9092
rect 107528 9052 107534 9064
rect 120718 9052 120724 9064
rect 120776 9052 120782 9104
rect 121914 9052 121920 9104
rect 121972 9092 121978 9104
rect 124214 9092 124220 9104
rect 121972 9064 124220 9092
rect 121972 9052 121978 9064
rect 124214 9052 124220 9064
rect 124272 9052 124278 9104
rect 126974 9092 126980 9104
rect 125566 9064 126836 9092
rect 126935 9064 126980 9092
rect 100803 8996 101260 9024
rect 100803 8993 100815 8996
rect 100757 8987 100815 8993
rect 90968 8928 94820 8956
rect 90968 8916 90974 8928
rect 71740 8860 75040 8888
rect 75288 8860 79916 8888
rect 71740 8848 71746 8860
rect 57330 8820 57336 8832
rect 56520 8792 57336 8820
rect 57330 8780 57336 8792
rect 57388 8780 57394 8832
rect 57514 8780 57520 8832
rect 57572 8820 57578 8832
rect 58250 8820 58256 8832
rect 57572 8792 58256 8820
rect 57572 8780 57578 8792
rect 58250 8780 58256 8792
rect 58308 8820 58314 8832
rect 59541 8823 59599 8829
rect 59541 8820 59553 8823
rect 58308 8792 59553 8820
rect 58308 8780 58314 8792
rect 59541 8789 59553 8792
rect 59587 8820 59599 8823
rect 59722 8820 59728 8832
rect 59587 8792 59728 8820
rect 59587 8789 59599 8792
rect 59541 8783 59599 8789
rect 59722 8780 59728 8792
rect 59780 8780 59786 8832
rect 61286 8780 61292 8832
rect 61344 8820 61350 8832
rect 61654 8820 61660 8832
rect 61344 8792 61660 8820
rect 61344 8780 61350 8792
rect 61654 8780 61660 8792
rect 61712 8780 61718 8832
rect 63497 8823 63555 8829
rect 63497 8789 63509 8823
rect 63543 8820 63555 8823
rect 63586 8820 63592 8832
rect 63543 8792 63592 8820
rect 63543 8789 63555 8792
rect 63497 8783 63555 8789
rect 63586 8780 63592 8792
rect 63644 8820 63650 8832
rect 65058 8820 65064 8832
rect 63644 8792 65064 8820
rect 63644 8780 63650 8792
rect 65058 8780 65064 8792
rect 65116 8780 65122 8832
rect 68281 8823 68339 8829
rect 68281 8789 68293 8823
rect 68327 8820 68339 8823
rect 68370 8820 68376 8832
rect 68327 8792 68376 8820
rect 68327 8789 68339 8792
rect 68281 8783 68339 8789
rect 68370 8780 68376 8792
rect 68428 8780 68434 8832
rect 73246 8780 73252 8832
rect 73304 8820 73310 8832
rect 74905 8823 74963 8829
rect 74905 8820 74917 8823
rect 73304 8792 74917 8820
rect 73304 8780 73310 8792
rect 74905 8789 74917 8792
rect 74951 8789 74963 8823
rect 75012 8820 75040 8860
rect 79962 8848 79968 8900
rect 80020 8888 80026 8900
rect 86494 8888 86500 8900
rect 80020 8860 86500 8888
rect 80020 8848 80026 8860
rect 86494 8848 86500 8860
rect 86552 8848 86558 8900
rect 86672 8891 86730 8897
rect 86672 8857 86684 8891
rect 86718 8888 86730 8891
rect 86718 8860 88380 8888
rect 86718 8857 86730 8860
rect 86672 8851 86730 8857
rect 88352 8832 88380 8860
rect 90450 8848 90456 8900
rect 90508 8848 90514 8900
rect 90726 8848 90732 8900
rect 90784 8888 90790 8900
rect 90784 8860 91692 8888
rect 90784 8848 90790 8860
rect 76006 8820 76012 8832
rect 75012 8792 76012 8820
rect 74905 8783 74963 8789
rect 76006 8780 76012 8792
rect 76064 8780 76070 8832
rect 76101 8823 76159 8829
rect 76101 8789 76113 8823
rect 76147 8820 76159 8823
rect 76282 8820 76288 8832
rect 76147 8792 76288 8820
rect 76147 8789 76159 8792
rect 76101 8783 76159 8789
rect 76282 8780 76288 8792
rect 76340 8780 76346 8832
rect 76374 8780 76380 8832
rect 76432 8820 76438 8832
rect 84010 8820 84016 8832
rect 76432 8792 84016 8820
rect 76432 8780 76438 8792
rect 84010 8780 84016 8792
rect 84068 8780 84074 8832
rect 84286 8780 84292 8832
rect 84344 8820 84350 8832
rect 87782 8820 87788 8832
rect 84344 8792 87788 8820
rect 84344 8780 84350 8792
rect 87782 8780 87788 8792
rect 87840 8780 87846 8832
rect 88334 8820 88340 8832
rect 88295 8792 88340 8820
rect 88334 8780 88340 8792
rect 88392 8780 88398 8832
rect 89438 8820 89444 8832
rect 89399 8792 89444 8820
rect 89438 8780 89444 8792
rect 89496 8780 89502 8832
rect 89622 8780 89628 8832
rect 89680 8820 89686 8832
rect 91557 8823 91615 8829
rect 91557 8820 91569 8823
rect 89680 8792 91569 8820
rect 89680 8780 89686 8792
rect 91557 8789 91569 8792
rect 91603 8789 91615 8823
rect 91664 8820 91692 8860
rect 92566 8848 92572 8900
rect 92624 8888 92630 8900
rect 93670 8897 93676 8900
rect 92670 8891 92728 8897
rect 92670 8888 92682 8891
rect 92624 8860 92682 8888
rect 92624 8848 92630 8860
rect 92670 8857 92682 8860
rect 92716 8857 92728 8891
rect 93664 8888 93676 8897
rect 93631 8860 93676 8888
rect 92670 8851 92728 8857
rect 93664 8851 93676 8860
rect 93670 8848 93676 8851
rect 93728 8848 93734 8900
rect 95418 8888 95424 8900
rect 93780 8860 95424 8888
rect 93780 8820 93808 8860
rect 95418 8848 95424 8860
rect 95476 8848 95482 8900
rect 96080 8888 96108 8987
rect 104618 8984 104624 9036
rect 104676 9024 104682 9036
rect 124769 9027 124827 9033
rect 104676 8996 123524 9024
rect 104676 8984 104682 8996
rect 96154 8916 96160 8968
rect 96212 8956 96218 8968
rect 96212 8928 97948 8956
rect 96212 8916 96218 8928
rect 97718 8888 97724 8900
rect 96080 8860 97724 8888
rect 97718 8848 97724 8860
rect 97776 8848 97782 8900
rect 97822 8891 97880 8897
rect 97822 8857 97834 8891
rect 97868 8857 97880 8891
rect 97920 8888 97948 8928
rect 97994 8916 98000 8968
rect 98052 8956 98058 8968
rect 98089 8959 98147 8965
rect 98089 8956 98101 8959
rect 98052 8928 98101 8956
rect 98052 8916 98058 8928
rect 98089 8925 98101 8928
rect 98135 8925 98147 8959
rect 98089 8919 98147 8925
rect 99466 8916 99472 8968
rect 99524 8956 99530 8968
rect 100490 8959 100548 8965
rect 100490 8956 100502 8959
rect 99524 8928 100502 8956
rect 99524 8916 99530 8928
rect 100490 8925 100502 8928
rect 100536 8925 100548 8959
rect 100490 8919 100548 8925
rect 107194 8916 107200 8968
rect 107252 8956 107258 8968
rect 107381 8959 107439 8965
rect 107381 8956 107393 8959
rect 107252 8928 107393 8956
rect 107252 8916 107258 8928
rect 107381 8925 107393 8928
rect 107427 8925 107439 8959
rect 107562 8956 107568 8968
rect 107523 8928 107568 8956
rect 107381 8919 107439 8925
rect 104253 8891 104311 8897
rect 104253 8888 104265 8891
rect 97920 8860 104265 8888
rect 97822 8851 97880 8857
rect 104253 8857 104265 8860
rect 104299 8888 104311 8891
rect 104618 8888 104624 8900
rect 104299 8860 104624 8888
rect 104299 8857 104311 8860
rect 104253 8851 104311 8857
rect 91664 8792 93808 8820
rect 91557 8783 91615 8789
rect 95050 8780 95056 8832
rect 95108 8820 95114 8832
rect 97626 8820 97632 8832
rect 95108 8792 97632 8820
rect 95108 8780 95114 8792
rect 97626 8780 97632 8792
rect 97684 8780 97690 8832
rect 97828 8820 97856 8851
rect 104618 8848 104624 8860
rect 104676 8848 104682 8900
rect 107396 8888 107424 8919
rect 107562 8916 107568 8928
rect 107620 8916 107626 8968
rect 107749 8959 107807 8965
rect 107749 8925 107761 8959
rect 107795 8956 107807 8959
rect 108393 8959 108451 8965
rect 108393 8956 108405 8959
rect 107795 8928 108405 8956
rect 107795 8925 107807 8928
rect 107749 8919 107807 8925
rect 108393 8925 108405 8928
rect 108439 8925 108451 8959
rect 108393 8919 108451 8925
rect 111061 8959 111119 8965
rect 111061 8925 111073 8959
rect 111107 8956 111119 8959
rect 111334 8956 111340 8968
rect 111107 8928 111340 8956
rect 111107 8925 111119 8928
rect 111061 8919 111119 8925
rect 111334 8916 111340 8928
rect 111392 8916 111398 8968
rect 112346 8956 112352 8968
rect 112307 8928 112352 8956
rect 112346 8916 112352 8928
rect 112404 8916 112410 8968
rect 118142 8956 118148 8968
rect 118103 8928 118148 8956
rect 118142 8916 118148 8928
rect 118200 8916 118206 8968
rect 119614 8916 119620 8968
rect 119672 8956 119678 8968
rect 120902 8956 120908 8968
rect 119672 8928 119717 8956
rect 120184 8928 120908 8956
rect 119672 8916 119678 8928
rect 107930 8888 107936 8900
rect 107396 8860 107936 8888
rect 107930 8848 107936 8860
rect 107988 8888 107994 8900
rect 108942 8888 108948 8900
rect 107988 8860 108948 8888
rect 107988 8848 107994 8860
rect 108942 8848 108948 8860
rect 109000 8848 109006 8900
rect 109218 8848 109224 8900
rect 109276 8888 109282 8900
rect 112364 8888 112392 8916
rect 116765 8891 116823 8897
rect 109276 8860 112208 8888
rect 112364 8860 116072 8888
rect 109276 8848 109282 8860
rect 98178 8820 98184 8832
rect 97828 8792 98184 8820
rect 98178 8780 98184 8792
rect 98236 8780 98242 8832
rect 99374 8780 99380 8832
rect 99432 8820 99438 8832
rect 108206 8820 108212 8832
rect 99432 8792 99477 8820
rect 108167 8792 108212 8820
rect 99432 8780 99438 8792
rect 108206 8780 108212 8792
rect 108264 8780 108270 8832
rect 110782 8780 110788 8832
rect 110840 8820 110846 8832
rect 110877 8823 110935 8829
rect 110877 8820 110889 8823
rect 110840 8792 110889 8820
rect 110840 8780 110846 8792
rect 110877 8789 110889 8792
rect 110923 8789 110935 8823
rect 112180 8820 112208 8860
rect 112533 8823 112591 8829
rect 112533 8820 112545 8823
rect 112180 8792 112545 8820
rect 110877 8783 110935 8789
rect 112533 8789 112545 8792
rect 112579 8820 112591 8823
rect 113085 8823 113143 8829
rect 113085 8820 113097 8823
rect 112579 8792 113097 8820
rect 112579 8789 112591 8792
rect 112533 8783 112591 8789
rect 113085 8789 113097 8792
rect 113131 8820 113143 8823
rect 113266 8820 113272 8832
rect 113131 8792 113272 8820
rect 113131 8789 113143 8792
rect 113085 8783 113143 8789
rect 113266 8780 113272 8792
rect 113324 8820 113330 8832
rect 115842 8820 115848 8832
rect 113324 8792 115848 8820
rect 113324 8780 113330 8792
rect 115842 8780 115848 8792
rect 115900 8820 115906 8832
rect 115937 8823 115995 8829
rect 115937 8820 115949 8823
rect 115900 8792 115949 8820
rect 115900 8780 115906 8792
rect 115937 8789 115949 8792
rect 115983 8789 115995 8823
rect 116044 8820 116072 8860
rect 116765 8857 116777 8891
rect 116811 8888 116823 8891
rect 117222 8888 117228 8900
rect 116811 8860 117228 8888
rect 116811 8857 116823 8860
rect 116765 8851 116823 8857
rect 117222 8848 117228 8860
rect 117280 8848 117286 8900
rect 118418 8848 118424 8900
rect 118476 8888 118482 8900
rect 119433 8891 119491 8897
rect 119433 8888 119445 8891
rect 118476 8860 119445 8888
rect 118476 8848 118482 8860
rect 119433 8857 119445 8860
rect 119479 8857 119491 8891
rect 119433 8851 119491 8857
rect 116946 8820 116952 8832
rect 116044 8792 116952 8820
rect 115937 8783 115995 8789
rect 116946 8780 116952 8792
rect 117004 8780 117010 8832
rect 117130 8780 117136 8832
rect 117188 8820 117194 8832
rect 117317 8823 117375 8829
rect 117317 8820 117329 8823
rect 117188 8792 117329 8820
rect 117188 8780 117194 8792
rect 117317 8789 117329 8792
rect 117363 8789 117375 8823
rect 117317 8783 117375 8789
rect 118697 8823 118755 8829
rect 118697 8789 118709 8823
rect 118743 8820 118755 8823
rect 118970 8820 118976 8832
rect 118743 8792 118976 8820
rect 118743 8789 118755 8792
rect 118697 8783 118755 8789
rect 118970 8780 118976 8792
rect 119028 8780 119034 8832
rect 119154 8780 119160 8832
rect 119212 8820 119218 8832
rect 120184 8829 120212 8928
rect 120902 8916 120908 8928
rect 120960 8916 120966 8968
rect 121822 8916 121828 8968
rect 121880 8956 121886 8968
rect 122653 8959 122711 8965
rect 122653 8956 122665 8959
rect 121880 8928 122665 8956
rect 121880 8916 121886 8928
rect 122653 8925 122665 8928
rect 122699 8925 122711 8959
rect 122653 8919 122711 8925
rect 122837 8959 122895 8965
rect 122837 8925 122849 8959
rect 122883 8956 122895 8959
rect 122883 8928 123432 8956
rect 122883 8925 122895 8928
rect 122837 8919 122895 8925
rect 120442 8848 120448 8900
rect 120500 8888 120506 8900
rect 120500 8860 121684 8888
rect 120500 8848 120506 8860
rect 120169 8823 120227 8829
rect 120169 8820 120181 8823
rect 119212 8792 120181 8820
rect 119212 8780 119218 8792
rect 120169 8789 120181 8792
rect 120215 8789 120227 8823
rect 120169 8783 120227 8789
rect 120258 8780 120264 8832
rect 120316 8820 120322 8832
rect 120721 8823 120779 8829
rect 120721 8820 120733 8823
rect 120316 8792 120733 8820
rect 120316 8780 120322 8792
rect 120721 8789 120733 8792
rect 120767 8789 120779 8823
rect 121362 8820 121368 8832
rect 121323 8792 121368 8820
rect 120721 8783 120779 8789
rect 121362 8780 121368 8792
rect 121420 8780 121426 8832
rect 121656 8820 121684 8860
rect 122374 8820 122380 8832
rect 121656 8792 122380 8820
rect 122374 8780 122380 8792
rect 122432 8780 122438 8832
rect 122466 8780 122472 8832
rect 122524 8820 122530 8832
rect 123404 8829 123432 8928
rect 123496 8888 123524 8996
rect 124769 8993 124781 9027
rect 124815 9024 124827 9027
rect 125566 9024 125594 9064
rect 124815 8996 125594 9024
rect 124815 8993 124827 8996
rect 124769 8987 124827 8993
rect 126606 8984 126612 9036
rect 126664 9024 126670 9036
rect 126808 9024 126836 9064
rect 126974 9052 126980 9064
rect 127032 9052 127038 9104
rect 129090 9092 129096 9104
rect 127452 9064 129096 9092
rect 127452 9024 127480 9064
rect 129090 9052 129096 9064
rect 129148 9052 129154 9104
rect 126664 8996 126709 9024
rect 126808 8996 127480 9024
rect 126664 8984 126670 8996
rect 127526 8984 127532 9036
rect 127584 9024 127590 9036
rect 129200 9033 129228 9132
rect 130930 9120 130936 9132
rect 130988 9120 130994 9172
rect 131022 9120 131028 9172
rect 131080 9160 131086 9172
rect 131669 9163 131727 9169
rect 131080 9132 131620 9160
rect 131080 9120 131086 9132
rect 130565 9095 130623 9101
rect 130565 9061 130577 9095
rect 130611 9092 130623 9095
rect 130838 9092 130844 9104
rect 130611 9064 130844 9092
rect 130611 9061 130623 9064
rect 130565 9055 130623 9061
rect 130838 9052 130844 9064
rect 130896 9052 130902 9104
rect 131114 9092 131120 9104
rect 131075 9064 131120 9092
rect 131114 9052 131120 9064
rect 131172 9052 131178 9104
rect 131592 9092 131620 9132
rect 131669 9129 131681 9163
rect 131715 9160 131727 9163
rect 131942 9160 131948 9172
rect 131715 9132 131948 9160
rect 131715 9129 131727 9132
rect 131669 9123 131727 9129
rect 131942 9120 131948 9132
rect 132000 9120 132006 9172
rect 134794 9160 134800 9172
rect 132420 9132 134800 9160
rect 132420 9092 132448 9132
rect 134794 9120 134800 9132
rect 134852 9120 134858 9172
rect 135070 9120 135076 9172
rect 135128 9160 135134 9172
rect 136450 9160 136456 9172
rect 135128 9132 136456 9160
rect 135128 9120 135134 9132
rect 136450 9120 136456 9132
rect 136508 9120 136514 9172
rect 136542 9120 136548 9172
rect 136600 9160 136606 9172
rect 137830 9160 137836 9172
rect 136600 9132 137836 9160
rect 136600 9120 136606 9132
rect 137830 9120 137836 9132
rect 137888 9160 137894 9172
rect 137888 9132 138060 9160
rect 137888 9120 137894 9132
rect 131592 9064 132448 9092
rect 132494 9052 132500 9104
rect 132552 9092 132558 9104
rect 137922 9092 137928 9104
rect 132552 9064 137928 9092
rect 132552 9052 132558 9064
rect 137922 9052 137928 9064
rect 137980 9052 137986 9104
rect 138032 9092 138060 9132
rect 138198 9120 138204 9172
rect 138256 9160 138262 9172
rect 145742 9160 145748 9172
rect 138256 9132 145748 9160
rect 138256 9120 138262 9132
rect 145742 9120 145748 9132
rect 145800 9120 145806 9172
rect 146018 9120 146024 9172
rect 146076 9160 146082 9172
rect 146076 9132 148732 9160
rect 146076 9120 146082 9132
rect 138109 9095 138167 9101
rect 138109 9092 138121 9095
rect 138032 9064 138121 9092
rect 138109 9061 138121 9064
rect 138155 9061 138167 9095
rect 138658 9092 138664 9104
rect 138619 9064 138664 9092
rect 138109 9055 138167 9061
rect 138658 9052 138664 9064
rect 138716 9052 138722 9104
rect 139305 9095 139363 9101
rect 139305 9061 139317 9095
rect 139351 9092 139363 9095
rect 139486 9092 139492 9104
rect 139351 9064 139492 9092
rect 139351 9061 139363 9064
rect 139305 9055 139363 9061
rect 139486 9052 139492 9064
rect 139544 9052 139550 9104
rect 139762 9052 139768 9104
rect 139820 9092 139826 9104
rect 139857 9095 139915 9101
rect 139857 9092 139869 9095
rect 139820 9064 139869 9092
rect 139820 9052 139826 9064
rect 139857 9061 139869 9064
rect 139903 9092 139915 9095
rect 140590 9092 140596 9104
rect 139903 9064 140596 9092
rect 139903 9061 139915 9064
rect 139857 9055 139915 9061
rect 140590 9052 140596 9064
rect 140648 9052 140654 9104
rect 140682 9052 140688 9104
rect 140740 9092 140746 9104
rect 143442 9092 143448 9104
rect 140740 9064 143448 9092
rect 140740 9052 140746 9064
rect 143442 9052 143448 9064
rect 143500 9052 143506 9104
rect 144638 9052 144644 9104
rect 144696 9092 144702 9104
rect 144917 9095 144975 9101
rect 144917 9092 144929 9095
rect 144696 9064 144929 9092
rect 144696 9052 144702 9064
rect 144917 9061 144929 9064
rect 144963 9092 144975 9095
rect 145098 9092 145104 9104
rect 144963 9064 145104 9092
rect 144963 9061 144975 9064
rect 144917 9055 144975 9061
rect 145098 9052 145104 9064
rect 145156 9052 145162 9104
rect 145466 9052 145472 9104
rect 145524 9092 145530 9104
rect 145653 9095 145711 9101
rect 145653 9092 145665 9095
rect 145524 9064 145665 9092
rect 145524 9052 145530 9064
rect 145653 9061 145665 9064
rect 145699 9061 145711 9095
rect 145653 9055 145711 9061
rect 147214 9052 147220 9104
rect 147272 9092 147278 9104
rect 148594 9092 148600 9104
rect 147272 9064 148600 9092
rect 147272 9052 147278 9064
rect 148594 9052 148600 9064
rect 148652 9052 148658 9104
rect 129185 9027 129243 9033
rect 127584 8996 128768 9024
rect 127584 8984 127590 8996
rect 123754 8916 123760 8968
rect 123812 8956 123818 8968
rect 126793 8959 126851 8965
rect 126793 8956 126805 8959
rect 123812 8950 126560 8956
rect 126716 8950 126805 8956
rect 123812 8928 126805 8950
rect 123812 8916 123818 8928
rect 126532 8922 126744 8928
rect 126793 8925 126805 8928
rect 126839 8956 126851 8959
rect 127621 8959 127679 8965
rect 127621 8956 127633 8959
rect 126839 8928 127633 8956
rect 126839 8925 126851 8928
rect 126793 8919 126851 8925
rect 127621 8925 127633 8928
rect 127667 8925 127679 8959
rect 127621 8919 127679 8925
rect 128740 8897 128768 8996
rect 129185 8993 129197 9027
rect 129231 8993 129243 9027
rect 137370 9024 137376 9036
rect 129185 8987 129243 8993
rect 131960 8996 137376 9024
rect 128814 8916 128820 8968
rect 128872 8956 128878 8968
rect 131666 8956 131672 8968
rect 128872 8928 131672 8956
rect 128872 8916 128878 8928
rect 131666 8916 131672 8928
rect 131724 8916 131730 8968
rect 128725 8891 128783 8897
rect 123496 8860 126376 8888
rect 123389 8823 123447 8829
rect 122524 8792 122569 8820
rect 122524 8780 122530 8792
rect 123389 8789 123401 8823
rect 123435 8820 123447 8823
rect 123846 8820 123852 8832
rect 123435 8792 123852 8820
rect 123435 8789 123447 8792
rect 123389 8783 123447 8789
rect 123846 8780 123852 8792
rect 123904 8780 123910 8832
rect 124217 8823 124275 8829
rect 124217 8789 124229 8823
rect 124263 8820 124275 8823
rect 124398 8820 124404 8832
rect 124263 8792 124404 8820
rect 124263 8789 124275 8792
rect 124217 8783 124275 8789
rect 124398 8780 124404 8792
rect 124456 8820 124462 8832
rect 125229 8823 125287 8829
rect 125229 8820 125241 8823
rect 124456 8792 125241 8820
rect 124456 8780 124462 8792
rect 125229 8789 125241 8792
rect 125275 8820 125287 8823
rect 125410 8820 125416 8832
rect 125275 8792 125416 8820
rect 125275 8789 125287 8792
rect 125229 8783 125287 8789
rect 125410 8780 125416 8792
rect 125468 8780 125474 8832
rect 125686 8780 125692 8832
rect 125744 8820 125750 8832
rect 125873 8823 125931 8829
rect 125873 8820 125885 8823
rect 125744 8792 125885 8820
rect 125744 8780 125750 8792
rect 125873 8789 125885 8792
rect 125919 8820 125931 8823
rect 126238 8820 126244 8832
rect 125919 8792 126244 8820
rect 125919 8789 125931 8792
rect 125873 8783 125931 8789
rect 126238 8780 126244 8792
rect 126296 8780 126302 8832
rect 126348 8820 126376 8860
rect 126716 8860 128676 8888
rect 126716 8820 126744 8860
rect 126348 8792 126744 8820
rect 127710 8780 127716 8832
rect 127768 8820 127774 8832
rect 128538 8820 128544 8832
rect 127768 8792 128544 8820
rect 127768 8780 127774 8792
rect 128538 8780 128544 8792
rect 128596 8780 128602 8832
rect 128648 8820 128676 8860
rect 128725 8857 128737 8891
rect 128771 8888 128783 8891
rect 129430 8891 129488 8897
rect 129430 8888 129442 8891
rect 128771 8860 129442 8888
rect 128771 8857 128783 8860
rect 128725 8851 128783 8857
rect 129430 8857 129442 8860
rect 129476 8857 129488 8891
rect 129430 8851 129488 8857
rect 129550 8848 129556 8900
rect 129608 8888 129614 8900
rect 130286 8888 130292 8900
rect 129608 8860 130292 8888
rect 129608 8848 129614 8860
rect 130286 8848 130292 8860
rect 130344 8848 130350 8900
rect 131960 8888 131988 8996
rect 137370 8984 137376 8996
rect 137428 8984 137434 9036
rect 137554 8984 137560 9036
rect 137612 9024 137618 9036
rect 139578 9024 139584 9036
rect 137612 8996 139584 9024
rect 137612 8984 137618 8996
rect 139578 8984 139584 8996
rect 139636 8984 139642 9036
rect 145834 9024 145840 9036
rect 140332 8996 143488 9024
rect 132957 8959 133015 8965
rect 132957 8956 132969 8959
rect 132144 8928 132969 8956
rect 132144 8900 132172 8928
rect 132957 8925 132969 8928
rect 133003 8925 133015 8959
rect 132957 8919 133015 8925
rect 133141 8959 133199 8965
rect 133141 8925 133153 8959
rect 133187 8956 133199 8959
rect 133506 8956 133512 8968
rect 133187 8928 133512 8956
rect 133187 8925 133199 8928
rect 133141 8919 133199 8925
rect 133506 8916 133512 8928
rect 133564 8916 133570 8968
rect 133690 8916 133696 8968
rect 133748 8956 133754 8968
rect 135070 8956 135076 8968
rect 133748 8928 135076 8956
rect 133748 8916 133754 8928
rect 135070 8916 135076 8928
rect 135128 8916 135134 8968
rect 135254 8916 135260 8968
rect 135312 8956 135318 8968
rect 135625 8959 135683 8965
rect 135625 8956 135637 8959
rect 135312 8928 135637 8956
rect 135312 8916 135318 8928
rect 135625 8925 135637 8928
rect 135671 8956 135683 8959
rect 135990 8956 135996 8968
rect 135671 8928 135996 8956
rect 135671 8925 135683 8928
rect 135625 8919 135683 8925
rect 135990 8916 135996 8928
rect 136048 8916 136054 8968
rect 136450 8916 136456 8968
rect 136508 8956 136514 8968
rect 137925 8959 137983 8965
rect 137925 8956 137937 8959
rect 136508 8928 137937 8956
rect 136508 8916 136514 8928
rect 137925 8925 137937 8928
rect 137971 8956 137983 8959
rect 138658 8956 138664 8968
rect 137971 8928 138664 8956
rect 137971 8925 137983 8928
rect 137925 8919 137983 8925
rect 138658 8916 138664 8928
rect 138716 8916 138722 8968
rect 140332 8965 140360 8996
rect 140317 8959 140375 8965
rect 140317 8925 140329 8959
rect 140363 8925 140375 8959
rect 140317 8919 140375 8925
rect 140958 8916 140964 8968
rect 141016 8956 141022 8968
rect 141016 8928 141061 8956
rect 141016 8916 141022 8928
rect 141510 8916 141516 8968
rect 141568 8956 141574 8968
rect 141697 8959 141755 8965
rect 141697 8956 141709 8959
rect 141568 8928 141709 8956
rect 141568 8916 141574 8928
rect 141697 8925 141709 8928
rect 141743 8925 141755 8959
rect 141970 8956 141976 8968
rect 141931 8928 141976 8956
rect 141697 8919 141755 8925
rect 141970 8916 141976 8928
rect 142028 8916 142034 8968
rect 143460 8956 143488 8996
rect 144380 8996 145840 9024
rect 143626 8956 143632 8968
rect 143460 8928 143632 8956
rect 143626 8916 143632 8928
rect 143684 8916 143690 8968
rect 144201 8959 144259 8965
rect 144201 8925 144213 8959
rect 144247 8956 144259 8959
rect 144380 8956 144408 8996
rect 145834 8984 145840 8996
rect 145892 8984 145898 9036
rect 147033 9027 147091 9033
rect 147033 8993 147045 9027
rect 147079 9024 147091 9027
rect 147122 9024 147128 9036
rect 147079 8996 147128 9024
rect 147079 8993 147091 8996
rect 147033 8987 147091 8993
rect 147122 8984 147128 8996
rect 147180 9024 147186 9036
rect 147490 9024 147496 9036
rect 147180 8996 147496 9024
rect 147180 8984 147186 8996
rect 147490 8984 147496 8996
rect 147548 8984 147554 9036
rect 148226 9024 148232 9036
rect 147600 8996 148232 9024
rect 144247 8928 144408 8956
rect 144457 8959 144515 8965
rect 144247 8925 144259 8928
rect 144201 8919 144259 8925
rect 144457 8925 144469 8959
rect 144503 8956 144515 8959
rect 144638 8956 144644 8968
rect 144503 8928 144644 8956
rect 144503 8925 144515 8928
rect 144457 8919 144515 8925
rect 144638 8916 144644 8928
rect 144696 8956 144702 8968
rect 144822 8956 144828 8968
rect 144696 8928 144828 8956
rect 144696 8916 144702 8928
rect 144822 8916 144828 8928
rect 144880 8916 144886 8968
rect 145006 8916 145012 8968
rect 145064 8956 145070 8968
rect 147398 8956 147404 8968
rect 145064 8928 147404 8956
rect 145064 8916 145070 8928
rect 147398 8916 147404 8928
rect 147456 8916 147462 8968
rect 147600 8956 147628 8996
rect 148226 8984 148232 8996
rect 148284 8984 148290 9036
rect 147508 8928 147628 8956
rect 132126 8888 132132 8900
rect 130764 8860 131988 8888
rect 132087 8860 132132 8888
rect 130764 8820 130792 8860
rect 132126 8848 132132 8860
rect 132184 8848 132190 8900
rect 137370 8888 137376 8900
rect 132236 8860 137376 8888
rect 128648 8792 130792 8820
rect 130838 8780 130844 8832
rect 130896 8820 130902 8832
rect 132236 8820 132264 8860
rect 137370 8848 137376 8860
rect 137428 8848 137434 8900
rect 140516 8860 141280 8888
rect 130896 8792 132264 8820
rect 132773 8823 132831 8829
rect 130896 8780 130902 8792
rect 132773 8789 132785 8823
rect 132819 8820 132831 8823
rect 132862 8820 132868 8832
rect 132819 8792 132868 8820
rect 132819 8789 132831 8792
rect 132773 8783 132831 8789
rect 132862 8780 132868 8792
rect 132920 8780 132926 8832
rect 133506 8780 133512 8832
rect 133564 8820 133570 8832
rect 133601 8823 133659 8829
rect 133601 8820 133613 8823
rect 133564 8792 133613 8820
rect 133564 8780 133570 8792
rect 133601 8789 133613 8792
rect 133647 8789 133659 8823
rect 133601 8783 133659 8789
rect 133782 8780 133788 8832
rect 133840 8820 133846 8832
rect 134153 8823 134211 8829
rect 134153 8820 134165 8823
rect 133840 8792 134165 8820
rect 133840 8780 133846 8792
rect 134153 8789 134165 8792
rect 134199 8789 134211 8823
rect 134153 8783 134211 8789
rect 135165 8823 135223 8829
rect 135165 8789 135177 8823
rect 135211 8820 135223 8823
rect 135254 8820 135260 8832
rect 135211 8792 135260 8820
rect 135211 8789 135223 8792
rect 135165 8783 135223 8789
rect 135254 8780 135260 8792
rect 135312 8780 135318 8832
rect 135530 8780 135536 8832
rect 135588 8820 135594 8832
rect 135809 8823 135867 8829
rect 135809 8820 135821 8823
rect 135588 8792 135821 8820
rect 135588 8780 135594 8792
rect 135809 8789 135821 8792
rect 135855 8789 135867 8823
rect 135809 8783 135867 8789
rect 135990 8780 135996 8832
rect 136048 8820 136054 8832
rect 136450 8820 136456 8832
rect 136048 8792 136456 8820
rect 136048 8780 136054 8792
rect 136450 8780 136456 8792
rect 136508 8780 136514 8832
rect 136910 8780 136916 8832
rect 136968 8820 136974 8832
rect 137281 8823 137339 8829
rect 137281 8820 137293 8823
rect 136968 8792 137293 8820
rect 136968 8780 136974 8792
rect 137281 8789 137293 8792
rect 137327 8789 137339 8823
rect 137281 8783 137339 8789
rect 137462 8780 137468 8832
rect 137520 8820 137526 8832
rect 139670 8820 139676 8832
rect 137520 8792 139676 8820
rect 137520 8780 137526 8792
rect 139670 8780 139676 8792
rect 139728 8780 139734 8832
rect 140516 8829 140544 8860
rect 140501 8823 140559 8829
rect 140501 8789 140513 8823
rect 140547 8789 140559 8823
rect 140501 8783 140559 8789
rect 140590 8780 140596 8832
rect 140648 8820 140654 8832
rect 141145 8823 141203 8829
rect 141145 8820 141157 8823
rect 140648 8792 141157 8820
rect 140648 8780 140654 8792
rect 141145 8789 141157 8792
rect 141191 8789 141203 8823
rect 141252 8820 141280 8860
rect 141326 8848 141332 8900
rect 141384 8888 141390 8900
rect 146788 8891 146846 8897
rect 141384 8860 146708 8888
rect 141384 8848 141390 8860
rect 142890 8820 142896 8832
rect 141252 8792 142896 8820
rect 141145 8783 141203 8789
rect 142890 8780 142896 8792
rect 142948 8780 142954 8832
rect 143074 8820 143080 8832
rect 143035 8792 143080 8820
rect 143074 8780 143080 8792
rect 143132 8780 143138 8832
rect 144546 8780 144552 8832
rect 144604 8820 144610 8832
rect 145926 8820 145932 8832
rect 144604 8792 145932 8820
rect 144604 8780 144610 8792
rect 145926 8780 145932 8792
rect 145984 8780 145990 8832
rect 146680 8820 146708 8860
rect 146788 8857 146800 8891
rect 146834 8888 146846 8891
rect 147122 8888 147128 8900
rect 146834 8860 147128 8888
rect 146834 8857 146846 8860
rect 146788 8851 146846 8857
rect 147122 8848 147128 8860
rect 147180 8848 147186 8900
rect 147508 8888 147536 8928
rect 147416 8860 147536 8888
rect 147416 8820 147444 8860
rect 146680 8792 147444 8820
rect 147490 8780 147496 8832
rect 147548 8820 147554 8832
rect 148318 8820 148324 8832
rect 147548 8792 148324 8820
rect 147548 8780 147554 8792
rect 148318 8780 148324 8792
rect 148376 8780 148382 8832
rect 148704 8820 148732 9132
rect 148778 9120 148784 9172
rect 148836 9160 148842 9172
rect 148836 9132 148881 9160
rect 148980 9132 153194 9160
rect 148836 9120 148842 9132
rect 148870 9052 148876 9104
rect 148928 9092 148934 9104
rect 148980 9092 149008 9132
rect 148928 9064 149008 9092
rect 148928 9052 148934 9064
rect 150434 9052 150440 9104
rect 150492 9092 150498 9104
rect 151814 9092 151820 9104
rect 150492 9064 151820 9092
rect 150492 9052 150498 9064
rect 151814 9052 151820 9064
rect 151872 9092 151878 9104
rect 152826 9092 152832 9104
rect 151872 9064 152832 9092
rect 151872 9052 151878 9064
rect 152826 9052 152832 9064
rect 152884 9052 152890 9104
rect 153166 9092 153194 9132
rect 153562 9120 153568 9172
rect 153620 9160 153626 9172
rect 154666 9160 154672 9172
rect 153620 9132 154672 9160
rect 153620 9120 153626 9132
rect 154666 9120 154672 9132
rect 154724 9120 154730 9172
rect 155405 9163 155463 9169
rect 155405 9129 155417 9163
rect 155451 9160 155463 9163
rect 157794 9160 157800 9172
rect 155451 9132 157800 9160
rect 155451 9129 155463 9132
rect 155405 9123 155463 9129
rect 157794 9120 157800 9132
rect 157852 9120 157858 9172
rect 153654 9092 153660 9104
rect 153166 9064 153660 9092
rect 153654 9052 153660 9064
rect 153712 9052 153718 9104
rect 153749 9095 153807 9101
rect 153749 9061 153761 9095
rect 153795 9092 153807 9095
rect 154758 9092 154764 9104
rect 153795 9064 154764 9092
rect 153795 9061 153807 9064
rect 153749 9055 153807 9061
rect 154758 9052 154764 9064
rect 154816 9052 154822 9104
rect 156874 9052 156880 9104
rect 156932 9092 156938 9104
rect 157521 9095 157579 9101
rect 157521 9092 157533 9095
rect 156932 9064 157533 9092
rect 156932 9052 156938 9064
rect 157521 9061 157533 9064
rect 157567 9061 157579 9095
rect 157521 9055 157579 9061
rect 150621 9027 150679 9033
rect 150621 8993 150633 9027
rect 150667 9024 150679 9027
rect 150667 8996 150940 9024
rect 150667 8993 150679 8996
rect 150621 8987 150679 8993
rect 149606 8916 149612 8968
rect 149664 8956 149670 8968
rect 150161 8959 150219 8965
rect 150161 8956 150173 8959
rect 149664 8928 150173 8956
rect 149664 8916 149670 8928
rect 150161 8925 150173 8928
rect 150207 8925 150219 8959
rect 150161 8919 150219 8925
rect 150250 8916 150256 8968
rect 150308 8956 150314 8968
rect 150805 8959 150863 8965
rect 150805 8956 150817 8959
rect 150308 8928 150817 8956
rect 150308 8916 150314 8928
rect 150805 8925 150817 8928
rect 150851 8925 150863 8959
rect 150912 8956 150940 8996
rect 151998 8984 152004 9036
rect 152056 9024 152062 9036
rect 152056 8996 153608 9024
rect 152056 8984 152062 8996
rect 151541 8959 151599 8965
rect 151541 8956 151553 8959
rect 150912 8928 151553 8956
rect 150805 8919 150863 8925
rect 151541 8925 151553 8928
rect 151587 8925 151599 8959
rect 151541 8919 151599 8925
rect 149916 8891 149974 8897
rect 149916 8857 149928 8891
rect 149962 8888 149974 8891
rect 150894 8888 150900 8900
rect 149962 8860 150900 8888
rect 149962 8857 149974 8860
rect 149916 8851 149974 8857
rect 150894 8848 150900 8860
rect 150952 8848 150958 8900
rect 150526 8820 150532 8832
rect 148704 8792 150532 8820
rect 150526 8780 150532 8792
rect 150584 8780 150590 8832
rect 150986 8820 150992 8832
rect 150947 8792 150992 8820
rect 150986 8780 150992 8792
rect 151044 8780 151050 8832
rect 151565 8820 151593 8919
rect 151630 8916 151636 8968
rect 151688 8956 151694 8968
rect 151817 8959 151875 8965
rect 151688 8928 151733 8956
rect 151688 8916 151694 8928
rect 151817 8925 151829 8959
rect 151863 8956 151875 8959
rect 152090 8956 152096 8968
rect 151863 8928 152096 8956
rect 151863 8925 151875 8928
rect 151817 8919 151875 8925
rect 152090 8916 152096 8928
rect 152148 8916 152154 8968
rect 152458 8956 152464 8968
rect 152419 8928 152464 8956
rect 152458 8916 152464 8928
rect 152516 8916 152522 8968
rect 152550 8916 152556 8968
rect 152608 8956 152614 8968
rect 153470 8956 153476 8968
rect 152608 8928 152653 8956
rect 153383 8928 153476 8956
rect 152608 8916 152614 8928
rect 153470 8916 153476 8928
rect 153528 8916 153534 8968
rect 153580 8965 153608 8996
rect 155034 8984 155040 9036
rect 155092 9024 155098 9036
rect 155954 9024 155960 9036
rect 155092 8996 155960 9024
rect 155092 8984 155098 8996
rect 153565 8959 153623 8965
rect 153565 8925 153577 8959
rect 153611 8925 153623 8959
rect 153565 8919 153623 8925
rect 153930 8916 153936 8968
rect 153988 8956 153994 8968
rect 154206 8956 154212 8968
rect 153988 8928 154212 8956
rect 153988 8916 153994 8928
rect 154206 8916 154212 8928
rect 154264 8916 154270 8968
rect 155144 8965 155172 8996
rect 155954 8984 155960 8996
rect 156012 8984 156018 9036
rect 154393 8959 154451 8965
rect 154393 8925 154405 8959
rect 154439 8925 154451 8959
rect 154393 8919 154451 8925
rect 155129 8959 155187 8965
rect 155129 8925 155141 8959
rect 155175 8925 155187 8959
rect 155129 8919 155187 8925
rect 151722 8848 151728 8900
rect 151780 8888 151786 8900
rect 152277 8891 152335 8897
rect 152277 8888 152289 8891
rect 151780 8860 152289 8888
rect 151780 8848 151786 8860
rect 152277 8857 152289 8860
rect 152323 8857 152335 8891
rect 153488 8888 153516 8916
rect 153654 8888 153660 8900
rect 152277 8851 152335 8857
rect 152384 8860 153660 8888
rect 152384 8820 152412 8860
rect 153654 8848 153660 8860
rect 153712 8848 153718 8900
rect 151565 8792 152412 8820
rect 152826 8780 152832 8832
rect 152884 8820 152890 8832
rect 154408 8820 154436 8919
rect 155218 8916 155224 8968
rect 155276 8956 155282 8968
rect 156046 8956 156052 8968
rect 155276 8928 155321 8956
rect 156007 8928 156052 8956
rect 155276 8916 155282 8928
rect 156046 8916 156052 8928
rect 156104 8916 156110 8968
rect 156138 8916 156144 8968
rect 156196 8956 156202 8968
rect 156196 8928 156241 8956
rect 156196 8916 156202 8928
rect 156322 8916 156328 8968
rect 156380 8956 156386 8968
rect 156693 8959 156751 8965
rect 156693 8956 156705 8959
rect 156380 8928 156705 8956
rect 156380 8916 156386 8928
rect 156693 8925 156705 8928
rect 156739 8925 156751 8959
rect 156693 8919 156751 8925
rect 156782 8916 156788 8968
rect 156840 8956 156846 8968
rect 156877 8959 156935 8965
rect 156877 8956 156889 8959
rect 156840 8928 156889 8956
rect 156840 8916 156846 8928
rect 156877 8925 156889 8928
rect 156923 8925 156935 8959
rect 157702 8956 157708 8968
rect 157663 8928 157708 8956
rect 156877 8919 156935 8925
rect 157702 8916 157708 8928
rect 157760 8916 157766 8968
rect 154577 8891 154635 8897
rect 154577 8857 154589 8891
rect 154623 8888 154635 8891
rect 158530 8888 158536 8900
rect 154623 8860 158536 8888
rect 154623 8857 154635 8860
rect 154577 8851 154635 8857
rect 158530 8848 158536 8860
rect 158588 8848 158594 8900
rect 152884 8792 154436 8820
rect 152884 8780 152890 8792
rect 155034 8780 155040 8832
rect 155092 8820 155098 8832
rect 155865 8823 155923 8829
rect 155865 8820 155877 8823
rect 155092 8792 155877 8820
rect 155092 8780 155098 8792
rect 155865 8789 155877 8792
rect 155911 8789 155923 8823
rect 155865 8783 155923 8789
rect 156874 8780 156880 8832
rect 156932 8820 156938 8832
rect 157061 8823 157119 8829
rect 157061 8820 157073 8823
rect 156932 8792 157073 8820
rect 156932 8780 156938 8792
rect 157061 8789 157073 8792
rect 157107 8789 157119 8823
rect 157061 8783 157119 8789
rect 1104 8730 159043 8752
rect 1104 8678 40394 8730
rect 40446 8678 40458 8730
rect 40510 8678 40522 8730
rect 40574 8678 40586 8730
rect 40638 8678 40650 8730
rect 40702 8678 79839 8730
rect 79891 8678 79903 8730
rect 79955 8678 79967 8730
rect 80019 8678 80031 8730
rect 80083 8678 80095 8730
rect 80147 8678 119284 8730
rect 119336 8678 119348 8730
rect 119400 8678 119412 8730
rect 119464 8678 119476 8730
rect 119528 8678 119540 8730
rect 119592 8678 158729 8730
rect 158781 8678 158793 8730
rect 158845 8678 158857 8730
rect 158909 8678 158921 8730
rect 158973 8678 158985 8730
rect 159037 8678 159043 8730
rect 1104 8656 159043 8678
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 5868 8588 11805 8616
rect 5868 8576 5874 8588
rect 11793 8585 11805 8588
rect 11839 8616 11851 8619
rect 12434 8616 12440 8628
rect 11839 8588 12440 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 12434 8576 12440 8588
rect 12492 8616 12498 8628
rect 12894 8616 12900 8628
rect 12492 8588 12900 8616
rect 12492 8576 12498 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 18230 8616 18236 8628
rect 13648 8588 18236 8616
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 5184 8480 5212 8576
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 13458 8551 13516 8557
rect 13458 8548 13470 8551
rect 13320 8520 13470 8548
rect 13320 8508 13326 8520
rect 13458 8517 13470 8520
rect 13504 8517 13516 8551
rect 13458 8511 13516 8517
rect 4571 8452 5212 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5592 8452 6009 8480
rect 5592 8440 5598 8452
rect 5997 8449 6009 8452
rect 6043 8480 6055 8483
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6043 8452 6745 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6733 8449 6745 8452
rect 6779 8480 6791 8483
rect 13648 8480 13676 8588
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 18690 8616 18696 8628
rect 18463 8588 18696 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 28534 8616 28540 8628
rect 27540 8588 28304 8616
rect 28495 8588 28540 8616
rect 19444 8548 19472 8576
rect 27540 8548 27568 8588
rect 14660 8520 19472 8548
rect 27172 8520 27568 8548
rect 28276 8548 28304 8588
rect 28534 8576 28540 8588
rect 28592 8576 28598 8628
rect 29546 8616 29552 8628
rect 29507 8588 29552 8616
rect 29546 8576 29552 8588
rect 29604 8576 29610 8628
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 33318 8616 33324 8628
rect 29696 8588 31754 8616
rect 33279 8588 33324 8616
rect 29696 8576 29702 8588
rect 28997 8551 29055 8557
rect 28997 8548 29009 8551
rect 28276 8520 29009 8548
rect 6779 8452 13676 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14660 8489 14688 8520
rect 14918 8489 14924 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13780 8452 14657 8480
rect 13780 8440 13786 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14912 8443 14924 8489
rect 14976 8480 14982 8492
rect 14976 8452 15012 8480
rect 14918 8440 14924 8443
rect 14976 8440 14982 8452
rect 16482 8440 16488 8492
rect 16540 8480 16546 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 16540 8452 17049 8480
rect 16540 8440 16546 8452
rect 17037 8449 17049 8452
rect 17083 8480 17095 8483
rect 17678 8480 17684 8492
rect 17083 8452 17684 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17862 8480 17868 8492
rect 17823 8452 17868 8480
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18288 8452 26280 8480
rect 18288 8440 18294 8452
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8412 3939 8415
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 3927 8384 4353 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 4341 8381 4353 8384
rect 4387 8412 4399 8415
rect 5626 8412 5632 8424
rect 4387 8384 5632 8412
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 16758 8412 16764 8424
rect 6917 8375 6975 8381
rect 16040 8384 16764 8412
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 5408 8316 6561 8344
rect 5408 8304 5414 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 6932 8344 6960 8375
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 6788 8316 7481 8344
rect 6788 8304 6794 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 4709 8279 4767 8285
rect 4709 8245 4721 8279
rect 4755 8276 4767 8279
rect 5074 8276 5080 8288
rect 4755 8248 5080 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 7484 8276 7512 8307
rect 8202 8304 8208 8356
rect 8260 8304 8266 8356
rect 11974 8304 11980 8356
rect 12032 8344 12038 8356
rect 16040 8353 16068 8384
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 17221 8415 17279 8421
rect 16908 8384 16953 8412
rect 16908 8372 16914 8384
rect 17221 8381 17233 8415
rect 17267 8412 17279 8415
rect 19794 8412 19800 8424
rect 17267 8384 19800 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 26252 8412 26280 8452
rect 26326 8440 26332 8492
rect 26384 8480 26390 8492
rect 27172 8489 27200 8520
rect 28997 8517 29009 8520
rect 29043 8548 29055 8551
rect 29086 8548 29092 8560
rect 29043 8520 29092 8548
rect 29043 8517 29055 8520
rect 28997 8511 29055 8517
rect 29086 8508 29092 8520
rect 29144 8548 29150 8560
rect 30101 8551 30159 8557
rect 30101 8548 30113 8551
rect 29144 8520 30113 8548
rect 29144 8508 29150 8520
rect 30101 8517 30113 8520
rect 30147 8548 30159 8551
rect 31018 8548 31024 8560
rect 30147 8520 31024 8548
rect 30147 8517 30159 8520
rect 30101 8511 30159 8517
rect 31018 8508 31024 8520
rect 31076 8508 31082 8560
rect 31726 8548 31754 8588
rect 33318 8576 33324 8588
rect 33376 8576 33382 8628
rect 34238 8576 34244 8628
rect 34296 8616 34302 8628
rect 35250 8616 35256 8628
rect 34296 8588 35256 8616
rect 34296 8576 34302 8588
rect 35250 8576 35256 8588
rect 35308 8576 35314 8628
rect 35894 8616 35900 8628
rect 35855 8588 35900 8616
rect 35894 8576 35900 8588
rect 35952 8576 35958 8628
rect 41046 8616 41052 8628
rect 36556 8588 41052 8616
rect 36556 8548 36584 8588
rect 41046 8576 41052 8588
rect 41104 8576 41110 8628
rect 41782 8576 41788 8628
rect 41840 8616 41846 8628
rect 45281 8619 45339 8625
rect 45281 8616 45293 8619
rect 41840 8588 45293 8616
rect 41840 8576 41846 8588
rect 45281 8585 45293 8588
rect 45327 8585 45339 8619
rect 45281 8579 45339 8585
rect 45462 8576 45468 8628
rect 45520 8616 45526 8628
rect 45646 8616 45652 8628
rect 45520 8588 45652 8616
rect 45520 8576 45526 8588
rect 45646 8576 45652 8588
rect 45704 8616 45710 8628
rect 45922 8616 45928 8628
rect 45704 8588 45928 8616
rect 45704 8576 45710 8588
rect 45922 8576 45928 8588
rect 45980 8576 45986 8628
rect 48777 8619 48835 8625
rect 48777 8616 48789 8619
rect 46308 8588 48789 8616
rect 37642 8548 37648 8560
rect 31726 8520 36584 8548
rect 36740 8520 37648 8548
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26384 8452 27169 8480
rect 26384 8440 26390 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27246 8440 27252 8492
rect 27304 8480 27310 8492
rect 27413 8483 27471 8489
rect 27413 8480 27425 8483
rect 27304 8452 27425 8480
rect 27304 8440 27310 8452
rect 27413 8449 27425 8452
rect 27459 8449 27471 8483
rect 27413 8443 27471 8449
rect 27706 8440 27712 8492
rect 27764 8480 27770 8492
rect 30466 8480 30472 8492
rect 27764 8452 30472 8480
rect 27764 8440 27770 8452
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 30840 8476 30898 8479
rect 30834 8464 30840 8476
rect 30804 8436 30840 8464
rect 30834 8424 30840 8436
rect 30892 8424 30898 8476
rect 33134 8440 33140 8492
rect 33192 8480 33198 8492
rect 33505 8483 33563 8489
rect 33505 8480 33517 8483
rect 33192 8452 33517 8480
rect 33192 8440 33198 8452
rect 33505 8449 33517 8452
rect 33551 8449 33563 8483
rect 35078 8483 35136 8489
rect 35078 8480 35090 8483
rect 33505 8443 33563 8449
rect 33612 8452 35090 8480
rect 20036 8384 22094 8412
rect 26252 8384 27200 8412
rect 20036 8372 20042 8384
rect 12345 8347 12403 8353
rect 12345 8344 12357 8347
rect 12032 8316 12357 8344
rect 12032 8304 12038 8316
rect 12345 8313 12357 8316
rect 12391 8313 12403 8347
rect 12345 8307 12403 8313
rect 16025 8347 16083 8353
rect 16025 8313 16037 8347
rect 16071 8313 16083 8347
rect 16025 8307 16083 8313
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 17681 8347 17739 8353
rect 17681 8344 17693 8347
rect 16540 8316 17693 8344
rect 16540 8304 16546 8316
rect 17681 8313 17693 8316
rect 17727 8313 17739 8347
rect 17681 8307 17739 8313
rect 17770 8304 17776 8356
rect 17828 8344 17834 8356
rect 21910 8344 21916 8356
rect 17828 8316 21916 8344
rect 17828 8304 17834 8316
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 22066 8344 22094 8384
rect 27062 8344 27068 8356
rect 22066 8316 27068 8344
rect 27062 8304 27068 8316
rect 27120 8304 27126 8356
rect 8220 8276 8248 8304
rect 8662 8276 8668 8288
rect 7484 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 14274 8276 14280 8288
rect 10744 8248 14280 8276
rect 10744 8236 10750 8248
rect 14274 8236 14280 8248
rect 14332 8276 14338 8288
rect 15746 8276 15752 8288
rect 14332 8248 15752 8276
rect 14332 8236 14338 8248
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 16942 8236 16948 8288
rect 17000 8276 17006 8288
rect 17310 8276 17316 8288
rect 17000 8248 17316 8276
rect 17000 8236 17006 8248
rect 17310 8236 17316 8248
rect 17368 8276 17374 8288
rect 18877 8279 18935 8285
rect 18877 8276 18889 8279
rect 17368 8248 18889 8276
rect 17368 8236 17374 8248
rect 18877 8245 18889 8248
rect 18923 8245 18935 8279
rect 18877 8239 18935 8245
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 24210 8276 24216 8288
rect 19024 8248 24216 8276
rect 19024 8236 19030 8248
rect 24210 8236 24216 8248
rect 24268 8236 24274 8288
rect 27172 8276 27200 8384
rect 28166 8372 28172 8424
rect 28224 8412 28230 8424
rect 29638 8412 29644 8424
rect 28224 8384 29644 8412
rect 28224 8372 28230 8384
rect 29638 8372 29644 8384
rect 29696 8372 29702 8424
rect 30558 8372 30564 8424
rect 30616 8412 30622 8424
rect 30653 8415 30711 8421
rect 30653 8412 30665 8415
rect 30616 8384 30665 8412
rect 30616 8372 30622 8384
rect 30653 8381 30665 8384
rect 30699 8381 30711 8415
rect 30653 8375 30711 8381
rect 31021 8415 31079 8421
rect 31021 8381 31033 8415
rect 31067 8412 31079 8415
rect 31110 8412 31116 8424
rect 31067 8384 31116 8412
rect 31067 8381 31079 8384
rect 31021 8375 31079 8381
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 31757 8415 31815 8421
rect 31757 8381 31769 8415
rect 31803 8412 31815 8415
rect 33612 8412 33640 8452
rect 35078 8449 35090 8452
rect 35124 8449 35136 8483
rect 35078 8443 35136 8449
rect 35250 8440 35256 8492
rect 35308 8480 35314 8492
rect 35345 8483 35403 8489
rect 35345 8480 35357 8483
rect 35308 8452 35357 8480
rect 35308 8440 35314 8452
rect 35345 8449 35357 8452
rect 35391 8449 35403 8483
rect 36538 8480 36544 8492
rect 36499 8452 36544 8480
rect 35345 8443 35403 8449
rect 36538 8440 36544 8452
rect 36596 8440 36602 8492
rect 36740 8489 36768 8520
rect 37642 8508 37648 8520
rect 37700 8548 37706 8560
rect 38470 8548 38476 8560
rect 37700 8520 38476 8548
rect 37700 8508 37706 8520
rect 38470 8508 38476 8520
rect 38528 8508 38534 8560
rect 38930 8557 38936 8560
rect 38924 8511 38936 8557
rect 38988 8548 38994 8560
rect 38988 8520 39024 8548
rect 38930 8508 38936 8511
rect 38988 8508 38994 8520
rect 39390 8508 39396 8560
rect 39448 8548 39454 8560
rect 40681 8551 40739 8557
rect 40681 8548 40693 8551
rect 39448 8520 40693 8548
rect 39448 8508 39454 8520
rect 40681 8517 40693 8520
rect 40727 8517 40739 8551
rect 46308 8548 46336 8588
rect 48777 8585 48789 8588
rect 48823 8585 48835 8619
rect 49418 8616 49424 8628
rect 49379 8588 49424 8616
rect 48777 8579 48835 8585
rect 49418 8576 49424 8588
rect 49476 8576 49482 8628
rect 51442 8616 51448 8628
rect 51403 8588 51448 8616
rect 51442 8576 51448 8588
rect 51500 8576 51506 8628
rect 53469 8619 53527 8625
rect 53469 8585 53481 8619
rect 53515 8616 53527 8619
rect 56045 8619 56103 8625
rect 56045 8616 56057 8619
rect 53515 8588 56057 8616
rect 53515 8585 53527 8588
rect 53469 8579 53527 8585
rect 56045 8585 56057 8588
rect 56091 8616 56103 8619
rect 56134 8616 56140 8628
rect 56091 8588 56140 8616
rect 56091 8585 56103 8588
rect 56045 8579 56103 8585
rect 56134 8576 56140 8588
rect 56192 8576 56198 8628
rect 59998 8616 60004 8628
rect 59959 8588 60004 8616
rect 59998 8576 60004 8588
rect 60056 8576 60062 8628
rect 61381 8619 61439 8625
rect 61381 8585 61393 8619
rect 61427 8616 61439 8619
rect 62206 8616 62212 8628
rect 61427 8588 62212 8616
rect 61427 8585 61439 8588
rect 61381 8579 61439 8585
rect 40681 8511 40739 8517
rect 44100 8520 46336 8548
rect 36725 8483 36783 8489
rect 36725 8449 36737 8483
rect 36771 8449 36783 8483
rect 37826 8480 37832 8492
rect 37787 8452 37832 8480
rect 36725 8443 36783 8449
rect 37826 8440 37832 8452
rect 37884 8440 37890 8492
rect 38010 8480 38016 8492
rect 37971 8452 38016 8480
rect 38010 8440 38016 8452
rect 38068 8440 38074 8492
rect 38654 8480 38660 8492
rect 38615 8452 38660 8480
rect 38654 8440 38660 8452
rect 38712 8440 38718 8492
rect 38764 8452 39712 8480
rect 31803 8384 33640 8412
rect 36556 8412 36584 8440
rect 36998 8412 37004 8424
rect 36556 8384 37004 8412
rect 31803 8381 31815 8384
rect 31757 8375 31815 8381
rect 31772 8344 31800 8375
rect 36998 8372 37004 8384
rect 37056 8412 37062 8424
rect 38764 8412 38792 8452
rect 37056 8384 38792 8412
rect 37056 8372 37062 8384
rect 33965 8347 34023 8353
rect 33965 8344 33977 8347
rect 28092 8316 31800 8344
rect 31864 8316 33977 8344
rect 28092 8276 28120 8316
rect 27172 8248 28120 8276
rect 31386 8236 31392 8288
rect 31444 8276 31450 8288
rect 31864 8276 31892 8316
rect 33965 8313 33977 8316
rect 34011 8313 34023 8347
rect 33965 8307 34023 8313
rect 36357 8347 36415 8353
rect 36357 8313 36369 8347
rect 36403 8344 36415 8347
rect 36538 8344 36544 8356
rect 36403 8316 36544 8344
rect 36403 8313 36415 8316
rect 36357 8307 36415 8313
rect 36538 8304 36544 8316
rect 36596 8304 36602 8356
rect 38197 8347 38255 8353
rect 38197 8313 38209 8347
rect 38243 8344 38255 8347
rect 38243 8316 38700 8344
rect 38243 8313 38255 8316
rect 38197 8307 38255 8313
rect 31444 8248 31892 8276
rect 32861 8279 32919 8285
rect 31444 8236 31450 8248
rect 32861 8245 32873 8279
rect 32907 8276 32919 8279
rect 32950 8276 32956 8288
rect 32907 8248 32956 8276
rect 32907 8245 32919 8248
rect 32861 8239 32919 8245
rect 32950 8236 32956 8248
rect 33008 8236 33014 8288
rect 38672 8276 38700 8316
rect 39298 8276 39304 8288
rect 38672 8248 39304 8276
rect 39298 8236 39304 8248
rect 39356 8236 39362 8288
rect 39684 8276 39712 8452
rect 41138 8440 41144 8492
rect 41196 8480 41202 8492
rect 41233 8483 41291 8489
rect 41233 8480 41245 8483
rect 41196 8452 41245 8480
rect 41196 8440 41202 8452
rect 41233 8449 41245 8452
rect 41279 8449 41291 8483
rect 41233 8443 41291 8449
rect 41417 8483 41475 8489
rect 41417 8449 41429 8483
rect 41463 8449 41475 8483
rect 41417 8443 41475 8449
rect 41509 8483 41567 8489
rect 41509 8449 41521 8483
rect 41555 8449 41567 8483
rect 41509 8443 41567 8449
rect 43737 8483 43795 8489
rect 43737 8449 43749 8483
rect 43783 8480 43795 8483
rect 44100 8480 44128 8520
rect 46382 8508 46388 8560
rect 46440 8557 46446 8560
rect 46440 8548 46452 8557
rect 50430 8548 50436 8560
rect 46440 8520 46485 8548
rect 48976 8520 50436 8548
rect 46440 8511 46452 8520
rect 46440 8508 46446 8511
rect 43783 8452 44128 8480
rect 43783 8449 43795 8452
rect 43737 8443 43795 8449
rect 40037 8347 40095 8353
rect 40037 8313 40049 8347
rect 40083 8344 40095 8347
rect 40770 8344 40776 8356
rect 40083 8316 40776 8344
rect 40083 8313 40095 8316
rect 40037 8307 40095 8313
rect 40770 8304 40776 8316
rect 40828 8304 40834 8356
rect 41230 8304 41236 8356
rect 41288 8344 41294 8356
rect 41432 8344 41460 8443
rect 41288 8316 41460 8344
rect 41524 8344 41552 8443
rect 44174 8440 44180 8492
rect 44232 8480 44238 8492
rect 44637 8483 44695 8489
rect 44637 8480 44649 8483
rect 44232 8452 44649 8480
rect 44232 8440 44238 8452
rect 44637 8449 44649 8452
rect 44683 8449 44695 8483
rect 44637 8443 44695 8449
rect 44726 8440 44732 8492
rect 44784 8480 44790 8492
rect 48317 8483 48375 8489
rect 48317 8480 48329 8483
rect 44784 8452 48329 8480
rect 44784 8440 44790 8452
rect 48317 8449 48329 8452
rect 48363 8480 48375 8483
rect 48866 8480 48872 8492
rect 48363 8452 48872 8480
rect 48363 8449 48375 8452
rect 48317 8443 48375 8449
rect 48866 8440 48872 8452
rect 48924 8440 48930 8492
rect 48976 8489 49004 8520
rect 50430 8508 50436 8520
rect 50488 8508 50494 8560
rect 53374 8508 53380 8560
rect 53432 8548 53438 8560
rect 55042 8551 55100 8557
rect 55042 8548 55054 8551
rect 53432 8520 55054 8548
rect 53432 8508 53438 8520
rect 55042 8517 55054 8520
rect 55088 8517 55100 8551
rect 55042 8511 55100 8517
rect 55214 8508 55220 8560
rect 55272 8548 55278 8560
rect 58066 8548 58072 8560
rect 55272 8520 58072 8548
rect 55272 8508 55278 8520
rect 58066 8508 58072 8520
rect 58124 8508 58130 8560
rect 58336 8551 58394 8557
rect 58336 8517 58348 8551
rect 58382 8548 58394 8551
rect 60826 8548 60832 8560
rect 58382 8520 60832 8548
rect 58382 8517 58394 8520
rect 58336 8511 58394 8517
rect 60826 8508 60832 8520
rect 60884 8508 60890 8560
rect 48961 8483 49019 8489
rect 48961 8449 48973 8483
rect 49007 8449 49019 8483
rect 48961 8443 49019 8449
rect 49142 8440 49148 8492
rect 49200 8480 49206 8492
rect 50534 8483 50592 8489
rect 50534 8480 50546 8483
rect 49200 8452 50546 8480
rect 49200 8440 49206 8452
rect 50534 8449 50546 8452
rect 50580 8449 50592 8483
rect 52178 8480 52184 8492
rect 52139 8452 52184 8480
rect 50534 8443 50592 8449
rect 52178 8440 52184 8452
rect 52236 8440 52242 8492
rect 52270 8440 52276 8492
rect 52328 8480 52334 8492
rect 52328 8452 52373 8480
rect 52328 8440 52334 8452
rect 52546 8440 52552 8492
rect 52604 8480 52610 8492
rect 55309 8483 55367 8489
rect 55309 8480 55321 8483
rect 52604 8452 55321 8480
rect 52604 8440 52610 8452
rect 55309 8449 55321 8452
rect 55355 8480 55367 8483
rect 55674 8480 55680 8492
rect 55355 8452 55680 8480
rect 55355 8449 55367 8452
rect 55309 8443 55367 8449
rect 55674 8440 55680 8452
rect 55732 8440 55738 8492
rect 56689 8483 56747 8489
rect 56689 8449 56701 8483
rect 56735 8480 56747 8483
rect 57149 8483 57207 8489
rect 57149 8480 57161 8483
rect 56735 8452 57161 8480
rect 56735 8449 56747 8452
rect 56689 8443 56747 8449
rect 57149 8449 57161 8452
rect 57195 8449 57207 8483
rect 57330 8480 57336 8492
rect 57291 8452 57336 8480
rect 57149 8443 57207 8449
rect 57330 8440 57336 8452
rect 57388 8440 57394 8492
rect 59814 8480 59820 8492
rect 57440 8452 59820 8480
rect 43990 8372 43996 8424
rect 44048 8412 44054 8424
rect 45370 8412 45376 8424
rect 44048 8384 45376 8412
rect 44048 8372 44054 8384
rect 45370 8372 45376 8384
rect 45428 8372 45434 8424
rect 46658 8372 46664 8424
rect 46716 8412 46722 8424
rect 49786 8412 49792 8424
rect 46716 8384 49792 8412
rect 46716 8372 46722 8384
rect 49786 8372 49792 8384
rect 49844 8372 49850 8424
rect 50801 8415 50859 8421
rect 50801 8381 50813 8415
rect 50847 8412 50859 8415
rect 51074 8412 51080 8424
rect 50847 8384 51080 8412
rect 50847 8381 50859 8384
rect 50801 8375 50859 8381
rect 51074 8372 51080 8384
rect 51132 8372 51138 8424
rect 51350 8372 51356 8424
rect 51408 8412 51414 8424
rect 52086 8412 52092 8424
rect 51408 8384 52092 8412
rect 51408 8372 51414 8384
rect 52086 8372 52092 8384
rect 52144 8372 52150 8424
rect 52730 8372 52736 8424
rect 52788 8412 52794 8424
rect 54110 8412 54116 8424
rect 52788 8384 54116 8412
rect 52788 8372 52794 8384
rect 54110 8372 54116 8384
rect 54168 8372 54174 8424
rect 57440 8412 57468 8452
rect 59814 8440 59820 8452
rect 59872 8440 59878 8492
rect 60642 8480 60648 8492
rect 60603 8452 60648 8480
rect 60642 8440 60648 8452
rect 60700 8440 60706 8492
rect 60737 8483 60795 8489
rect 60737 8449 60749 8483
rect 60783 8480 60795 8483
rect 61396 8480 61424 8579
rect 62206 8576 62212 8588
rect 62264 8576 62270 8628
rect 62666 8616 62672 8628
rect 62627 8588 62672 8616
rect 62666 8576 62672 8588
rect 62724 8576 62730 8628
rect 63773 8619 63831 8625
rect 63773 8585 63785 8619
rect 63819 8616 63831 8619
rect 65150 8616 65156 8628
rect 63819 8588 65156 8616
rect 63819 8585 63831 8588
rect 63773 8579 63831 8585
rect 65150 8576 65156 8588
rect 65208 8576 65214 8628
rect 67450 8616 67456 8628
rect 67411 8588 67456 8616
rect 67450 8576 67456 8588
rect 67508 8576 67514 8628
rect 69750 8616 69756 8628
rect 69711 8588 69756 8616
rect 69750 8576 69756 8588
rect 69808 8576 69814 8628
rect 69842 8576 69848 8628
rect 69900 8616 69906 8628
rect 83918 8616 83924 8628
rect 69900 8588 83924 8616
rect 69900 8576 69906 8588
rect 83918 8576 83924 8588
rect 83976 8576 83982 8628
rect 84010 8576 84016 8628
rect 84068 8616 84074 8628
rect 88981 8619 89039 8625
rect 84068 8588 88932 8616
rect 84068 8576 84074 8588
rect 64230 8548 64236 8560
rect 64191 8520 64236 8548
rect 64230 8508 64236 8520
rect 64288 8508 64294 8560
rect 85206 8548 85212 8560
rect 65536 8520 85212 8548
rect 60783 8452 61424 8480
rect 60783 8449 60795 8452
rect 60737 8443 60795 8449
rect 55324 8384 57468 8412
rect 42058 8344 42064 8356
rect 41524 8316 42064 8344
rect 41288 8304 41294 8316
rect 42058 8304 42064 8316
rect 42116 8304 42122 8356
rect 44082 8304 44088 8356
rect 44140 8344 44146 8356
rect 44453 8347 44511 8353
rect 44453 8344 44465 8347
rect 44140 8316 44465 8344
rect 44140 8304 44146 8316
rect 44453 8313 44465 8316
rect 44499 8313 44511 8347
rect 44453 8307 44511 8313
rect 50982 8304 50988 8356
rect 51040 8344 51046 8356
rect 51997 8347 52055 8353
rect 51997 8344 52009 8347
rect 51040 8316 52009 8344
rect 51040 8304 51046 8316
rect 51997 8313 52009 8316
rect 52043 8313 52055 8347
rect 53926 8344 53932 8356
rect 53887 8316 53932 8344
rect 51997 8307 52055 8313
rect 53926 8304 53932 8316
rect 53984 8304 53990 8356
rect 41782 8276 41788 8288
rect 39684 8248 41788 8276
rect 41782 8236 41788 8248
rect 41840 8236 41846 8288
rect 42334 8236 42340 8288
rect 42392 8276 42398 8288
rect 42613 8279 42671 8285
rect 42613 8276 42625 8279
rect 42392 8248 42625 8276
rect 42392 8236 42398 8248
rect 42613 8245 42625 8248
rect 42659 8276 42671 8279
rect 46014 8276 46020 8288
rect 42659 8248 46020 8276
rect 42659 8245 42671 8248
rect 42613 8239 42671 8245
rect 46014 8236 46020 8248
rect 46072 8236 46078 8288
rect 46750 8236 46756 8288
rect 46808 8276 46814 8288
rect 47026 8276 47032 8288
rect 46808 8248 47032 8276
rect 46808 8236 46814 8248
rect 47026 8236 47032 8248
rect 47084 8276 47090 8288
rect 47121 8279 47179 8285
rect 47121 8276 47133 8279
rect 47084 8248 47133 8276
rect 47084 8236 47090 8248
rect 47121 8245 47133 8248
rect 47167 8245 47179 8279
rect 47121 8239 47179 8245
rect 51902 8236 51908 8288
rect 51960 8276 51966 8288
rect 54202 8276 54208 8288
rect 51960 8248 54208 8276
rect 51960 8236 51966 8248
rect 54202 8236 54208 8248
rect 54260 8236 54266 8288
rect 54570 8236 54576 8288
rect 54628 8276 54634 8288
rect 55324 8276 55352 8384
rect 57514 8372 57520 8424
rect 57572 8412 57578 8424
rect 58069 8415 58127 8421
rect 57572 8384 57617 8412
rect 57572 8372 57578 8384
rect 58069 8381 58081 8415
rect 58115 8381 58127 8415
rect 58069 8375 58127 8381
rect 56042 8304 56048 8356
rect 56100 8344 56106 8356
rect 56505 8347 56563 8353
rect 56505 8344 56517 8347
rect 56100 8316 56517 8344
rect 56100 8304 56106 8316
rect 56505 8313 56517 8316
rect 56551 8313 56563 8347
rect 56505 8307 56563 8313
rect 54628 8248 55352 8276
rect 58084 8276 58112 8375
rect 59722 8372 59728 8424
rect 59780 8412 59786 8424
rect 60752 8412 60780 8443
rect 59780 8384 60780 8412
rect 59780 8372 59786 8384
rect 59449 8347 59507 8353
rect 59449 8313 59461 8347
rect 59495 8344 59507 8347
rect 65536 8344 65564 8520
rect 85206 8508 85212 8520
rect 85264 8508 85270 8560
rect 87874 8508 87880 8560
rect 87932 8557 87938 8560
rect 87932 8548 87944 8557
rect 88904 8548 88932 8588
rect 88981 8585 88993 8619
rect 89027 8616 89039 8619
rect 89346 8616 89352 8628
rect 89027 8588 89352 8616
rect 89027 8585 89039 8588
rect 88981 8579 89039 8585
rect 89346 8576 89352 8588
rect 89404 8576 89410 8628
rect 89438 8576 89444 8628
rect 89496 8616 89502 8628
rect 117314 8616 117320 8628
rect 89496 8588 117320 8616
rect 89496 8576 89502 8588
rect 117314 8576 117320 8588
rect 117372 8616 117378 8628
rect 117409 8619 117467 8625
rect 117409 8616 117421 8619
rect 117372 8588 117421 8616
rect 117372 8576 117378 8588
rect 117409 8585 117421 8588
rect 117455 8585 117467 8619
rect 117409 8579 117467 8585
rect 117498 8576 117504 8628
rect 117556 8616 117562 8628
rect 121914 8616 121920 8628
rect 117556 8588 121920 8616
rect 117556 8576 117562 8588
rect 121914 8576 121920 8588
rect 121972 8576 121978 8628
rect 122377 8619 122435 8625
rect 122377 8585 122389 8619
rect 122423 8585 122435 8619
rect 130565 8619 130623 8625
rect 122377 8579 122435 8585
rect 122475 8588 130516 8616
rect 90910 8548 90916 8560
rect 87932 8520 87977 8548
rect 88904 8520 90916 8548
rect 87932 8511 87944 8520
rect 87932 8508 87938 8511
rect 90910 8508 90916 8520
rect 90968 8508 90974 8560
rect 92474 8508 92480 8560
rect 92532 8548 92538 8560
rect 108666 8548 108672 8560
rect 92532 8520 108672 8548
rect 92532 8508 92538 8520
rect 108666 8508 108672 8520
rect 108724 8508 108730 8560
rect 112165 8551 112223 8557
rect 112165 8548 112177 8551
rect 109696 8520 112177 8548
rect 67634 8480 67640 8492
rect 67595 8452 67640 8480
rect 67634 8440 67640 8452
rect 67692 8440 67698 8492
rect 68640 8483 68698 8489
rect 68640 8449 68652 8483
rect 68686 8480 68698 8483
rect 70210 8480 70216 8492
rect 68686 8452 70216 8480
rect 68686 8449 68698 8452
rect 68640 8443 68698 8449
rect 70210 8440 70216 8452
rect 70268 8440 70274 8492
rect 72326 8440 72332 8492
rect 72384 8480 72390 8492
rect 76018 8483 76076 8489
rect 76018 8480 76030 8483
rect 72384 8452 76030 8480
rect 72384 8440 72390 8452
rect 76018 8449 76030 8452
rect 76064 8449 76076 8483
rect 76018 8443 76076 8449
rect 76285 8483 76343 8489
rect 76285 8449 76297 8483
rect 76331 8480 76343 8483
rect 76466 8480 76472 8492
rect 76331 8452 76472 8480
rect 76331 8449 76343 8452
rect 76285 8443 76343 8449
rect 76466 8440 76472 8452
rect 76524 8440 76530 8492
rect 76558 8440 76564 8492
rect 76616 8480 76622 8492
rect 76745 8483 76803 8489
rect 76745 8480 76757 8483
rect 76616 8452 76757 8480
rect 76616 8440 76622 8452
rect 76745 8449 76757 8452
rect 76791 8449 76803 8483
rect 76745 8443 76803 8449
rect 77012 8483 77070 8489
rect 77012 8449 77024 8483
rect 77058 8480 77070 8483
rect 83642 8480 83648 8492
rect 77058 8452 83648 8480
rect 77058 8449 77070 8452
rect 77012 8443 77070 8449
rect 83642 8440 83648 8452
rect 83700 8440 83706 8492
rect 83826 8480 83832 8492
rect 83787 8452 83832 8480
rect 83826 8440 83832 8452
rect 83884 8440 83890 8492
rect 88153 8483 88211 8489
rect 84028 8452 88104 8480
rect 67818 8412 67824 8424
rect 67731 8384 67824 8412
rect 67818 8372 67824 8384
rect 67876 8372 67882 8424
rect 68370 8412 68376 8424
rect 68331 8384 68376 8412
rect 68370 8372 68376 8384
rect 68428 8372 68434 8424
rect 73338 8372 73344 8424
rect 73396 8412 73402 8424
rect 73396 8384 74948 8412
rect 73396 8372 73402 8384
rect 59495 8316 65564 8344
rect 59495 8313 59507 8316
rect 59449 8307 59507 8313
rect 65886 8304 65892 8356
rect 65944 8344 65950 8356
rect 66901 8347 66959 8353
rect 66901 8344 66913 8347
rect 65944 8316 66913 8344
rect 65944 8304 65950 8316
rect 66901 8313 66913 8316
rect 66947 8344 66959 8347
rect 67836 8344 67864 8372
rect 66947 8316 67864 8344
rect 66947 8313 66959 8316
rect 66901 8307 66959 8313
rect 73154 8304 73160 8356
rect 73212 8344 73218 8356
rect 74920 8353 74948 8384
rect 73525 8347 73583 8353
rect 73525 8344 73537 8347
rect 73212 8316 73537 8344
rect 73212 8304 73218 8316
rect 73525 8313 73537 8316
rect 73571 8313 73583 8347
rect 73525 8307 73583 8313
rect 74905 8347 74963 8353
rect 74905 8313 74917 8347
rect 74951 8313 74963 8347
rect 74905 8307 74963 8313
rect 78125 8347 78183 8353
rect 78125 8313 78137 8347
rect 78171 8344 78183 8347
rect 78858 8344 78864 8356
rect 78171 8316 78864 8344
rect 78171 8313 78183 8316
rect 78125 8307 78183 8313
rect 78858 8304 78864 8316
rect 78916 8344 78922 8356
rect 80330 8344 80336 8356
rect 78916 8316 80336 8344
rect 78916 8304 78922 8316
rect 80330 8304 80336 8316
rect 80388 8304 80394 8356
rect 84028 8353 84056 8452
rect 88076 8412 88104 8452
rect 88153 8449 88165 8483
rect 88199 8480 88211 8483
rect 88426 8480 88432 8492
rect 88199 8452 88432 8480
rect 88199 8449 88211 8452
rect 88153 8443 88211 8449
rect 88426 8440 88432 8452
rect 88484 8440 88490 8492
rect 90082 8440 90088 8492
rect 90140 8489 90146 8492
rect 90140 8480 90152 8489
rect 90140 8452 90185 8480
rect 90140 8443 90152 8452
rect 90140 8440 90146 8443
rect 90450 8440 90456 8492
rect 90508 8480 90514 8492
rect 91002 8480 91008 8492
rect 90508 8452 91008 8480
rect 90508 8440 90514 8452
rect 91002 8440 91008 8452
rect 91060 8440 91066 8492
rect 91922 8440 91928 8492
rect 91980 8489 91986 8492
rect 92198 8489 92204 8492
rect 91980 8443 91992 8489
rect 92194 8443 92204 8489
rect 92256 8480 92262 8492
rect 92256 8452 92294 8480
rect 91980 8440 91986 8443
rect 92198 8440 92204 8443
rect 92256 8440 92262 8452
rect 92382 8440 92388 8492
rect 92440 8480 92446 8492
rect 92440 8452 94268 8480
rect 92440 8440 92446 8452
rect 88886 8412 88892 8424
rect 88076 8384 88892 8412
rect 88886 8372 88892 8384
rect 88944 8372 88950 8424
rect 90358 8412 90364 8424
rect 90319 8384 90364 8412
rect 90358 8372 90364 8384
rect 90416 8412 90422 8424
rect 90910 8412 90916 8424
rect 90416 8384 90916 8412
rect 90416 8372 90422 8384
rect 90910 8372 90916 8384
rect 90968 8372 90974 8424
rect 92290 8372 92296 8424
rect 92348 8412 92354 8424
rect 92348 8384 93348 8412
rect 92348 8372 92354 8384
rect 93320 8356 93348 8384
rect 94038 8372 94044 8424
rect 94096 8412 94102 8424
rect 94133 8415 94191 8421
rect 94133 8412 94145 8415
rect 94096 8384 94145 8412
rect 94096 8372 94102 8384
rect 94133 8381 94145 8384
rect 94179 8381 94191 8415
rect 94240 8412 94268 8452
rect 94314 8440 94320 8492
rect 94372 8480 94378 8492
rect 98178 8480 98184 8492
rect 94372 8452 94417 8480
rect 98139 8452 98184 8480
rect 94372 8440 94378 8452
rect 98178 8440 98184 8452
rect 98236 8480 98242 8492
rect 98236 8452 100984 8480
rect 98236 8440 98242 8452
rect 100386 8412 100392 8424
rect 94240 8384 100392 8412
rect 94133 8375 94191 8381
rect 100386 8372 100392 8384
rect 100444 8372 100450 8424
rect 100956 8412 100984 8452
rect 101030 8440 101036 8492
rect 101088 8480 101094 8492
rect 107013 8483 107071 8489
rect 107013 8480 107025 8483
rect 101088 8452 107025 8480
rect 101088 8440 101094 8452
rect 107013 8449 107025 8452
rect 107059 8480 107071 8483
rect 107562 8480 107568 8492
rect 107059 8452 107568 8480
rect 107059 8449 107071 8452
rect 107013 8443 107071 8449
rect 107562 8440 107568 8452
rect 107620 8440 107626 8492
rect 107930 8440 107936 8492
rect 107988 8480 107994 8492
rect 108301 8483 108359 8489
rect 108301 8480 108313 8483
rect 107988 8452 108313 8480
rect 107988 8440 107994 8452
rect 108301 8449 108313 8452
rect 108347 8449 108359 8483
rect 108301 8443 108359 8449
rect 108482 8440 108488 8492
rect 108540 8480 108546 8492
rect 108945 8483 109003 8489
rect 108945 8480 108957 8483
rect 108540 8452 108957 8480
rect 108540 8440 108546 8452
rect 108945 8449 108957 8452
rect 108991 8449 109003 8483
rect 108945 8443 109003 8449
rect 109126 8440 109132 8492
rect 109184 8480 109190 8492
rect 109586 8480 109592 8492
rect 109184 8452 109592 8480
rect 109184 8440 109190 8452
rect 109586 8440 109592 8452
rect 109644 8440 109650 8492
rect 107286 8412 107292 8424
rect 100956 8384 107292 8412
rect 107286 8372 107292 8384
rect 107344 8372 107350 8424
rect 107378 8372 107384 8424
rect 107436 8412 107442 8424
rect 109696 8412 109724 8520
rect 112165 8517 112177 8520
rect 112211 8548 112223 8551
rect 112346 8548 112352 8560
rect 112211 8520 112352 8548
rect 112211 8517 112223 8520
rect 112165 8511 112223 8517
rect 112346 8508 112352 8520
rect 112404 8508 112410 8560
rect 115290 8548 115296 8560
rect 115251 8520 115296 8548
rect 115290 8508 115296 8520
rect 115348 8508 115354 8560
rect 120712 8551 120770 8557
rect 115400 8520 120672 8548
rect 109856 8483 109914 8489
rect 109856 8449 109868 8483
rect 109902 8480 109914 8483
rect 109902 8452 111564 8480
rect 109902 8449 109914 8452
rect 109856 8443 109914 8449
rect 111536 8421 111564 8452
rect 112714 8440 112720 8492
rect 112772 8480 112778 8492
rect 112809 8483 112867 8489
rect 112809 8480 112821 8483
rect 112772 8452 112821 8480
rect 112772 8440 112778 8452
rect 112809 8449 112821 8452
rect 112855 8480 112867 8483
rect 115400 8480 115428 8520
rect 112855 8452 115428 8480
rect 112855 8449 112867 8452
rect 112809 8443 112867 8449
rect 115566 8440 115572 8492
rect 115624 8480 115630 8492
rect 115624 8452 117268 8480
rect 115624 8440 115630 8452
rect 107436 8384 109724 8412
rect 111521 8415 111579 8421
rect 107436 8372 107442 8384
rect 111521 8381 111533 8415
rect 111567 8412 111579 8415
rect 114186 8412 114192 8424
rect 111567 8384 114192 8412
rect 111567 8381 111579 8384
rect 111521 8375 111579 8381
rect 114186 8372 114192 8384
rect 114244 8372 114250 8424
rect 116397 8415 116455 8421
rect 116397 8381 116409 8415
rect 116443 8412 116455 8415
rect 116670 8412 116676 8424
rect 116443 8384 116676 8412
rect 116443 8381 116455 8384
rect 116397 8375 116455 8381
rect 116670 8372 116676 8384
rect 116728 8372 116734 8424
rect 117240 8412 117268 8452
rect 117314 8440 117320 8492
rect 117372 8480 117378 8492
rect 118145 8483 118203 8489
rect 118145 8480 118157 8483
rect 117372 8452 118157 8480
rect 117372 8440 117378 8452
rect 118145 8449 118157 8452
rect 118191 8449 118203 8483
rect 118970 8480 118976 8492
rect 118931 8452 118976 8480
rect 118145 8443 118203 8449
rect 118970 8440 118976 8452
rect 119028 8440 119034 8492
rect 120644 8480 120672 8520
rect 120712 8517 120724 8551
rect 120758 8548 120770 8551
rect 122392 8548 122420 8579
rect 120758 8520 122420 8548
rect 120758 8517 120770 8520
rect 120712 8511 120770 8517
rect 122475 8480 122503 8588
rect 130286 8548 130292 8560
rect 122944 8520 130292 8548
rect 120644 8452 122503 8480
rect 122561 8483 122619 8489
rect 122561 8449 122573 8483
rect 122607 8480 122619 8483
rect 122834 8480 122840 8492
rect 122607 8452 122840 8480
rect 122607 8449 122619 8452
rect 122561 8443 122619 8449
rect 122834 8440 122840 8452
rect 122892 8440 122898 8492
rect 117498 8412 117504 8424
rect 117240 8384 117504 8412
rect 117498 8372 117504 8384
rect 117556 8372 117562 8424
rect 117590 8372 117596 8424
rect 117648 8412 117654 8424
rect 117961 8415 118019 8421
rect 117961 8412 117973 8415
rect 117648 8384 117973 8412
rect 117648 8372 117654 8384
rect 117961 8381 117973 8384
rect 118007 8381 118019 8415
rect 118326 8412 118332 8424
rect 118287 8384 118332 8412
rect 117961 8375 118019 8381
rect 118326 8372 118332 8384
rect 118384 8372 118390 8424
rect 118510 8372 118516 8424
rect 118568 8412 118574 8424
rect 118789 8415 118847 8421
rect 118789 8412 118801 8415
rect 118568 8384 118801 8412
rect 118568 8372 118574 8384
rect 118789 8381 118801 8384
rect 118835 8381 118847 8415
rect 119154 8412 119160 8424
rect 119115 8384 119160 8412
rect 118789 8375 118847 8381
rect 119154 8372 119160 8384
rect 119212 8412 119218 8424
rect 119893 8415 119951 8421
rect 119893 8412 119905 8415
rect 119212 8384 119905 8412
rect 119212 8372 119218 8384
rect 119893 8381 119905 8384
rect 119939 8412 119951 8415
rect 119982 8412 119988 8424
rect 119939 8384 119988 8412
rect 119939 8381 119951 8384
rect 119893 8375 119951 8381
rect 119982 8372 119988 8384
rect 120040 8372 120046 8424
rect 120445 8415 120503 8421
rect 120445 8381 120457 8415
rect 120491 8381 120503 8415
rect 122944 8412 122972 8520
rect 130286 8508 130292 8520
rect 130344 8508 130350 8560
rect 123294 8489 123300 8492
rect 123288 8480 123300 8489
rect 123255 8452 123300 8480
rect 123288 8443 123300 8452
rect 123294 8440 123300 8443
rect 123352 8440 123358 8492
rect 123570 8440 123576 8492
rect 123628 8480 123634 8492
rect 126517 8483 126575 8489
rect 126517 8480 126529 8483
rect 123628 8452 126529 8480
rect 123628 8440 123634 8452
rect 126517 8449 126529 8452
rect 126563 8449 126575 8483
rect 126517 8443 126575 8449
rect 126606 8440 126612 8492
rect 126664 8480 126670 8492
rect 127250 8480 127256 8492
rect 126664 8452 127256 8480
rect 126664 8440 126670 8452
rect 127250 8440 127256 8452
rect 127308 8440 127314 8492
rect 127342 8440 127348 8492
rect 127400 8480 127406 8492
rect 128541 8483 128599 8489
rect 128541 8480 128553 8483
rect 127400 8452 128553 8480
rect 127400 8440 127406 8452
rect 128541 8449 128553 8452
rect 128587 8449 128599 8483
rect 130381 8483 130439 8489
rect 128541 8443 128599 8449
rect 128648 8452 128952 8480
rect 120445 8375 120503 8381
rect 121840 8384 122972 8412
rect 84013 8347 84071 8353
rect 84013 8313 84025 8347
rect 84059 8313 84071 8347
rect 84013 8307 84071 8313
rect 86494 8304 86500 8356
rect 86552 8344 86558 8356
rect 86773 8347 86831 8353
rect 86773 8344 86785 8347
rect 86552 8316 86785 8344
rect 86552 8304 86558 8316
rect 86773 8313 86785 8316
rect 86819 8313 86831 8347
rect 86773 8307 86831 8313
rect 92198 8304 92204 8356
rect 92256 8344 92262 8356
rect 93302 8344 93308 8356
rect 92256 8316 92796 8344
rect 93263 8316 93308 8344
rect 92256 8304 92262 8316
rect 59078 8276 59084 8288
rect 58084 8248 59084 8276
rect 54628 8236 54634 8248
rect 59078 8236 59084 8248
rect 59136 8236 59142 8288
rect 59998 8236 60004 8288
rect 60056 8276 60062 8288
rect 60461 8279 60519 8285
rect 60461 8276 60473 8279
rect 60056 8248 60473 8276
rect 60056 8236 60062 8248
rect 60461 8245 60473 8248
rect 60507 8245 60519 8279
rect 60461 8239 60519 8245
rect 65242 8236 65248 8288
rect 65300 8276 65306 8288
rect 65521 8279 65579 8285
rect 65521 8276 65533 8279
rect 65300 8248 65533 8276
rect 65300 8236 65306 8248
rect 65521 8245 65533 8248
rect 65567 8245 65579 8279
rect 74350 8276 74356 8288
rect 74311 8248 74356 8276
rect 65521 8239 65579 8245
rect 74350 8236 74356 8248
rect 74408 8236 74414 8288
rect 75086 8236 75092 8288
rect 75144 8276 75150 8288
rect 83918 8276 83924 8288
rect 75144 8248 83924 8276
rect 75144 8236 75150 8248
rect 83918 8236 83924 8248
rect 83976 8236 83982 8288
rect 84102 8236 84108 8288
rect 84160 8276 84166 8288
rect 90726 8276 90732 8288
rect 84160 8248 90732 8276
rect 84160 8236 84166 8248
rect 90726 8236 90732 8248
rect 90784 8236 90790 8288
rect 90818 8236 90824 8288
rect 90876 8276 90882 8288
rect 92382 8276 92388 8288
rect 90876 8248 92388 8276
rect 90876 8236 90882 8248
rect 92382 8236 92388 8248
rect 92440 8236 92446 8288
rect 92768 8285 92796 8316
rect 93302 8304 93308 8316
rect 93360 8304 93366 8356
rect 94501 8347 94559 8353
rect 94501 8313 94513 8347
rect 94547 8344 94559 8347
rect 95326 8344 95332 8356
rect 94547 8316 95332 8344
rect 94547 8313 94559 8316
rect 94501 8307 94559 8313
rect 95326 8304 95332 8316
rect 95384 8304 95390 8356
rect 95418 8304 95424 8356
rect 95476 8344 95482 8356
rect 101674 8344 101680 8356
rect 95476 8316 101680 8344
rect 95476 8304 95482 8316
rect 101674 8304 101680 8316
rect 101732 8304 101738 8356
rect 104250 8304 104256 8356
rect 104308 8344 104314 8356
rect 108117 8347 108175 8353
rect 108117 8344 108129 8347
rect 104308 8316 108129 8344
rect 104308 8304 104314 8316
rect 108117 8313 108129 8316
rect 108163 8313 108175 8347
rect 108117 8307 108175 8313
rect 110969 8347 111027 8353
rect 110969 8313 110981 8347
rect 111015 8344 111027 8347
rect 112806 8344 112812 8356
rect 111015 8316 112812 8344
rect 111015 8313 111027 8316
rect 110969 8307 111027 8313
rect 112806 8304 112812 8316
rect 112864 8304 112870 8356
rect 115845 8347 115903 8353
rect 115845 8313 115857 8347
rect 115891 8344 115903 8347
rect 115891 8316 117728 8344
rect 115891 8313 115903 8316
rect 115845 8307 115903 8313
rect 92753 8279 92811 8285
rect 92753 8245 92765 8279
rect 92799 8276 92811 8279
rect 97534 8276 97540 8288
rect 92799 8248 97540 8276
rect 92799 8245 92811 8248
rect 92753 8239 92811 8245
rect 97534 8236 97540 8248
rect 97592 8236 97598 8288
rect 98270 8236 98276 8288
rect 98328 8276 98334 8288
rect 101858 8276 101864 8288
rect 98328 8248 101864 8276
rect 98328 8236 98334 8248
rect 101858 8236 101864 8248
rect 101916 8236 101922 8288
rect 108666 8236 108672 8288
rect 108724 8276 108730 8288
rect 108761 8279 108819 8285
rect 108761 8276 108773 8279
rect 108724 8248 108773 8276
rect 108724 8236 108730 8248
rect 108761 8245 108773 8248
rect 108807 8245 108819 8279
rect 108761 8239 108819 8245
rect 112070 8236 112076 8288
rect 112128 8276 112134 8288
rect 115934 8276 115940 8288
rect 112128 8248 115940 8276
rect 112128 8236 112134 8248
rect 115934 8236 115940 8248
rect 115992 8236 115998 8288
rect 116026 8236 116032 8288
rect 116084 8276 116090 8288
rect 116857 8279 116915 8285
rect 116857 8276 116869 8279
rect 116084 8248 116869 8276
rect 116084 8236 116090 8248
rect 116857 8245 116869 8248
rect 116903 8276 116915 8279
rect 117498 8276 117504 8288
rect 116903 8248 117504 8276
rect 116903 8245 116915 8248
rect 116857 8239 116915 8245
rect 117498 8236 117504 8248
rect 117556 8236 117562 8288
rect 117700 8276 117728 8316
rect 119430 8304 119436 8356
rect 119488 8344 119494 8356
rect 120460 8344 120488 8375
rect 121840 8353 121868 8384
rect 123018 8372 123024 8424
rect 123076 8412 123082 8424
rect 125134 8412 125140 8424
rect 123076 8384 123121 8412
rect 124048 8384 125140 8412
rect 123076 8372 123082 8384
rect 119488 8316 120488 8344
rect 119488 8304 119494 8316
rect 120166 8276 120172 8288
rect 117700 8248 120172 8276
rect 120166 8236 120172 8248
rect 120224 8236 120230 8288
rect 120460 8276 120488 8316
rect 121825 8347 121883 8353
rect 121825 8313 121837 8347
rect 121871 8313 121883 8347
rect 121825 8307 121883 8313
rect 122006 8304 122012 8356
rect 122064 8344 122070 8356
rect 123036 8344 123064 8372
rect 124048 8344 124076 8384
rect 125134 8372 125140 8384
rect 125192 8372 125198 8424
rect 126146 8372 126152 8424
rect 126204 8412 126210 8424
rect 126624 8412 126652 8440
rect 126790 8412 126796 8424
rect 126204 8384 126652 8412
rect 126751 8384 126796 8412
rect 126204 8372 126210 8384
rect 126790 8372 126796 8384
rect 126848 8372 126854 8424
rect 127618 8372 127624 8424
rect 127676 8412 127682 8424
rect 128648 8412 128676 8452
rect 127676 8384 128676 8412
rect 128817 8415 128875 8421
rect 127676 8372 127682 8384
rect 128817 8381 128829 8415
rect 128863 8381 128875 8415
rect 128924 8412 128952 8452
rect 130381 8449 130393 8483
rect 130427 8449 130439 8483
rect 130488 8480 130516 8588
rect 130565 8585 130577 8619
rect 130611 8585 130623 8619
rect 130565 8579 130623 8585
rect 130580 8548 130608 8579
rect 131298 8576 131304 8628
rect 131356 8616 131362 8628
rect 131577 8619 131635 8625
rect 131577 8616 131589 8619
rect 131356 8588 131589 8616
rect 131356 8576 131362 8588
rect 131577 8585 131589 8588
rect 131623 8585 131635 8619
rect 131577 8579 131635 8585
rect 131666 8576 131672 8628
rect 131724 8616 131730 8628
rect 132310 8616 132316 8628
rect 131724 8588 132316 8616
rect 131724 8576 131730 8588
rect 132310 8576 132316 8588
rect 132368 8576 132374 8628
rect 132770 8576 132776 8628
rect 132828 8616 132834 8628
rect 135717 8619 135775 8625
rect 135717 8616 135729 8619
rect 132828 8588 135729 8616
rect 132828 8576 132834 8588
rect 135717 8585 135729 8588
rect 135763 8616 135775 8619
rect 143350 8616 143356 8628
rect 135763 8588 143356 8616
rect 135763 8585 135775 8588
rect 135717 8579 135775 8585
rect 143350 8576 143356 8588
rect 143408 8576 143414 8628
rect 144914 8616 144920 8628
rect 143552 8588 144920 8616
rect 133662 8551 133720 8557
rect 133662 8548 133674 8551
rect 130580 8520 133674 8548
rect 133662 8517 133674 8520
rect 133708 8517 133720 8551
rect 143552 8548 143580 8588
rect 144914 8576 144920 8588
rect 144972 8576 144978 8628
rect 145009 8619 145067 8625
rect 145009 8585 145021 8619
rect 145055 8616 145067 8619
rect 146018 8616 146024 8628
rect 145055 8588 146024 8616
rect 145055 8585 145067 8588
rect 145009 8579 145067 8585
rect 146018 8576 146024 8588
rect 146076 8576 146082 8628
rect 147766 8576 147772 8628
rect 147824 8616 147830 8628
rect 149701 8619 149759 8625
rect 147824 8588 149652 8616
rect 147824 8576 147830 8588
rect 148226 8548 148232 8560
rect 133662 8511 133720 8517
rect 135732 8520 141188 8548
rect 135732 8492 135760 8520
rect 132402 8480 132408 8492
rect 130488 8452 132408 8480
rect 130381 8443 130439 8449
rect 130396 8412 130424 8443
rect 132402 8440 132408 8452
rect 132460 8440 132466 8492
rect 132701 8483 132759 8489
rect 132701 8449 132713 8483
rect 132747 8480 132759 8483
rect 135346 8480 135352 8492
rect 132747 8452 135352 8480
rect 132747 8449 132759 8452
rect 132701 8443 132759 8449
rect 135346 8440 135352 8452
rect 135404 8440 135410 8492
rect 135714 8440 135720 8492
rect 135772 8440 135778 8492
rect 137465 8483 137523 8489
rect 137465 8449 137477 8483
rect 137511 8480 137523 8483
rect 137830 8480 137836 8492
rect 137511 8452 137836 8480
rect 137511 8449 137523 8452
rect 137465 8443 137523 8449
rect 137830 8440 137836 8452
rect 137888 8440 137894 8492
rect 138198 8440 138204 8492
rect 138256 8480 138262 8492
rect 140501 8483 140559 8489
rect 138256 8452 139992 8480
rect 138256 8440 138262 8452
rect 128924 8384 130424 8412
rect 132957 8415 133015 8421
rect 128817 8375 128875 8381
rect 132957 8381 132969 8415
rect 133003 8412 133015 8415
rect 133138 8412 133144 8424
rect 133003 8384 133144 8412
rect 133003 8381 133015 8384
rect 132957 8375 133015 8381
rect 122064 8316 123064 8344
rect 123956 8316 124076 8344
rect 124401 8347 124459 8353
rect 122064 8304 122070 8316
rect 121454 8276 121460 8288
rect 120460 8248 121460 8276
rect 121454 8236 121460 8248
rect 121512 8236 121518 8288
rect 123294 8236 123300 8288
rect 123352 8276 123358 8288
rect 123956 8276 123984 8316
rect 124401 8313 124413 8347
rect 124447 8344 124459 8347
rect 127710 8344 127716 8356
rect 124447 8316 127716 8344
rect 124447 8313 124459 8316
rect 124401 8307 124459 8313
rect 127710 8304 127716 8316
rect 127768 8304 127774 8356
rect 128081 8347 128139 8353
rect 128081 8313 128093 8347
rect 128127 8344 128139 8347
rect 128354 8344 128360 8356
rect 128127 8316 128360 8344
rect 128127 8313 128139 8316
rect 128081 8307 128139 8313
rect 128354 8304 128360 8316
rect 128412 8304 128418 8356
rect 128446 8304 128452 8356
rect 128504 8344 128510 8356
rect 128832 8344 128860 8375
rect 133138 8372 133144 8384
rect 133196 8372 133202 8424
rect 133417 8415 133475 8421
rect 133417 8381 133429 8415
rect 133463 8381 133475 8415
rect 133417 8375 133475 8381
rect 128504 8316 128860 8344
rect 128504 8304 128510 8316
rect 130286 8304 130292 8356
rect 130344 8344 130350 8356
rect 131942 8344 131948 8356
rect 130344 8316 131948 8344
rect 130344 8304 130350 8316
rect 131942 8304 131948 8316
rect 132000 8304 132006 8356
rect 123352 8248 123984 8276
rect 123352 8236 123358 8248
rect 124122 8236 124128 8288
rect 124180 8276 124186 8288
rect 129642 8276 129648 8288
rect 124180 8248 129648 8276
rect 124180 8236 124186 8248
rect 129642 8236 129648 8248
rect 129700 8236 129706 8288
rect 130654 8236 130660 8288
rect 130712 8276 130718 8288
rect 131025 8279 131083 8285
rect 131025 8276 131037 8279
rect 130712 8248 131037 8276
rect 130712 8236 130718 8248
rect 131025 8245 131037 8248
rect 131071 8276 131083 8279
rect 131298 8276 131304 8288
rect 131071 8248 131304 8276
rect 131071 8245 131083 8248
rect 131025 8239 131083 8245
rect 131298 8236 131304 8248
rect 131356 8236 131362 8288
rect 133432 8276 133460 8375
rect 134702 8372 134708 8424
rect 134760 8412 134766 8424
rect 136910 8412 136916 8424
rect 134760 8384 135254 8412
rect 136871 8384 136916 8412
rect 134760 8372 134766 8384
rect 134797 8347 134855 8353
rect 134797 8344 134809 8347
rect 134352 8316 134809 8344
rect 133782 8276 133788 8288
rect 133432 8248 133788 8276
rect 133782 8236 133788 8248
rect 133840 8236 133846 8288
rect 134058 8236 134064 8288
rect 134116 8276 134122 8288
rect 134352 8276 134380 8316
rect 134797 8313 134809 8316
rect 134843 8313 134855 8347
rect 134797 8307 134855 8313
rect 134116 8248 134380 8276
rect 135226 8276 135254 8384
rect 136910 8372 136916 8384
rect 136968 8372 136974 8424
rect 137186 8372 137192 8424
rect 137244 8412 137250 8424
rect 139397 8415 139455 8421
rect 137244 8384 138704 8412
rect 137244 8372 137250 8384
rect 135714 8304 135720 8356
rect 135772 8344 135778 8356
rect 138017 8347 138075 8353
rect 138017 8344 138029 8347
rect 135772 8316 138029 8344
rect 135772 8304 135778 8316
rect 138017 8313 138029 8316
rect 138063 8344 138075 8347
rect 138566 8344 138572 8356
rect 138063 8316 138572 8344
rect 138063 8313 138075 8316
rect 138017 8307 138075 8313
rect 138566 8304 138572 8316
rect 138624 8304 138630 8356
rect 138676 8344 138704 8384
rect 139397 8381 139409 8415
rect 139443 8412 139455 8415
rect 139854 8412 139860 8424
rect 139443 8384 139860 8412
rect 139443 8381 139455 8384
rect 139397 8375 139455 8381
rect 139854 8372 139860 8384
rect 139912 8372 139918 8424
rect 139964 8421 139992 8452
rect 140501 8449 140513 8483
rect 140547 8480 140559 8483
rect 140547 8452 141096 8480
rect 140547 8449 140559 8452
rect 140501 8443 140559 8449
rect 139949 8415 140007 8421
rect 139949 8381 139961 8415
rect 139995 8412 140007 8415
rect 140958 8412 140964 8424
rect 139995 8384 140964 8412
rect 139995 8381 140007 8384
rect 139949 8375 140007 8381
rect 140958 8372 140964 8384
rect 141016 8372 141022 8424
rect 140682 8344 140688 8356
rect 138676 8316 140544 8344
rect 140643 8316 140688 8344
rect 136361 8279 136419 8285
rect 136361 8276 136373 8279
rect 135226 8248 136373 8276
rect 134116 8236 134122 8248
rect 136361 8245 136373 8248
rect 136407 8276 136419 8279
rect 137462 8276 137468 8288
rect 136407 8248 137468 8276
rect 136407 8245 136419 8248
rect 136361 8239 136419 8245
rect 137462 8236 137468 8248
rect 137520 8236 137526 8288
rect 138658 8236 138664 8288
rect 138716 8276 138722 8288
rect 139762 8276 139768 8288
rect 138716 8248 139768 8276
rect 138716 8236 138722 8248
rect 139762 8236 139768 8248
rect 139820 8236 139826 8288
rect 140516 8276 140544 8316
rect 140682 8304 140688 8316
rect 140740 8304 140746 8356
rect 140590 8276 140596 8288
rect 140516 8248 140596 8276
rect 140590 8236 140596 8248
rect 140648 8236 140654 8288
rect 141068 8276 141096 8452
rect 141160 8353 141188 8520
rect 141436 8520 143580 8548
rect 143644 8520 148232 8548
rect 141326 8480 141332 8492
rect 141287 8452 141332 8480
rect 141326 8440 141332 8452
rect 141384 8440 141390 8492
rect 141436 8412 141464 8520
rect 141510 8440 141516 8492
rect 141568 8480 141574 8492
rect 142902 8483 142960 8489
rect 142902 8480 142914 8483
rect 141568 8452 142914 8480
rect 141568 8440 141574 8452
rect 142902 8449 142914 8452
rect 142948 8449 142960 8483
rect 142902 8443 142960 8449
rect 143074 8440 143080 8492
rect 143132 8480 143138 8492
rect 143169 8483 143227 8489
rect 143169 8480 143181 8483
rect 143132 8452 143181 8480
rect 143132 8440 143138 8452
rect 143169 8449 143181 8452
rect 143215 8480 143227 8483
rect 143258 8480 143264 8492
rect 143215 8452 143264 8480
rect 143215 8449 143227 8452
rect 143169 8443 143227 8449
rect 143258 8440 143264 8452
rect 143316 8480 143322 8492
rect 143644 8489 143672 8520
rect 143902 8489 143908 8492
rect 143629 8483 143687 8489
rect 143629 8480 143641 8483
rect 143316 8452 143641 8480
rect 143316 8440 143322 8452
rect 143629 8449 143641 8452
rect 143675 8449 143687 8483
rect 143896 8480 143908 8489
rect 143863 8452 143908 8480
rect 143629 8443 143687 8449
rect 143896 8443 143908 8452
rect 143902 8440 143908 8443
rect 143960 8440 143966 8492
rect 145650 8480 145656 8492
rect 145611 8452 145656 8480
rect 145650 8440 145656 8452
rect 145708 8440 145714 8492
rect 145920 8483 145978 8489
rect 145920 8449 145932 8483
rect 145966 8480 145978 8483
rect 147398 8480 147404 8492
rect 145966 8452 147404 8480
rect 145966 8449 145978 8452
rect 145920 8443 145978 8449
rect 147398 8440 147404 8452
rect 147456 8440 147462 8492
rect 147508 8489 147536 8520
rect 148226 8508 148232 8520
rect 148284 8508 148290 8560
rect 148318 8508 148324 8560
rect 148376 8548 148382 8560
rect 148686 8548 148692 8560
rect 148376 8520 148692 8548
rect 148376 8508 148382 8520
rect 148686 8508 148692 8520
rect 148744 8508 148750 8560
rect 149624 8548 149652 8588
rect 149701 8585 149713 8619
rect 149747 8616 149759 8619
rect 149882 8616 149888 8628
rect 149747 8588 149888 8616
rect 149747 8585 149759 8588
rect 149701 8579 149759 8585
rect 149882 8576 149888 8588
rect 149940 8576 149946 8628
rect 150802 8616 150808 8628
rect 150763 8588 150808 8616
rect 150802 8576 150808 8588
rect 150860 8576 150866 8628
rect 150894 8576 150900 8628
rect 150952 8616 150958 8628
rect 151078 8616 151084 8628
rect 150952 8588 151084 8616
rect 150952 8576 150958 8588
rect 151078 8576 151084 8588
rect 151136 8616 151142 8628
rect 155310 8616 155316 8628
rect 151136 8588 154344 8616
rect 155271 8588 155316 8616
rect 151136 8576 151142 8588
rect 151630 8548 151636 8560
rect 149624 8520 151636 8548
rect 151630 8508 151636 8520
rect 151688 8508 151694 8560
rect 153746 8548 153752 8560
rect 151740 8520 153752 8548
rect 147493 8483 147551 8489
rect 147493 8449 147505 8483
rect 147539 8449 147551 8483
rect 147493 8443 147551 8449
rect 147760 8483 147818 8489
rect 147760 8449 147772 8483
rect 147806 8480 147818 8483
rect 147806 8452 149468 8480
rect 147806 8449 147818 8452
rect 147760 8443 147818 8449
rect 141252 8384 141464 8412
rect 141145 8347 141203 8353
rect 141145 8313 141157 8347
rect 141191 8313 141203 8347
rect 141145 8307 141203 8313
rect 141252 8276 141280 8384
rect 141602 8372 141608 8424
rect 141660 8412 141666 8424
rect 141970 8412 141976 8424
rect 141660 8384 141976 8412
rect 141660 8372 141666 8384
rect 141970 8372 141976 8384
rect 142028 8372 142034 8424
rect 144914 8372 144920 8424
rect 144972 8412 144978 8424
rect 145558 8412 145564 8424
rect 144972 8384 145564 8412
rect 144972 8372 144978 8384
rect 145558 8372 145564 8384
rect 145616 8372 145622 8424
rect 147122 8372 147128 8424
rect 147180 8412 147186 8424
rect 147180 8384 147444 8412
rect 147180 8372 147186 8384
rect 147416 8356 147444 8384
rect 148962 8372 148968 8424
rect 149020 8412 149026 8424
rect 149333 8415 149391 8421
rect 149333 8412 149345 8415
rect 149020 8384 149345 8412
rect 149020 8372 149026 8384
rect 149333 8381 149345 8384
rect 149379 8381 149391 8415
rect 149440 8412 149468 8452
rect 149514 8440 149520 8492
rect 149572 8480 149578 8492
rect 149572 8452 149617 8480
rect 149572 8440 149578 8452
rect 149882 8440 149888 8492
rect 149940 8480 149946 8492
rect 150989 8483 151047 8489
rect 150989 8480 151001 8483
rect 149940 8452 151001 8480
rect 149940 8440 149946 8452
rect 150989 8449 151001 8452
rect 151035 8449 151047 8483
rect 150989 8443 151047 8449
rect 151170 8440 151176 8492
rect 151228 8480 151234 8492
rect 151740 8480 151768 8520
rect 153746 8508 153752 8520
rect 153804 8548 153810 8560
rect 154206 8548 154212 8560
rect 153804 8520 153884 8548
rect 153804 8508 153810 8520
rect 151228 8452 151768 8480
rect 151228 8440 151234 8452
rect 151814 8440 151820 8492
rect 151872 8480 151878 8492
rect 152826 8480 152832 8492
rect 151872 8452 152832 8480
rect 151872 8440 151878 8452
rect 152826 8440 152832 8452
rect 152884 8440 152890 8492
rect 153856 8489 153884 8520
rect 153948 8520 154212 8548
rect 153841 8483 153899 8489
rect 153841 8449 153853 8483
rect 153887 8449 153899 8483
rect 153841 8443 153899 8449
rect 149440 8384 150112 8412
rect 149333 8375 149391 8381
rect 141786 8344 141792 8356
rect 141747 8316 141792 8344
rect 141786 8304 141792 8316
rect 141844 8304 141850 8356
rect 147033 8347 147091 8353
rect 147033 8313 147045 8347
rect 147079 8344 147091 8347
rect 147214 8344 147220 8356
rect 147079 8316 147220 8344
rect 147079 8313 147091 8316
rect 147033 8307 147091 8313
rect 147214 8304 147220 8316
rect 147272 8304 147278 8356
rect 147398 8304 147404 8356
rect 147456 8304 147462 8356
rect 148873 8347 148931 8353
rect 148873 8313 148885 8347
rect 148919 8344 148931 8347
rect 149054 8344 149060 8356
rect 148919 8316 149060 8344
rect 148919 8313 148931 8316
rect 148873 8307 148931 8313
rect 149054 8304 149060 8316
rect 149112 8304 149118 8356
rect 149348 8344 149376 8375
rect 150084 8344 150112 8384
rect 150158 8372 150164 8424
rect 150216 8412 150222 8424
rect 150894 8412 150900 8424
rect 150216 8384 150900 8412
rect 150216 8372 150222 8384
rect 150894 8372 150900 8384
rect 150952 8372 150958 8424
rect 151998 8412 152004 8424
rect 151959 8384 152004 8412
rect 151998 8372 152004 8384
rect 152056 8372 152062 8424
rect 152274 8412 152280 8424
rect 152235 8384 152280 8412
rect 152274 8372 152280 8384
rect 152332 8372 152338 8424
rect 153010 8344 153016 8356
rect 149348 8316 149560 8344
rect 150084 8316 153016 8344
rect 141068 8248 141280 8276
rect 142062 8236 142068 8288
rect 142120 8276 142126 8288
rect 144914 8276 144920 8288
rect 142120 8248 144920 8276
rect 142120 8236 142126 8248
rect 144914 8236 144920 8248
rect 144972 8236 144978 8288
rect 146018 8236 146024 8288
rect 146076 8276 146082 8288
rect 149422 8276 149428 8288
rect 146076 8248 149428 8276
rect 146076 8236 146082 8248
rect 149422 8236 149428 8248
rect 149480 8236 149486 8288
rect 149532 8276 149560 8316
rect 153010 8304 153016 8316
rect 153068 8304 153074 8356
rect 150161 8279 150219 8285
rect 150161 8276 150173 8279
rect 149532 8248 150173 8276
rect 150161 8245 150173 8248
rect 150207 8245 150219 8279
rect 150161 8239 150219 8245
rect 151078 8236 151084 8288
rect 151136 8276 151142 8288
rect 152921 8279 152979 8285
rect 152921 8276 152933 8279
rect 151136 8248 152933 8276
rect 151136 8236 151142 8248
rect 152921 8245 152933 8248
rect 152967 8276 152979 8279
rect 153470 8276 153476 8288
rect 152967 8248 153476 8276
rect 152967 8245 152979 8248
rect 152921 8239 152979 8245
rect 153470 8236 153476 8248
rect 153528 8236 153534 8288
rect 153654 8276 153660 8288
rect 153615 8248 153660 8276
rect 153654 8236 153660 8248
rect 153712 8236 153718 8288
rect 153948 8276 153976 8520
rect 154206 8508 154212 8520
rect 154264 8508 154270 8560
rect 154316 8548 154344 8588
rect 155310 8576 155316 8588
rect 155368 8576 155374 8628
rect 155954 8576 155960 8628
rect 156012 8616 156018 8628
rect 156782 8616 156788 8628
rect 156012 8588 156788 8616
rect 156012 8576 156018 8588
rect 156782 8576 156788 8588
rect 156840 8576 156846 8628
rect 156966 8576 156972 8628
rect 157024 8576 157030 8628
rect 156984 8548 157012 8576
rect 154316 8520 156184 8548
rect 154298 8440 154304 8492
rect 154356 8480 154362 8492
rect 156156 8489 156184 8520
rect 156340 8520 157012 8548
rect 156340 8489 156368 8520
rect 154669 8483 154727 8489
rect 154669 8480 154681 8483
rect 154356 8452 154681 8480
rect 154356 8440 154362 8452
rect 154669 8449 154681 8452
rect 154715 8449 154727 8483
rect 154669 8443 154727 8449
rect 156141 8483 156199 8489
rect 156141 8449 156153 8483
rect 156187 8449 156199 8483
rect 156141 8443 156199 8449
rect 156325 8483 156383 8489
rect 156325 8449 156337 8483
rect 156371 8449 156383 8483
rect 156782 8480 156788 8492
rect 156743 8452 156788 8480
rect 156325 8443 156383 8449
rect 154025 8415 154083 8421
rect 154025 8381 154037 8415
rect 154071 8412 154083 8415
rect 154206 8412 154212 8424
rect 154071 8384 154212 8412
rect 154071 8381 154083 8384
rect 154025 8375 154083 8381
rect 154206 8372 154212 8384
rect 154264 8412 154270 8424
rect 154264 8384 154712 8412
rect 154264 8372 154270 8384
rect 154482 8344 154488 8356
rect 154443 8316 154488 8344
rect 154482 8304 154488 8316
rect 154540 8304 154546 8356
rect 154684 8344 154712 8384
rect 154758 8372 154764 8424
rect 154816 8412 154822 8424
rect 154853 8415 154911 8421
rect 154853 8412 154865 8415
rect 154816 8384 154865 8412
rect 154816 8372 154822 8384
rect 154853 8381 154865 8384
rect 154899 8412 154911 8415
rect 155770 8412 155776 8424
rect 154899 8384 155776 8412
rect 154899 8381 154911 8384
rect 154853 8375 154911 8381
rect 155770 8372 155776 8384
rect 155828 8412 155834 8424
rect 156340 8412 156368 8443
rect 156782 8440 156788 8452
rect 156840 8440 156846 8492
rect 156966 8480 156972 8492
rect 156927 8452 156972 8480
rect 156966 8440 156972 8452
rect 157024 8440 157030 8492
rect 158070 8480 158076 8492
rect 158031 8452 158076 8480
rect 158070 8440 158076 8452
rect 158128 8440 158134 8492
rect 155828 8384 156368 8412
rect 155828 8372 155834 8384
rect 155954 8344 155960 8356
rect 154684 8316 155816 8344
rect 155915 8316 155960 8344
rect 154298 8276 154304 8288
rect 153948 8248 154304 8276
rect 154298 8236 154304 8248
rect 154356 8276 154362 8288
rect 155402 8276 155408 8288
rect 154356 8248 155408 8276
rect 154356 8236 154362 8248
rect 155402 8236 155408 8248
rect 155460 8236 155466 8288
rect 155788 8276 155816 8316
rect 155954 8304 155960 8316
rect 156012 8304 156018 8356
rect 156138 8344 156144 8356
rect 156064 8316 156144 8344
rect 156064 8276 156092 8316
rect 156138 8304 156144 8316
rect 156196 8304 156202 8356
rect 157153 8347 157211 8353
rect 157153 8313 157165 8347
rect 157199 8344 157211 8347
rect 157334 8344 157340 8356
rect 157199 8316 157340 8344
rect 157199 8313 157211 8316
rect 157153 8307 157211 8313
rect 157334 8304 157340 8316
rect 157392 8304 157398 8356
rect 157518 8304 157524 8356
rect 157576 8344 157582 8356
rect 158070 8344 158076 8356
rect 157576 8316 158076 8344
rect 157576 8304 157582 8316
rect 158070 8304 158076 8316
rect 158128 8304 158134 8356
rect 158254 8344 158260 8356
rect 158215 8316 158260 8344
rect 158254 8304 158260 8316
rect 158312 8304 158318 8356
rect 155788 8248 156092 8276
rect 1104 8186 158884 8208
rect 1104 8134 20672 8186
rect 20724 8134 20736 8186
rect 20788 8134 20800 8186
rect 20852 8134 20864 8186
rect 20916 8134 20928 8186
rect 20980 8134 60117 8186
rect 60169 8134 60181 8186
rect 60233 8134 60245 8186
rect 60297 8134 60309 8186
rect 60361 8134 60373 8186
rect 60425 8134 99562 8186
rect 99614 8134 99626 8186
rect 99678 8134 99690 8186
rect 99742 8134 99754 8186
rect 99806 8134 99818 8186
rect 99870 8134 139007 8186
rect 139059 8134 139071 8186
rect 139123 8134 139135 8186
rect 139187 8134 139199 8186
rect 139251 8134 139263 8186
rect 139315 8134 158884 8186
rect 1104 8112 158884 8134
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 10686 8072 10692 8084
rect 6411 8044 10692 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 12894 8072 12900 8084
rect 12807 8044 12900 8072
rect 12894 8032 12900 8044
rect 12952 8072 12958 8084
rect 13722 8072 13728 8084
rect 12952 8044 13728 8072
rect 12952 8032 12958 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 14332 8044 14381 8072
rect 14332 8032 14338 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 17862 8072 17868 8084
rect 15335 8044 17868 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18598 8072 18604 8084
rect 18559 8044 18604 8072
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 21545 8075 21603 8081
rect 21545 8041 21557 8075
rect 21591 8072 21603 8075
rect 22186 8072 22192 8084
rect 21591 8044 22192 8072
rect 21591 8041 21603 8044
rect 21545 8035 21603 8041
rect 22186 8032 22192 8044
rect 22244 8072 22250 8084
rect 23382 8072 23388 8084
rect 22244 8044 23388 8072
rect 22244 8032 22250 8044
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 26053 8075 26111 8081
rect 26053 8041 26065 8075
rect 26099 8072 26111 8075
rect 27246 8072 27252 8084
rect 26099 8044 27252 8072
rect 26099 8041 26111 8044
rect 26053 8035 26111 8041
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 31018 8072 31024 8084
rect 30979 8044 31024 8072
rect 31018 8032 31024 8044
rect 31076 8032 31082 8084
rect 31570 8072 31576 8084
rect 31531 8044 31576 8072
rect 31570 8032 31576 8044
rect 31628 8032 31634 8084
rect 31726 8044 35480 8072
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 8004 5779 8007
rect 5767 7976 17172 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 5442 7936 5448 7948
rect 5000 7908 5448 7936
rect 5000 7877 5028 7908
rect 5442 7896 5448 7908
rect 5500 7936 5506 7948
rect 5736 7936 5764 7967
rect 5500 7908 5764 7936
rect 12345 7939 12403 7945
rect 5500 7896 5506 7908
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12391 7908 14872 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 14844 7880 14872 7908
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 15896 7908 16896 7936
rect 15896 7896 15902 7908
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5626 7868 5632 7880
rect 5215 7840 5632 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5626 7828 5632 7840
rect 5684 7868 5690 7880
rect 5994 7868 6000 7880
rect 5684 7840 6000 7868
rect 5684 7828 5690 7840
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 6181 7831 6239 7837
rect 6196 7800 6224 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14884 7840 14933 7868
rect 14884 7828 14890 7840
rect 14921 7837 14933 7840
rect 14967 7868 14979 7871
rect 15010 7868 15016 7880
rect 14967 7840 15016 7868
rect 14967 7837 14979 7840
rect 14921 7831 14979 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 16114 7868 16120 7880
rect 16075 7840 16120 7868
rect 15105 7831 15163 7837
rect 6638 7800 6644 7812
rect 6196 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7800 6702 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6696 7772 7021 7800
rect 6696 7760 6702 7772
rect 7009 7769 7021 7772
rect 7055 7800 7067 7803
rect 8386 7800 8392 7812
rect 7055 7772 8392 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 8386 7760 8392 7772
rect 8444 7800 8450 7812
rect 8444 7772 13676 7800
rect 8444 7760 8450 7772
rect 4798 7732 4804 7744
rect 4759 7704 4804 7732
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 13354 7732 13360 7744
rect 13315 7704 13360 7732
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13648 7732 13676 7772
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 15120 7800 15148 7831
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 13780 7772 15148 7800
rect 13780 7760 13786 7772
rect 15470 7760 15476 7812
rect 15528 7800 15534 7812
rect 16868 7800 16896 7908
rect 17144 7868 17172 7976
rect 24210 7964 24216 8016
rect 24268 8004 24274 8016
rect 31726 8004 31754 8044
rect 32490 8004 32496 8016
rect 24268 7976 31754 8004
rect 32403 7976 32496 8004
rect 24268 7964 24274 7976
rect 32490 7964 32496 7976
rect 32548 8004 32554 8016
rect 33226 8004 33232 8016
rect 32548 7976 33232 8004
rect 32548 7964 32554 7976
rect 33226 7964 33232 7976
rect 33284 7964 33290 8016
rect 18966 7936 18972 7948
rect 18064 7908 18972 7936
rect 18064 7868 18092 7908
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 35452 7936 35480 8044
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 36173 8075 36231 8081
rect 36173 8072 36185 8075
rect 35952 8044 36185 8072
rect 35952 8032 35958 8044
rect 36173 8041 36185 8044
rect 36219 8041 36231 8075
rect 36173 8035 36231 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36725 8075 36783 8081
rect 36725 8072 36737 8075
rect 36688 8044 36737 8072
rect 36688 8032 36694 8044
rect 36725 8041 36737 8044
rect 36771 8041 36783 8075
rect 36725 8035 36783 8041
rect 37274 8032 37280 8084
rect 37332 8072 37338 8084
rect 38381 8075 38439 8081
rect 38381 8072 38393 8075
rect 37332 8044 38393 8072
rect 37332 8032 37338 8044
rect 38381 8041 38393 8044
rect 38427 8041 38439 8075
rect 38381 8035 38439 8041
rect 38562 8032 38568 8084
rect 38620 8072 38626 8084
rect 41690 8072 41696 8084
rect 38620 8044 40264 8072
rect 38620 8032 38626 8044
rect 35529 8007 35587 8013
rect 35529 7973 35541 8007
rect 35575 8004 35587 8007
rect 38930 8004 38936 8016
rect 35575 7976 38936 8004
rect 35575 7973 35587 7976
rect 35529 7967 35587 7973
rect 38930 7964 38936 7976
rect 38988 7964 38994 8016
rect 39114 8004 39120 8016
rect 39075 7976 39120 8004
rect 39114 7964 39120 7976
rect 39172 7964 39178 8016
rect 37550 7936 37556 7948
rect 35452 7908 37556 7936
rect 37550 7896 37556 7908
rect 37608 7896 37614 7948
rect 37737 7939 37795 7945
rect 37737 7905 37749 7939
rect 37783 7936 37795 7939
rect 37826 7936 37832 7948
rect 37783 7908 37832 7936
rect 37783 7905 37795 7908
rect 37737 7899 37795 7905
rect 37826 7896 37832 7908
rect 37884 7896 37890 7948
rect 40037 7939 40095 7945
rect 40037 7936 40049 7939
rect 38580 7908 40049 7936
rect 17144 7840 18092 7868
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18196 7840 19012 7868
rect 18196 7828 18202 7840
rect 17874 7803 17932 7809
rect 17874 7800 17886 7803
rect 15528 7772 16804 7800
rect 16868 7772 17886 7800
rect 15528 7760 15534 7772
rect 13998 7732 14004 7744
rect 13648 7704 14004 7732
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 16298 7732 16304 7744
rect 16259 7704 16304 7732
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16776 7741 16804 7772
rect 17874 7769 17886 7772
rect 17920 7769 17932 7803
rect 17874 7763 17932 7769
rect 18984 7744 19012 7840
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22097 7871 22155 7877
rect 22097 7868 22109 7871
rect 21324 7840 22109 7868
rect 21324 7828 21330 7840
rect 22097 7837 22109 7840
rect 22143 7837 22155 7871
rect 25866 7868 25872 7880
rect 25827 7840 25872 7868
rect 22097 7831 22155 7837
rect 25866 7828 25872 7840
rect 25924 7828 25930 7880
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7868 31815 7871
rect 33594 7868 33600 7880
rect 31803 7840 33600 7868
rect 31803 7837 31815 7840
rect 31757 7831 31815 7837
rect 33594 7828 33600 7840
rect 33652 7828 33658 7880
rect 33778 7828 33784 7880
rect 33836 7868 33842 7880
rect 34333 7871 34391 7877
rect 34333 7868 34345 7871
rect 33836 7840 34345 7868
rect 33836 7828 33842 7840
rect 34333 7837 34345 7840
rect 34379 7837 34391 7871
rect 35342 7868 35348 7880
rect 35303 7840 35348 7868
rect 34333 7831 34391 7837
rect 35342 7828 35348 7840
rect 35400 7828 35406 7880
rect 36906 7868 36912 7880
rect 36867 7840 36912 7868
rect 36906 7828 36912 7840
rect 36964 7828 36970 7880
rect 38580 7877 38608 7908
rect 40037 7905 40049 7908
rect 40083 7905 40095 7939
rect 40037 7899 40095 7905
rect 38565 7871 38623 7877
rect 38565 7837 38577 7871
rect 38611 7837 38623 7871
rect 39298 7868 39304 7880
rect 39259 7840 39304 7868
rect 38565 7831 38623 7837
rect 39298 7828 39304 7840
rect 39356 7828 39362 7880
rect 40236 7877 40264 8044
rect 41432 8044 41696 8072
rect 41432 7945 41460 8044
rect 41690 8032 41696 8044
rect 41748 8032 41754 8084
rect 42794 8072 42800 8084
rect 42755 8044 42800 8072
rect 42794 8032 42800 8044
rect 42852 8032 42858 8084
rect 42978 8032 42984 8084
rect 43036 8072 43042 8084
rect 43257 8075 43315 8081
rect 43257 8072 43269 8075
rect 43036 8044 43269 8072
rect 43036 8032 43042 8044
rect 43257 8041 43269 8044
rect 43303 8041 43315 8075
rect 45370 8072 45376 8084
rect 45331 8044 45376 8072
rect 43257 8035 43315 8041
rect 45370 8032 45376 8044
rect 45428 8032 45434 8084
rect 45462 8032 45468 8084
rect 45520 8072 45526 8084
rect 45520 8044 46161 8072
rect 45520 8032 45526 8044
rect 46133 8004 46161 8044
rect 46198 8032 46204 8084
rect 46256 8072 46262 8084
rect 46661 8075 46719 8081
rect 46661 8072 46673 8075
rect 46256 8044 46673 8072
rect 46256 8032 46262 8044
rect 46661 8041 46673 8044
rect 46707 8041 46719 8075
rect 46661 8035 46719 8041
rect 48130 8032 48136 8084
rect 48188 8072 48194 8084
rect 48593 8075 48651 8081
rect 48593 8072 48605 8075
rect 48188 8044 48605 8072
rect 48188 8032 48194 8044
rect 48593 8041 48605 8044
rect 48639 8072 48651 8075
rect 49142 8072 49148 8084
rect 48639 8044 49148 8072
rect 48639 8041 48651 8044
rect 48593 8035 48651 8041
rect 49142 8032 49148 8044
rect 49200 8032 49206 8084
rect 49237 8075 49295 8081
rect 49237 8041 49249 8075
rect 49283 8072 49295 8075
rect 49510 8072 49516 8084
rect 49283 8044 49516 8072
rect 49283 8041 49295 8044
rect 49237 8035 49295 8041
rect 49510 8032 49516 8044
rect 49568 8032 49574 8084
rect 49694 8032 49700 8084
rect 49752 8072 49758 8084
rect 55861 8075 55919 8081
rect 49752 8044 54248 8072
rect 49752 8032 49758 8044
rect 46133 7976 46244 8004
rect 41417 7939 41475 7945
rect 41417 7905 41429 7939
rect 41463 7905 41475 7939
rect 45462 7936 45468 7948
rect 41417 7899 41475 7905
rect 44560 7908 45468 7936
rect 40221 7871 40279 7877
rect 40221 7837 40233 7871
rect 40267 7837 40279 7871
rect 40221 7831 40279 7837
rect 40405 7871 40463 7877
rect 40405 7837 40417 7871
rect 40451 7868 40463 7871
rect 40770 7868 40776 7880
rect 40451 7840 40776 7868
rect 40451 7837 40463 7840
rect 40405 7831 40463 7837
rect 40770 7828 40776 7840
rect 40828 7868 40834 7880
rect 40865 7871 40923 7877
rect 40865 7868 40877 7871
rect 40828 7840 40877 7868
rect 40828 7828 40834 7840
rect 40865 7837 40877 7840
rect 40911 7837 40923 7871
rect 40865 7831 40923 7837
rect 41684 7871 41742 7877
rect 41684 7837 41696 7871
rect 41730 7868 41742 7871
rect 42610 7868 42616 7880
rect 41730 7840 42616 7868
rect 41730 7837 41742 7840
rect 41684 7831 41742 7837
rect 42610 7828 42616 7840
rect 42668 7868 42674 7880
rect 44560 7868 44588 7908
rect 45462 7896 45468 7908
rect 45520 7896 45526 7948
rect 42668 7840 44588 7868
rect 42668 7828 42674 7840
rect 44634 7828 44640 7880
rect 44692 7868 44698 7880
rect 45830 7868 45836 7880
rect 44692 7840 44737 7868
rect 45791 7840 45836 7868
rect 44692 7828 44698 7840
rect 45830 7828 45836 7840
rect 45888 7828 45894 7880
rect 46014 7828 46020 7880
rect 46072 7868 46078 7880
rect 46216 7868 46244 7976
rect 49326 7964 49332 8016
rect 49384 8004 49390 8016
rect 50985 8007 51043 8013
rect 50985 8004 50997 8007
rect 49384 7976 50997 8004
rect 49384 7964 49390 7976
rect 50985 7973 50997 7976
rect 51031 7973 51043 8007
rect 50985 7967 51043 7973
rect 53009 8007 53067 8013
rect 53009 7973 53021 8007
rect 53055 7973 53067 8007
rect 54220 8004 54248 8044
rect 55861 8041 55873 8075
rect 55907 8072 55919 8075
rect 56134 8072 56140 8084
rect 55907 8044 56140 8072
rect 55907 8041 55919 8044
rect 55861 8035 55919 8041
rect 56134 8032 56140 8044
rect 56192 8032 56198 8084
rect 56778 8032 56784 8084
rect 56836 8072 56842 8084
rect 56873 8075 56931 8081
rect 56873 8072 56885 8075
rect 56836 8044 56885 8072
rect 56836 8032 56842 8044
rect 56873 8041 56885 8044
rect 56919 8041 56931 8075
rect 59538 8072 59544 8084
rect 59499 8044 59544 8072
rect 56873 8035 56931 8041
rect 59538 8032 59544 8044
rect 59596 8032 59602 8084
rect 63313 8075 63371 8081
rect 63313 8072 63325 8075
rect 60706 8044 63325 8072
rect 57425 8007 57483 8013
rect 57425 8004 57437 8007
rect 54220 7976 57437 8004
rect 53009 7967 53067 7973
rect 57425 7973 57437 7976
rect 57471 7973 57483 8007
rect 57425 7967 57483 7973
rect 47026 7896 47032 7948
rect 47084 7936 47090 7948
rect 47213 7939 47271 7945
rect 47213 7936 47225 7939
rect 47084 7908 47225 7936
rect 47084 7896 47090 7908
rect 47213 7905 47225 7908
rect 47259 7936 47271 7939
rect 48041 7939 48099 7945
rect 48041 7936 48053 7939
rect 47259 7908 48053 7936
rect 47259 7905 47271 7908
rect 47213 7899 47271 7905
rect 48041 7905 48053 7908
rect 48087 7905 48099 7939
rect 48041 7899 48099 7905
rect 50338 7896 50344 7948
rect 50396 7936 50402 7948
rect 50433 7939 50491 7945
rect 50433 7936 50445 7939
rect 50396 7908 50445 7936
rect 50396 7896 50402 7908
rect 50433 7905 50445 7908
rect 50479 7936 50491 7939
rect 51350 7936 51356 7948
rect 50479 7908 51356 7936
rect 50479 7905 50491 7908
rect 50433 7899 50491 7905
rect 51350 7896 51356 7908
rect 51408 7896 51414 7948
rect 52365 7939 52423 7945
rect 52365 7905 52377 7939
rect 52411 7936 52423 7939
rect 52546 7936 52552 7948
rect 52411 7908 52552 7936
rect 52411 7905 52423 7908
rect 52365 7899 52423 7905
rect 52546 7896 52552 7908
rect 52604 7896 52610 7948
rect 53024 7936 53052 7967
rect 58802 7964 58808 8016
rect 58860 8004 58866 8016
rect 60706 8004 60734 8044
rect 63313 8041 63325 8044
rect 63359 8041 63371 8075
rect 66714 8072 66720 8084
rect 63313 8035 63371 8041
rect 63420 8044 66720 8072
rect 61194 8004 61200 8016
rect 58860 7976 60734 8004
rect 61155 7976 61200 8004
rect 58860 7964 58866 7976
rect 61194 7964 61200 7976
rect 61252 7964 61258 8016
rect 53024 7908 57744 7936
rect 47397 7871 47455 7877
rect 47397 7868 47409 7871
rect 46072 7840 46115 7868
rect 46216 7840 47409 7868
rect 46072 7828 46078 7840
rect 47397 7837 47409 7840
rect 47443 7837 47455 7871
rect 51810 7868 51816 7880
rect 47397 7831 47455 7837
rect 47504 7840 51816 7868
rect 20432 7803 20490 7809
rect 20432 7769 20444 7803
rect 20478 7800 20490 7803
rect 21082 7800 21088 7812
rect 20478 7772 21088 7800
rect 20478 7769 20490 7772
rect 20432 7763 20490 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 27890 7760 27896 7812
rect 27948 7800 27954 7812
rect 32858 7800 32864 7812
rect 27948 7772 32864 7800
rect 27948 7760 27954 7772
rect 32858 7760 32864 7772
rect 32916 7760 32922 7812
rect 34054 7800 34060 7812
rect 34112 7809 34118 7812
rect 34024 7772 34060 7800
rect 34054 7760 34060 7772
rect 34112 7763 34124 7809
rect 34112 7760 34118 7763
rect 36630 7760 36636 7812
rect 36688 7800 36694 7812
rect 39114 7800 39120 7812
rect 36688 7772 39120 7800
rect 36688 7760 36694 7772
rect 39114 7760 39120 7772
rect 39172 7760 39178 7812
rect 39224 7772 41414 7800
rect 16761 7735 16819 7741
rect 16761 7701 16773 7735
rect 16807 7701 16819 7735
rect 16761 7695 16819 7701
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19024 7704 19441 7732
rect 19024 7692 19030 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 23014 7732 23020 7744
rect 22327 7704 23020 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 30558 7692 30564 7744
rect 30616 7732 30622 7744
rect 32490 7732 32496 7744
rect 30616 7704 32496 7732
rect 30616 7692 30622 7704
rect 32490 7692 32496 7704
rect 32548 7692 32554 7744
rect 32950 7732 32956 7744
rect 32911 7704 32956 7732
rect 32950 7692 32956 7704
rect 33008 7692 33014 7744
rect 33962 7692 33968 7744
rect 34020 7732 34026 7744
rect 39224 7732 39252 7772
rect 34020 7704 39252 7732
rect 41386 7732 41414 7772
rect 42886 7760 42892 7812
rect 42944 7800 42950 7812
rect 44370 7803 44428 7809
rect 44370 7800 44382 7803
rect 42944 7772 44382 7800
rect 42944 7760 42950 7772
rect 44370 7769 44382 7772
rect 44416 7769 44428 7803
rect 47504 7800 47532 7840
rect 51810 7828 51816 7840
rect 51868 7828 51874 7880
rect 52454 7828 52460 7880
rect 52512 7868 52518 7880
rect 52825 7871 52883 7877
rect 52825 7868 52837 7871
rect 52512 7840 52837 7868
rect 52512 7828 52518 7840
rect 52825 7837 52837 7840
rect 52871 7837 52883 7871
rect 54110 7868 54116 7880
rect 54071 7840 54116 7868
rect 52825 7831 52883 7837
rect 54110 7828 54116 7840
rect 54168 7828 54174 7880
rect 54202 7828 54208 7880
rect 54260 7868 54266 7880
rect 54938 7868 54944 7880
rect 54260 7840 54305 7868
rect 54899 7840 54944 7868
rect 54260 7828 54266 7840
rect 54938 7828 54944 7840
rect 54996 7828 55002 7880
rect 57716 7868 57744 7908
rect 59538 7896 59544 7948
rect 59596 7936 59602 7948
rect 61562 7936 61568 7948
rect 59596 7908 61568 7936
rect 59596 7896 59602 7908
rect 61562 7896 61568 7908
rect 61620 7896 61626 7948
rect 63420 7936 63448 8044
rect 66714 8032 66720 8044
rect 66772 8032 66778 8084
rect 68922 8072 68928 8084
rect 68883 8044 68928 8072
rect 68922 8032 68928 8044
rect 68980 8032 68986 8084
rect 74813 8075 74871 8081
rect 74813 8041 74825 8075
rect 74859 8072 74871 8075
rect 75270 8072 75276 8084
rect 74859 8044 75276 8072
rect 74859 8041 74871 8044
rect 74813 8035 74871 8041
rect 75270 8032 75276 8044
rect 75328 8032 75334 8084
rect 76558 8032 76564 8084
rect 76616 8072 76622 8084
rect 76745 8075 76803 8081
rect 76745 8072 76757 8075
rect 76616 8044 76757 8072
rect 76616 8032 76622 8044
rect 76745 8041 76757 8044
rect 76791 8041 76803 8075
rect 80606 8072 80612 8084
rect 80567 8044 80612 8072
rect 76745 8035 76803 8041
rect 80606 8032 80612 8044
rect 80664 8032 80670 8084
rect 83918 8032 83924 8084
rect 83976 8072 83982 8084
rect 84473 8075 84531 8081
rect 84473 8072 84485 8075
rect 83976 8044 84485 8072
rect 83976 8032 83982 8044
rect 84473 8041 84485 8044
rect 84519 8041 84531 8075
rect 112070 8072 112076 8084
rect 84473 8035 84531 8041
rect 84856 8044 112076 8072
rect 64966 7964 64972 8016
rect 65024 8004 65030 8016
rect 65886 8004 65892 8016
rect 65024 7976 65892 8004
rect 65024 7964 65030 7976
rect 65886 7964 65892 7976
rect 65944 7964 65950 8016
rect 73614 7964 73620 8016
rect 73672 8004 73678 8016
rect 84856 8004 84884 8044
rect 112070 8032 112076 8044
rect 112128 8032 112134 8084
rect 112162 8032 112168 8084
rect 112220 8072 112226 8084
rect 112220 8044 119568 8072
rect 112220 8032 112226 8044
rect 73672 7976 84884 8004
rect 86957 8007 87015 8013
rect 73672 7964 73678 7976
rect 86957 7973 86969 8007
rect 87003 8004 87015 8007
rect 87003 7976 89714 8004
rect 87003 7973 87015 7976
rect 86957 7967 87015 7973
rect 66993 7939 67051 7945
rect 66993 7936 67005 7939
rect 62500 7908 63448 7936
rect 65260 7908 67005 7936
rect 58805 7871 58863 7877
rect 57716 7840 58756 7868
rect 44370 7763 44428 7769
rect 44468 7772 47532 7800
rect 44468 7732 44496 7772
rect 49510 7760 49516 7812
rect 49568 7800 49574 7812
rect 49568 7772 49924 7800
rect 49568 7760 49574 7772
rect 41386 7704 44496 7732
rect 46201 7735 46259 7741
rect 34020 7692 34026 7704
rect 46201 7701 46213 7735
rect 46247 7732 46259 7735
rect 46658 7732 46664 7744
rect 46247 7704 46664 7732
rect 46247 7701 46259 7704
rect 46201 7695 46259 7701
rect 46658 7692 46664 7704
rect 46716 7692 46722 7744
rect 47581 7735 47639 7741
rect 47581 7701 47593 7735
rect 47627 7732 47639 7735
rect 47946 7732 47952 7744
rect 47627 7704 47952 7732
rect 47627 7701 47639 7704
rect 47581 7695 47639 7701
rect 47946 7692 47952 7704
rect 48004 7692 48010 7744
rect 49786 7732 49792 7744
rect 49747 7704 49792 7732
rect 49786 7692 49792 7704
rect 49844 7692 49850 7744
rect 49896 7732 49924 7772
rect 50614 7760 50620 7812
rect 50672 7800 50678 7812
rect 52098 7803 52156 7809
rect 52098 7800 52110 7803
rect 50672 7772 52110 7800
rect 50672 7760 50678 7772
rect 52098 7769 52110 7772
rect 52144 7769 52156 7803
rect 52098 7763 52156 7769
rect 52270 7760 52276 7812
rect 52328 7800 52334 7812
rect 56321 7803 56379 7809
rect 56321 7800 56333 7803
rect 52328 7772 56333 7800
rect 52328 7760 52334 7772
rect 56321 7769 56333 7772
rect 56367 7800 56379 7803
rect 58538 7803 58596 7809
rect 58538 7800 58550 7803
rect 56367 7772 58550 7800
rect 56367 7769 56379 7772
rect 56321 7763 56379 7769
rect 58538 7769 58550 7772
rect 58584 7769 58596 7803
rect 58728 7800 58756 7840
rect 58805 7837 58817 7871
rect 58851 7868 58863 7871
rect 59078 7868 59084 7880
rect 58851 7840 59084 7868
rect 58851 7837 58863 7840
rect 58805 7831 58863 7837
rect 59078 7828 59084 7840
rect 59136 7828 59142 7880
rect 62321 7871 62379 7877
rect 62321 7837 62333 7871
rect 62367 7868 62379 7871
rect 62500 7868 62528 7908
rect 65260 7880 65288 7908
rect 66993 7905 67005 7908
rect 67039 7936 67051 7939
rect 67545 7939 67603 7945
rect 67545 7936 67557 7939
rect 67039 7908 67557 7936
rect 67039 7905 67051 7908
rect 66993 7899 67051 7905
rect 67545 7905 67557 7908
rect 67591 7905 67603 7939
rect 67545 7899 67603 7905
rect 62367 7840 62528 7868
rect 62577 7871 62635 7877
rect 62367 7837 62379 7840
rect 62321 7831 62379 7837
rect 62577 7837 62589 7871
rect 62623 7868 62635 7871
rect 62666 7868 62672 7880
rect 62623 7840 62672 7868
rect 62623 7837 62635 7840
rect 62577 7831 62635 7837
rect 62666 7828 62672 7840
rect 62724 7868 62730 7880
rect 64693 7871 64751 7877
rect 64693 7868 64705 7871
rect 62724 7840 64705 7868
rect 62724 7828 62730 7840
rect 64693 7837 64705 7840
rect 64739 7868 64751 7871
rect 65242 7868 65248 7880
rect 64739 7840 65248 7868
rect 64739 7837 64751 7840
rect 64693 7831 64751 7837
rect 65242 7828 65248 7840
rect 65300 7828 65306 7880
rect 66073 7871 66131 7877
rect 66073 7868 66085 7871
rect 65812 7840 66085 7868
rect 59262 7800 59268 7812
rect 58728 7772 59268 7800
rect 58538 7763 58596 7769
rect 59262 7760 59268 7772
rect 59320 7760 59326 7812
rect 60918 7760 60924 7812
rect 60976 7800 60982 7812
rect 64426 7803 64484 7809
rect 64426 7800 64438 7803
rect 60976 7772 64438 7800
rect 60976 7760 60982 7772
rect 64426 7769 64438 7772
rect 64472 7769 64484 7803
rect 64426 7763 64484 7769
rect 51902 7732 51908 7744
rect 49896 7704 51908 7732
rect 51902 7692 51908 7704
rect 51960 7692 51966 7744
rect 53742 7692 53748 7744
rect 53800 7732 53806 7744
rect 53929 7735 53987 7741
rect 53929 7732 53941 7735
rect 53800 7704 53941 7732
rect 53800 7692 53806 7704
rect 53929 7701 53941 7704
rect 53975 7701 53987 7735
rect 54754 7732 54760 7744
rect 54715 7704 54760 7732
rect 53929 7695 53987 7701
rect 54754 7692 54760 7704
rect 54812 7692 54818 7744
rect 60737 7735 60795 7741
rect 60737 7701 60749 7735
rect 60783 7732 60795 7735
rect 60826 7732 60832 7744
rect 60783 7704 60832 7732
rect 60783 7701 60795 7704
rect 60737 7695 60795 7701
rect 60826 7692 60832 7704
rect 60884 7692 60890 7744
rect 65245 7735 65303 7741
rect 65245 7701 65257 7735
rect 65291 7732 65303 7735
rect 65812 7732 65840 7840
rect 66073 7837 66085 7840
rect 66119 7868 66131 7871
rect 66898 7868 66904 7880
rect 66119 7840 66904 7868
rect 66119 7837 66131 7840
rect 66073 7831 66131 7837
rect 66898 7828 66904 7840
rect 66956 7828 66962 7880
rect 67560 7868 67588 7899
rect 80422 7896 80428 7948
rect 80480 7936 80486 7948
rect 85853 7939 85911 7945
rect 80480 7908 84884 7936
rect 80480 7896 80486 7908
rect 72053 7871 72111 7877
rect 72053 7868 72065 7871
rect 67560 7840 72065 7868
rect 72053 7837 72065 7840
rect 72099 7868 72111 7871
rect 72605 7871 72663 7877
rect 72605 7868 72617 7871
rect 72099 7840 72617 7868
rect 72099 7837 72111 7840
rect 72053 7831 72111 7837
rect 72605 7837 72617 7840
rect 72651 7837 72663 7871
rect 72605 7831 72663 7837
rect 72872 7871 72930 7877
rect 72872 7837 72884 7871
rect 72918 7868 72930 7871
rect 73246 7868 73252 7880
rect 72918 7840 73252 7868
rect 72918 7837 72930 7840
rect 72872 7831 72930 7837
rect 73246 7828 73252 7840
rect 73304 7828 73310 7880
rect 74350 7828 74356 7880
rect 74408 7868 74414 7880
rect 74445 7871 74503 7877
rect 74445 7868 74457 7871
rect 74408 7840 74457 7868
rect 74408 7828 74414 7840
rect 74445 7837 74457 7840
rect 74491 7837 74503 7871
rect 74445 7831 74503 7837
rect 74626 7828 74632 7880
rect 74684 7868 74690 7880
rect 75546 7868 75552 7880
rect 74684 7840 75552 7868
rect 74684 7828 74690 7840
rect 75546 7828 75552 7840
rect 75604 7828 75610 7880
rect 76282 7868 76288 7880
rect 76243 7840 76288 7868
rect 76282 7828 76288 7840
rect 76340 7828 76346 7880
rect 80606 7828 80612 7880
rect 80664 7868 80670 7880
rect 81253 7871 81311 7877
rect 81253 7868 81265 7871
rect 80664 7840 81265 7868
rect 80664 7828 80670 7840
rect 81253 7837 81265 7840
rect 81299 7837 81311 7871
rect 84856 7868 84884 7908
rect 85853 7905 85865 7939
rect 85899 7936 85911 7939
rect 86402 7936 86408 7948
rect 85899 7908 86408 7936
rect 85899 7905 85911 7908
rect 85853 7899 85911 7905
rect 86402 7896 86408 7908
rect 86460 7896 86466 7948
rect 87874 7936 87880 7948
rect 87616 7908 87880 7936
rect 87616 7877 87644 7908
rect 87874 7896 87880 7908
rect 87932 7896 87938 7948
rect 89686 7936 89714 7976
rect 90082 7964 90088 8016
rect 90140 8004 90146 8016
rect 90453 8007 90511 8013
rect 90453 8004 90465 8007
rect 90140 7976 90465 8004
rect 90140 7964 90146 7976
rect 90453 7973 90465 7976
rect 90499 8004 90511 8007
rect 90634 8004 90640 8016
rect 90499 7976 90640 8004
rect 90499 7973 90511 7976
rect 90453 7967 90511 7973
rect 90634 7964 90640 7976
rect 90692 7964 90698 8016
rect 90726 7964 90732 8016
rect 90784 8004 90790 8016
rect 91557 8007 91615 8013
rect 91557 8004 91569 8007
rect 90784 7976 91569 8004
rect 90784 7964 90790 7976
rect 91557 7973 91569 7976
rect 91603 7973 91615 8007
rect 91557 7967 91615 7973
rect 92934 7964 92940 8016
rect 92992 8004 92998 8016
rect 93489 8007 93547 8013
rect 93489 8004 93501 8007
rect 92992 7976 93501 8004
rect 92992 7964 92998 7976
rect 93489 7973 93501 7976
rect 93535 8004 93547 8007
rect 98270 8004 98276 8016
rect 93535 7976 98276 8004
rect 93535 7973 93547 7976
rect 93489 7967 93547 7973
rect 98270 7964 98276 7976
rect 98328 7964 98334 8016
rect 99745 8007 99803 8013
rect 99745 7973 99757 8007
rect 99791 8004 99803 8007
rect 100110 8004 100116 8016
rect 99791 7976 100116 8004
rect 99791 7973 99803 7976
rect 99745 7967 99803 7973
rect 100110 7964 100116 7976
rect 100168 7964 100174 8016
rect 110414 7964 110420 8016
rect 110472 8004 110478 8016
rect 110509 8007 110567 8013
rect 110509 8004 110521 8007
rect 110472 7976 110521 8004
rect 110472 7964 110478 7976
rect 110509 7973 110521 7976
rect 110555 7973 110567 8007
rect 110509 7967 110567 7973
rect 112530 7964 112536 8016
rect 112588 8004 112594 8016
rect 112625 8007 112683 8013
rect 112625 8004 112637 8007
rect 112588 7976 112637 8004
rect 112588 7964 112594 7976
rect 112625 7973 112637 7976
rect 112671 7973 112683 8007
rect 112625 7967 112683 7973
rect 117130 7964 117136 8016
rect 117188 8004 117194 8016
rect 119430 8004 119436 8016
rect 117188 7976 119436 8004
rect 117188 7964 117194 7976
rect 119430 7964 119436 7976
rect 119488 7964 119494 8016
rect 91370 7936 91376 7948
rect 89686 7908 91376 7936
rect 91370 7896 91376 7908
rect 91428 7896 91434 7948
rect 93762 7896 93768 7948
rect 93820 7936 93826 7948
rect 93820 7908 98500 7936
rect 93820 7896 93826 7908
rect 86773 7871 86831 7877
rect 84856 7840 85712 7868
rect 81253 7831 81311 7837
rect 67082 7760 67088 7812
rect 67140 7800 67146 7812
rect 67790 7803 67848 7809
rect 67790 7800 67802 7803
rect 67140 7772 67802 7800
rect 67140 7760 67146 7772
rect 67790 7769 67802 7772
rect 67836 7769 67848 7803
rect 67790 7763 67848 7769
rect 81434 7760 81440 7812
rect 81492 7800 81498 7812
rect 85574 7800 85580 7812
rect 85632 7809 85638 7812
rect 81492 7772 82676 7800
rect 85544 7772 85580 7800
rect 81492 7760 81498 7772
rect 65291 7704 65840 7732
rect 73985 7735 74043 7741
rect 65291 7701 65303 7704
rect 65245 7695 65303 7701
rect 73985 7701 73997 7735
rect 74031 7732 74043 7735
rect 75546 7732 75552 7744
rect 74031 7704 75552 7732
rect 74031 7701 74043 7704
rect 73985 7695 74043 7701
rect 75546 7692 75552 7704
rect 75604 7692 75610 7744
rect 76006 7692 76012 7744
rect 76064 7732 76070 7744
rect 76101 7735 76159 7741
rect 76101 7732 76113 7735
rect 76064 7704 76113 7732
rect 76064 7692 76070 7704
rect 76101 7701 76113 7704
rect 76147 7701 76159 7735
rect 76101 7695 76159 7701
rect 81250 7692 81256 7744
rect 81308 7732 81314 7744
rect 82541 7735 82599 7741
rect 82541 7732 82553 7735
rect 81308 7704 82553 7732
rect 81308 7692 81314 7704
rect 82541 7701 82553 7704
rect 82587 7701 82599 7735
rect 82648 7732 82676 7772
rect 85574 7760 85580 7772
rect 85632 7763 85644 7809
rect 85684 7800 85712 7840
rect 86773 7837 86785 7871
rect 86819 7868 86831 7871
rect 87417 7871 87475 7877
rect 87417 7868 87429 7871
rect 86819 7840 87429 7868
rect 86819 7837 86831 7840
rect 86773 7831 86831 7837
rect 87417 7837 87429 7840
rect 87463 7837 87475 7871
rect 87417 7831 87475 7837
rect 87601 7871 87659 7877
rect 87601 7837 87613 7871
rect 87647 7837 87659 7871
rect 87601 7831 87659 7837
rect 87690 7828 87696 7880
rect 87748 7868 87754 7880
rect 87748 7840 87793 7868
rect 87748 7828 87754 7840
rect 89622 7828 89628 7880
rect 89680 7868 89686 7880
rect 90818 7868 90824 7880
rect 89680 7840 90824 7868
rect 89680 7828 89686 7840
rect 90818 7828 90824 7840
rect 90876 7828 90882 7880
rect 91002 7828 91008 7880
rect 91060 7868 91066 7880
rect 92382 7868 92388 7880
rect 91060 7840 92388 7868
rect 91060 7828 91066 7840
rect 92382 7828 92388 7840
rect 92440 7828 92446 7880
rect 92937 7871 92995 7877
rect 92937 7837 92949 7871
rect 92983 7868 92995 7871
rect 93026 7868 93032 7880
rect 92983 7840 93032 7868
rect 92983 7837 92995 7840
rect 92937 7831 92995 7837
rect 93026 7828 93032 7840
rect 93084 7828 93090 7880
rect 95326 7868 95332 7880
rect 95287 7840 95332 7868
rect 95326 7828 95332 7840
rect 95384 7828 95390 7880
rect 98086 7828 98092 7880
rect 98144 7868 98150 7880
rect 98365 7871 98423 7877
rect 98365 7868 98377 7871
rect 98144 7840 98377 7868
rect 98144 7828 98150 7840
rect 98365 7837 98377 7840
rect 98411 7837 98423 7871
rect 98472 7868 98500 7908
rect 101416 7908 109264 7936
rect 101416 7868 101444 7908
rect 98472 7840 101444 7868
rect 98365 7831 98423 7837
rect 105354 7828 105360 7880
rect 105412 7868 105418 7880
rect 105725 7871 105783 7877
rect 105725 7868 105737 7871
rect 105412 7840 105737 7868
rect 105412 7828 105418 7840
rect 105725 7837 105737 7840
rect 105771 7837 105783 7871
rect 109126 7868 109132 7880
rect 109087 7840 109132 7868
rect 105725 7831 105783 7837
rect 109126 7828 109132 7840
rect 109184 7828 109190 7880
rect 109236 7868 109264 7908
rect 110340 7908 112760 7936
rect 110340 7868 110368 7908
rect 112732 7880 112760 7908
rect 117590 7896 117596 7948
rect 117648 7936 117654 7948
rect 118602 7936 118608 7948
rect 117648 7908 118608 7936
rect 117648 7896 117654 7908
rect 118602 7896 118608 7908
rect 118660 7896 118666 7948
rect 119540 7936 119568 8044
rect 121270 8032 121276 8084
rect 121328 8072 121334 8084
rect 124030 8072 124036 8084
rect 121328 8044 124036 8072
rect 121328 8032 121334 8044
rect 124030 8032 124036 8044
rect 124088 8032 124094 8084
rect 124950 8032 124956 8084
rect 125008 8072 125014 8084
rect 125321 8075 125379 8081
rect 125321 8072 125333 8075
rect 125008 8044 125333 8072
rect 125008 8032 125014 8044
rect 125321 8041 125333 8044
rect 125367 8041 125379 8075
rect 125321 8035 125379 8041
rect 127158 8032 127164 8084
rect 127216 8072 127222 8084
rect 127621 8075 127679 8081
rect 127621 8072 127633 8075
rect 127216 8044 127633 8072
rect 127216 8032 127222 8044
rect 127621 8041 127633 8044
rect 127667 8041 127679 8075
rect 127621 8035 127679 8041
rect 127728 8044 129044 8072
rect 121822 7964 121828 8016
rect 121880 8004 121886 8016
rect 122469 8007 122527 8013
rect 122469 8004 122481 8007
rect 121880 7976 122481 8004
rect 121880 7964 121886 7976
rect 122469 7973 122481 7976
rect 122515 7973 122527 8007
rect 122469 7967 122527 7973
rect 123018 7964 123024 8016
rect 123076 8004 123082 8016
rect 123294 8004 123300 8016
rect 123076 7976 123300 8004
rect 123076 7964 123082 7976
rect 123294 7964 123300 7976
rect 123352 8004 123358 8016
rect 127728 8004 127756 8044
rect 123352 7976 127756 8004
rect 123352 7964 123358 7976
rect 121641 7939 121699 7945
rect 121641 7936 121653 7939
rect 119540 7908 121653 7936
rect 109236 7840 110368 7868
rect 110966 7828 110972 7880
rect 111024 7828 111030 7880
rect 111058 7828 111064 7880
rect 111116 7868 111122 7880
rect 111153 7871 111211 7877
rect 111153 7868 111165 7871
rect 111116 7840 111165 7868
rect 111116 7828 111122 7840
rect 111153 7837 111165 7840
rect 111199 7837 111211 7871
rect 111153 7831 111211 7837
rect 112714 7828 112720 7880
rect 112772 7868 112778 7880
rect 112809 7871 112867 7877
rect 112809 7868 112821 7871
rect 112772 7840 112821 7868
rect 112772 7828 112778 7840
rect 112809 7837 112821 7840
rect 112855 7837 112867 7871
rect 112809 7831 112867 7837
rect 112898 7828 112904 7880
rect 112956 7868 112962 7880
rect 112956 7840 113001 7868
rect 112956 7828 112962 7840
rect 113082 7828 113088 7880
rect 113140 7868 113146 7880
rect 113729 7871 113787 7877
rect 113729 7868 113741 7871
rect 113140 7840 113741 7868
rect 113140 7828 113146 7840
rect 113729 7837 113741 7840
rect 113775 7868 113787 7871
rect 115569 7871 115627 7877
rect 115569 7868 115581 7871
rect 113775 7840 115581 7868
rect 113775 7837 113787 7840
rect 113729 7831 113787 7837
rect 115569 7837 115581 7840
rect 115615 7868 115627 7871
rect 117130 7868 117136 7880
rect 115615 7840 117136 7868
rect 115615 7837 115627 7840
rect 115569 7831 115627 7837
rect 117130 7828 117136 7840
rect 117188 7828 117194 7880
rect 117406 7828 117412 7880
rect 117464 7868 117470 7880
rect 117869 7871 117927 7877
rect 117869 7868 117881 7871
rect 117464 7840 117881 7868
rect 117464 7828 117470 7840
rect 117869 7837 117881 7840
rect 117915 7837 117927 7871
rect 117869 7831 117927 7837
rect 118694 7828 118700 7880
rect 118752 7868 118758 7880
rect 118789 7871 118847 7877
rect 118789 7868 118801 7871
rect 118752 7840 118801 7868
rect 118752 7828 118758 7840
rect 118789 7837 118801 7840
rect 118835 7837 118847 7871
rect 118789 7831 118847 7837
rect 119433 7871 119491 7877
rect 119433 7837 119445 7871
rect 119479 7868 119491 7871
rect 119540 7868 119568 7908
rect 121641 7905 121653 7908
rect 121687 7905 121699 7939
rect 121641 7899 121699 7905
rect 123404 7908 124352 7936
rect 119479 7840 119568 7868
rect 121656 7868 121684 7899
rect 123404 7868 123432 7908
rect 123941 7871 123999 7877
rect 123941 7868 123953 7871
rect 121656 7840 123432 7868
rect 123496 7840 123953 7868
rect 119479 7837 119491 7840
rect 119433 7831 119491 7837
rect 90726 7800 90732 7812
rect 85684 7772 90732 7800
rect 85632 7760 85638 7763
rect 90726 7760 90732 7772
rect 90784 7760 90790 7812
rect 92658 7760 92664 7812
rect 92716 7809 92722 7812
rect 92716 7800 92728 7809
rect 98454 7800 98460 7812
rect 92716 7772 92761 7800
rect 92952 7772 98460 7800
rect 92716 7763 92728 7772
rect 92716 7760 92722 7763
rect 92952 7744 92980 7772
rect 98454 7760 98460 7772
rect 98512 7760 98518 7812
rect 98632 7803 98690 7809
rect 98632 7769 98644 7803
rect 98678 7800 98690 7803
rect 98678 7772 98960 7800
rect 98678 7769 98690 7772
rect 98632 7763 98690 7769
rect 90818 7732 90824 7744
rect 82648 7704 90824 7732
rect 82541 7695 82599 7701
rect 90818 7692 90824 7704
rect 90876 7692 90882 7744
rect 91370 7692 91376 7744
rect 91428 7732 91434 7744
rect 92474 7732 92480 7744
rect 91428 7704 92480 7732
rect 91428 7692 91434 7704
rect 92474 7692 92480 7704
rect 92532 7692 92538 7744
rect 92934 7692 92940 7744
rect 92992 7692 92998 7744
rect 94038 7732 94044 7744
rect 93999 7704 94044 7732
rect 94038 7692 94044 7704
rect 94096 7732 94102 7744
rect 95050 7732 95056 7744
rect 94096 7704 95056 7732
rect 94096 7692 94102 7704
rect 95050 7692 95056 7704
rect 95108 7692 95114 7744
rect 95142 7692 95148 7744
rect 95200 7732 95206 7744
rect 97810 7732 97816 7744
rect 95200 7704 95245 7732
rect 97771 7704 97816 7732
rect 95200 7692 95206 7704
rect 97810 7692 97816 7704
rect 97868 7692 97874 7744
rect 98932 7732 98960 7772
rect 99190 7760 99196 7812
rect 99248 7800 99254 7812
rect 104894 7800 104900 7812
rect 99248 7772 104900 7800
rect 99248 7760 99254 7772
rect 104894 7760 104900 7772
rect 104952 7760 104958 7812
rect 106734 7760 106740 7812
rect 106792 7800 106798 7812
rect 107286 7800 107292 7812
rect 106792 7772 107292 7800
rect 106792 7760 106798 7772
rect 107286 7760 107292 7772
rect 107344 7800 107350 7812
rect 109396 7803 109454 7809
rect 107344 7772 109264 7800
rect 107344 7760 107350 7772
rect 100294 7732 100300 7744
rect 98932 7704 100300 7732
rect 100294 7692 100300 7704
rect 100352 7692 100358 7744
rect 105909 7735 105967 7741
rect 105909 7701 105921 7735
rect 105955 7732 105967 7735
rect 107194 7732 107200 7744
rect 105955 7704 107200 7732
rect 105955 7701 105967 7704
rect 105909 7695 105967 7701
rect 107194 7692 107200 7704
rect 107252 7692 107258 7744
rect 109236 7732 109264 7772
rect 109396 7769 109408 7803
rect 109442 7800 109454 7803
rect 109770 7800 109776 7812
rect 109442 7772 109776 7800
rect 109442 7769 109454 7772
rect 109396 7763 109454 7769
rect 109770 7760 109776 7772
rect 109828 7760 109834 7812
rect 109862 7760 109868 7812
rect 109920 7800 109926 7812
rect 110984 7800 111012 7828
rect 112990 7800 112996 7812
rect 109920 7772 110920 7800
rect 110984 7772 112996 7800
rect 109920 7760 109926 7772
rect 110690 7732 110696 7744
rect 109236 7704 110696 7732
rect 110690 7692 110696 7704
rect 110748 7692 110754 7744
rect 110892 7732 110920 7772
rect 112990 7760 112996 7772
rect 113048 7760 113054 7812
rect 113996 7803 114054 7809
rect 113996 7769 114008 7803
rect 114042 7800 114054 7803
rect 115474 7800 115480 7812
rect 114042 7772 115480 7800
rect 114042 7769 114054 7772
rect 113996 7763 114054 7769
rect 115474 7760 115480 7772
rect 115532 7760 115538 7812
rect 116210 7800 116216 7812
rect 116171 7772 116216 7800
rect 116210 7760 116216 7772
rect 116268 7760 116274 7812
rect 116302 7760 116308 7812
rect 116360 7800 116366 7812
rect 121181 7803 121239 7809
rect 116360 7772 117728 7800
rect 116360 7760 116366 7772
rect 110969 7735 111027 7741
rect 110969 7732 110981 7735
rect 110892 7704 110981 7732
rect 110969 7701 110981 7704
rect 111015 7701 111027 7735
rect 110969 7695 111027 7701
rect 114830 7692 114836 7744
rect 114888 7732 114894 7744
rect 115109 7735 115167 7741
rect 115109 7732 115121 7735
rect 114888 7704 115121 7732
rect 114888 7692 114894 7704
rect 115109 7701 115121 7704
rect 115155 7701 115167 7735
rect 115109 7695 115167 7701
rect 116765 7735 116823 7741
rect 116765 7701 116777 7735
rect 116811 7732 116823 7735
rect 117038 7732 117044 7744
rect 116811 7704 117044 7732
rect 116811 7701 116823 7704
rect 116765 7695 116823 7701
rect 117038 7692 117044 7704
rect 117096 7692 117102 7744
rect 117700 7741 117728 7772
rect 121181 7769 121193 7803
rect 121227 7800 121239 7803
rect 121454 7800 121460 7812
rect 121227 7772 121460 7800
rect 121227 7769 121239 7772
rect 121181 7763 121239 7769
rect 121454 7760 121460 7772
rect 121512 7800 121518 7812
rect 121638 7800 121644 7812
rect 121512 7772 121644 7800
rect 121512 7760 121518 7772
rect 121638 7760 121644 7772
rect 121696 7760 121702 7812
rect 122466 7760 122472 7812
rect 122524 7800 122530 7812
rect 122653 7803 122711 7809
rect 122653 7800 122665 7803
rect 122524 7772 122665 7800
rect 122524 7760 122530 7772
rect 122653 7769 122665 7772
rect 122699 7769 122711 7803
rect 123496 7800 123524 7840
rect 123941 7837 123953 7840
rect 123987 7837 123999 7871
rect 124214 7868 124220 7880
rect 124175 7840 124220 7868
rect 123941 7831 123999 7837
rect 124214 7828 124220 7840
rect 124272 7828 124278 7880
rect 124324 7868 124352 7908
rect 124398 7896 124404 7948
rect 124456 7936 124462 7948
rect 127066 7936 127072 7948
rect 124456 7908 127072 7936
rect 124456 7896 124462 7908
rect 127066 7896 127072 7908
rect 127124 7896 127130 7948
rect 129016 7945 129044 8044
rect 130286 8032 130292 8084
rect 130344 8072 130350 8084
rect 130344 8044 135852 8072
rect 130344 8032 130350 8044
rect 129642 7964 129648 8016
rect 129700 8004 129706 8016
rect 129700 7976 130056 8004
rect 129700 7964 129706 7976
rect 129001 7939 129059 7945
rect 129001 7905 129013 7939
rect 129047 7905 129059 7939
rect 129001 7899 129059 7905
rect 129752 7877 129780 7976
rect 130028 7936 130056 7976
rect 130378 7964 130384 8016
rect 130436 8004 130442 8016
rect 132129 8007 132187 8013
rect 132129 8004 132141 8007
rect 130436 7976 132141 8004
rect 130436 7964 130442 7976
rect 132129 7973 132141 7976
rect 132175 8004 132187 8007
rect 134334 8004 134340 8016
rect 132175 7976 134340 8004
rect 132175 7973 132187 7976
rect 132129 7967 132187 7973
rect 134334 7964 134340 7976
rect 134392 7964 134398 8016
rect 132773 7939 132831 7945
rect 130028 7908 131528 7936
rect 129737 7871 129795 7877
rect 124324 7840 129688 7868
rect 122653 7763 122711 7769
rect 122760 7772 123524 7800
rect 117685 7735 117743 7741
rect 117685 7701 117697 7735
rect 117731 7701 117743 7735
rect 117685 7695 117743 7701
rect 118973 7735 119031 7741
rect 118973 7701 118985 7735
rect 119019 7732 119031 7735
rect 122760 7732 122788 7772
rect 124030 7760 124036 7812
rect 124088 7800 124094 7812
rect 128734 7803 128792 7809
rect 124088 7772 127756 7800
rect 124088 7760 124094 7772
rect 119019 7704 122788 7732
rect 119019 7701 119031 7704
rect 118973 7695 119031 7701
rect 122834 7692 122840 7744
rect 122892 7732 122898 7744
rect 123202 7732 123208 7744
rect 122892 7704 123208 7732
rect 122892 7692 122898 7704
rect 123202 7692 123208 7704
rect 123260 7692 123266 7744
rect 125870 7732 125876 7744
rect 125831 7704 125876 7732
rect 125870 7692 125876 7704
rect 125928 7692 125934 7744
rect 126238 7692 126244 7744
rect 126296 7732 126302 7744
rect 126425 7735 126483 7741
rect 126425 7732 126437 7735
rect 126296 7704 126437 7732
rect 126296 7692 126302 7704
rect 126425 7701 126437 7704
rect 126471 7701 126483 7735
rect 127066 7732 127072 7744
rect 127027 7704 127072 7732
rect 126425 7695 126483 7701
rect 127066 7692 127072 7704
rect 127124 7692 127130 7744
rect 127728 7732 127756 7772
rect 128734 7769 128746 7803
rect 128780 7800 128792 7803
rect 129274 7800 129280 7812
rect 128780 7772 129280 7800
rect 128780 7769 128792 7772
rect 128734 7763 128792 7769
rect 129274 7760 129280 7772
rect 129332 7760 129338 7812
rect 129660 7800 129688 7840
rect 129737 7837 129749 7871
rect 129783 7837 129795 7871
rect 129737 7831 129795 7837
rect 129918 7828 129924 7880
rect 129976 7868 129982 7880
rect 130102 7868 130108 7880
rect 129976 7840 130021 7868
rect 130063 7840 130108 7868
rect 129976 7828 129982 7840
rect 130102 7828 130108 7840
rect 130160 7828 130166 7880
rect 130654 7868 130660 7880
rect 130615 7840 130660 7868
rect 130654 7828 130660 7840
rect 130712 7828 130718 7880
rect 131500 7877 131528 7908
rect 132773 7905 132785 7939
rect 132819 7936 132831 7939
rect 132862 7936 132868 7948
rect 132819 7908 132868 7936
rect 132819 7905 132831 7908
rect 132773 7899 132831 7905
rect 132862 7896 132868 7908
rect 132920 7896 132926 7948
rect 132954 7896 132960 7948
rect 133012 7936 133018 7948
rect 133049 7939 133107 7945
rect 133049 7936 133061 7939
rect 133012 7908 133061 7936
rect 133012 7896 133018 7908
rect 133049 7905 133061 7908
rect 133095 7905 133107 7939
rect 133049 7899 133107 7905
rect 133138 7896 133144 7948
rect 133196 7936 133202 7948
rect 133598 7936 133604 7948
rect 133196 7908 133604 7936
rect 133196 7896 133202 7908
rect 133598 7896 133604 7908
rect 133656 7936 133662 7948
rect 134794 7936 134800 7948
rect 133656 7908 134800 7936
rect 133656 7896 133662 7908
rect 134794 7896 134800 7908
rect 134852 7896 134858 7948
rect 135824 7936 135852 8044
rect 136450 8032 136456 8084
rect 136508 8072 136514 8084
rect 137373 8075 137431 8081
rect 137373 8072 137385 8075
rect 136508 8044 137385 8072
rect 136508 8032 136514 8044
rect 137373 8041 137385 8044
rect 137419 8072 137431 8075
rect 137830 8072 137836 8084
rect 137419 8044 137836 8072
rect 137419 8041 137431 8044
rect 137373 8035 137431 8041
rect 137830 8032 137836 8044
rect 137888 8072 137894 8084
rect 138198 8072 138204 8084
rect 137888 8044 138204 8072
rect 137888 8032 137894 8044
rect 138198 8032 138204 8044
rect 138256 8032 138262 8084
rect 138566 8032 138572 8084
rect 138624 8072 138630 8084
rect 142982 8072 142988 8084
rect 138624 8044 142988 8072
rect 138624 8032 138630 8044
rect 138658 7936 138664 7948
rect 135824 7908 138664 7936
rect 138658 7896 138664 7908
rect 138716 7896 138722 7948
rect 140148 7945 140176 8044
rect 142982 8032 142988 8044
rect 143040 8032 143046 8084
rect 143092 8044 144592 8072
rect 140222 7964 140228 8016
rect 140280 8004 140286 8016
rect 141418 8004 141424 8016
rect 140280 7976 141188 8004
rect 141379 7976 141424 8004
rect 140280 7964 140286 7976
rect 140133 7939 140191 7945
rect 140133 7905 140145 7939
rect 140179 7905 140191 7939
rect 141050 7936 141056 7948
rect 140133 7899 140191 7905
rect 140608 7908 141056 7936
rect 130749 7871 130807 7877
rect 130749 7837 130761 7871
rect 130795 7837 130807 7871
rect 130749 7831 130807 7837
rect 131485 7871 131543 7877
rect 131485 7837 131497 7871
rect 131531 7868 131543 7871
rect 133506 7868 133512 7880
rect 131531 7840 133512 7868
rect 131531 7837 131543 7840
rect 131485 7831 131543 7837
rect 130562 7800 130568 7812
rect 129660 7772 130568 7800
rect 130562 7760 130568 7772
rect 130620 7760 130626 7812
rect 130764 7732 130792 7831
rect 133506 7828 133512 7840
rect 133564 7828 133570 7880
rect 133782 7828 133788 7880
rect 133840 7868 133846 7880
rect 135714 7868 135720 7880
rect 133840 7840 135720 7868
rect 133840 7828 133846 7840
rect 135714 7828 135720 7840
rect 135772 7868 135778 7880
rect 135809 7871 135867 7877
rect 135809 7868 135821 7871
rect 135772 7840 135821 7868
rect 135772 7828 135778 7840
rect 135809 7837 135821 7840
rect 135855 7837 135867 7871
rect 135809 7831 135867 7837
rect 138109 7871 138167 7877
rect 138109 7837 138121 7871
rect 138155 7868 138167 7871
rect 140608 7868 140636 7908
rect 141050 7896 141056 7908
rect 141108 7896 141114 7948
rect 138155 7840 140636 7868
rect 138155 7837 138167 7840
rect 138109 7831 138167 7837
rect 140682 7828 140688 7880
rect 140740 7868 140746 7880
rect 140777 7871 140835 7877
rect 140777 7868 140789 7871
rect 140740 7840 140789 7868
rect 140740 7828 140746 7840
rect 140777 7837 140789 7840
rect 140823 7837 140835 7871
rect 140777 7831 140835 7837
rect 140961 7871 141019 7877
rect 140961 7837 140973 7871
rect 141007 7868 141019 7871
rect 141160 7868 141188 7976
rect 141418 7964 141424 7976
rect 141476 7964 141482 8016
rect 141326 7896 141332 7948
rect 141384 7936 141390 7948
rect 143092 7936 143120 8044
rect 144457 8007 144515 8013
rect 144457 7973 144469 8007
rect 144503 7973 144515 8007
rect 144564 8004 144592 8044
rect 144730 8032 144736 8084
rect 144788 8072 144794 8084
rect 149882 8072 149888 8084
rect 144788 8044 147674 8072
rect 144788 8032 144794 8044
rect 144917 8007 144975 8013
rect 144917 8004 144929 8007
rect 144564 7976 144929 8004
rect 144457 7967 144515 7973
rect 144917 7973 144929 7976
rect 144963 8004 144975 8007
rect 145190 8004 145196 8016
rect 144963 7976 145196 8004
rect 144963 7973 144975 7976
rect 144917 7967 144975 7973
rect 141384 7908 143120 7936
rect 141384 7896 141390 7908
rect 141007 7840 141188 7868
rect 141605 7871 141663 7877
rect 141007 7837 141019 7840
rect 140961 7831 141019 7837
rect 141605 7837 141617 7871
rect 141651 7868 141663 7871
rect 142982 7868 142988 7880
rect 141651 7840 142988 7868
rect 141651 7837 141663 7840
rect 141605 7831 141663 7837
rect 142982 7828 142988 7840
rect 143040 7828 143046 7880
rect 143074 7828 143080 7880
rect 143132 7868 143138 7880
rect 144362 7868 144368 7880
rect 143132 7840 143177 7868
rect 143276 7840 144368 7868
rect 143132 7828 143138 7840
rect 135346 7800 135352 7812
rect 132880 7772 135352 7800
rect 127728 7704 130792 7732
rect 130933 7735 130991 7741
rect 130933 7701 130945 7735
rect 130979 7732 130991 7735
rect 132880 7732 132908 7772
rect 135346 7760 135352 7772
rect 135404 7760 135410 7812
rect 135564 7803 135622 7809
rect 135564 7769 135576 7803
rect 135610 7800 135622 7803
rect 136358 7800 136364 7812
rect 135610 7772 136364 7800
rect 135610 7769 135622 7772
rect 135564 7763 135622 7769
rect 136358 7760 136364 7772
rect 136416 7760 136422 7812
rect 137738 7760 137744 7812
rect 137796 7800 137802 7812
rect 137796 7772 138612 7800
rect 137796 7760 137802 7772
rect 130979 7704 132908 7732
rect 130979 7701 130991 7704
rect 130933 7695 130991 7701
rect 132954 7692 132960 7744
rect 133012 7732 133018 7744
rect 133690 7732 133696 7744
rect 133012 7704 133696 7732
rect 133012 7692 133018 7704
rect 133690 7692 133696 7704
rect 133748 7692 133754 7744
rect 134426 7732 134432 7744
rect 134387 7704 134432 7732
rect 134426 7692 134432 7704
rect 134484 7692 134490 7744
rect 137370 7692 137376 7744
rect 137428 7732 137434 7744
rect 137925 7735 137983 7741
rect 137925 7732 137937 7735
rect 137428 7704 137937 7732
rect 137428 7692 137434 7704
rect 137925 7701 137937 7704
rect 137971 7701 137983 7735
rect 138584 7732 138612 7772
rect 139854 7760 139860 7812
rect 139912 7809 139918 7812
rect 139912 7800 139924 7809
rect 139912 7772 139957 7800
rect 139912 7763 139924 7772
rect 139912 7760 139918 7763
rect 140406 7760 140412 7812
rect 140464 7800 140470 7812
rect 140464 7772 140728 7800
rect 140464 7760 140470 7772
rect 138753 7735 138811 7741
rect 138753 7732 138765 7735
rect 138584 7704 138765 7732
rect 137925 7695 137983 7701
rect 138753 7701 138765 7704
rect 138799 7701 138811 7735
rect 138753 7695 138811 7701
rect 139762 7692 139768 7744
rect 139820 7732 139826 7744
rect 140593 7735 140651 7741
rect 140593 7732 140605 7735
rect 139820 7704 140605 7732
rect 139820 7692 139826 7704
rect 140593 7701 140605 7704
rect 140639 7701 140651 7735
rect 140700 7732 140728 7772
rect 141050 7760 141056 7812
rect 141108 7800 141114 7812
rect 142157 7803 142215 7809
rect 142157 7800 142169 7803
rect 141108 7772 142169 7800
rect 141108 7760 141114 7772
rect 142157 7769 142169 7772
rect 142203 7800 142215 7803
rect 143276 7800 143304 7840
rect 144362 7828 144368 7840
rect 144420 7828 144426 7880
rect 144472 7868 144500 7967
rect 145190 7964 145196 7976
rect 145248 7964 145254 8016
rect 147214 7964 147220 8016
rect 147272 7964 147278 8016
rect 147646 8004 147674 8044
rect 148244 8044 149888 8072
rect 148134 8004 148140 8016
rect 147646 7976 148140 8004
rect 148134 7964 148140 7976
rect 148192 7964 148198 8016
rect 146754 7896 146760 7948
rect 146812 7936 146818 7948
rect 147030 7936 147036 7948
rect 146812 7908 147036 7936
rect 146812 7896 146818 7908
rect 147030 7896 147036 7908
rect 147088 7896 147094 7948
rect 147125 7939 147183 7945
rect 147125 7905 147137 7939
rect 147171 7936 147183 7939
rect 147232 7936 147260 7964
rect 147171 7908 147260 7936
rect 147493 7939 147551 7945
rect 147171 7905 147183 7908
rect 147125 7899 147183 7905
rect 147493 7905 147505 7939
rect 147539 7936 147551 7939
rect 148244 7936 148272 8044
rect 149882 8032 149888 8044
rect 149940 8032 149946 8084
rect 150158 8032 150164 8084
rect 150216 8072 150222 8084
rect 151814 8072 151820 8084
rect 150216 8044 151820 8072
rect 150216 8032 150222 8044
rect 151814 8032 151820 8044
rect 151872 8032 151878 8084
rect 152093 8075 152151 8081
rect 152093 8041 152105 8075
rect 152139 8072 152151 8075
rect 152274 8072 152280 8084
rect 152139 8044 152280 8072
rect 152139 8041 152151 8044
rect 152093 8035 152151 8041
rect 152274 8032 152280 8044
rect 152332 8032 152338 8084
rect 152366 8032 152372 8084
rect 152424 8072 152430 8084
rect 154758 8072 154764 8084
rect 152424 8044 154764 8072
rect 152424 8032 152430 8044
rect 154758 8032 154764 8044
rect 154816 8032 154822 8084
rect 155862 8032 155868 8084
rect 155920 8072 155926 8084
rect 157245 8075 157303 8081
rect 157245 8072 157257 8075
rect 155920 8044 157257 8072
rect 155920 8032 155926 8044
rect 157245 8041 157257 8044
rect 157291 8041 157303 8075
rect 157245 8035 157303 8041
rect 149238 7964 149244 8016
rect 149296 8004 149302 8016
rect 150345 8007 150403 8013
rect 150345 8004 150357 8007
rect 149296 7976 150357 8004
rect 149296 7964 149302 7976
rect 150345 7973 150357 7976
rect 150391 8004 150403 8007
rect 154298 8004 154304 8016
rect 150391 7976 154304 8004
rect 150391 7973 150403 7976
rect 150345 7967 150403 7973
rect 154298 7964 154304 7976
rect 154356 7964 154362 8016
rect 147539 7908 148272 7936
rect 147539 7905 147551 7908
rect 147493 7899 147551 7905
rect 150894 7896 150900 7948
rect 150952 7936 150958 7948
rect 150952 7908 152596 7936
rect 150952 7896 150958 7908
rect 146297 7871 146355 7877
rect 144472 7840 146248 7868
rect 142203 7772 143304 7800
rect 143344 7803 143402 7809
rect 142203 7769 142215 7772
rect 142157 7763 142215 7769
rect 143344 7769 143356 7803
rect 143390 7800 143402 7803
rect 145742 7800 145748 7812
rect 143390 7772 145748 7800
rect 143390 7769 143402 7772
rect 143344 7763 143402 7769
rect 145742 7760 145748 7772
rect 145800 7760 145806 7812
rect 146030 7803 146088 7809
rect 146030 7769 146042 7803
rect 146076 7769 146088 7803
rect 146220 7800 146248 7840
rect 146297 7837 146309 7871
rect 146343 7868 146355 7871
rect 146386 7868 146392 7880
rect 146343 7840 146392 7868
rect 146343 7837 146355 7840
rect 146297 7831 146355 7837
rect 146386 7828 146392 7840
rect 146444 7828 146450 7880
rect 147306 7868 147312 7880
rect 147267 7840 147312 7868
rect 147306 7828 147312 7840
rect 147364 7828 147370 7880
rect 147950 7868 147956 7880
rect 147416 7840 147956 7868
rect 146220 7772 146892 7800
rect 146030 7763 146088 7769
rect 142246 7732 142252 7744
rect 140700 7704 142252 7732
rect 140593 7695 140651 7701
rect 142246 7692 142252 7704
rect 142304 7692 142310 7744
rect 142430 7732 142436 7744
rect 142391 7704 142436 7732
rect 142430 7692 142436 7704
rect 142488 7692 142494 7744
rect 142982 7692 142988 7744
rect 143040 7732 143046 7744
rect 144638 7732 144644 7744
rect 143040 7704 144644 7732
rect 143040 7692 143046 7704
rect 144638 7692 144644 7704
rect 144696 7692 144702 7744
rect 146036 7732 146064 7763
rect 146294 7732 146300 7744
rect 146036 7704 146300 7732
rect 146294 7692 146300 7704
rect 146352 7692 146358 7744
rect 146864 7732 146892 7772
rect 147122 7760 147128 7812
rect 147180 7800 147186 7812
rect 147416 7800 147444 7840
rect 147950 7828 147956 7840
rect 148008 7828 148014 7880
rect 148226 7868 148232 7880
rect 148139 7840 148232 7868
rect 148226 7828 148232 7840
rect 148284 7868 148290 7880
rect 148962 7868 148968 7880
rect 148284 7840 148968 7868
rect 148284 7828 148290 7840
rect 148962 7828 148968 7840
rect 149020 7828 149026 7880
rect 149072 7840 150296 7868
rect 148318 7800 148324 7812
rect 147180 7772 147444 7800
rect 147784 7772 148324 7800
rect 147180 7760 147186 7772
rect 147784 7732 147812 7772
rect 148318 7760 148324 7772
rect 148376 7760 148382 7812
rect 148496 7803 148554 7809
rect 148496 7769 148508 7803
rect 148542 7800 148554 7803
rect 148870 7800 148876 7812
rect 148542 7772 148876 7800
rect 148542 7769 148554 7772
rect 148496 7763 148554 7769
rect 148870 7760 148876 7772
rect 148928 7760 148934 7812
rect 146864 7704 147812 7732
rect 148134 7692 148140 7744
rect 148192 7732 148198 7744
rect 149072 7732 149100 7840
rect 149330 7760 149336 7812
rect 149388 7800 149394 7812
rect 150158 7800 150164 7812
rect 149388 7772 150164 7800
rect 149388 7760 149394 7772
rect 150158 7760 150164 7772
rect 150216 7760 150222 7812
rect 150268 7800 150296 7840
rect 150526 7828 150532 7880
rect 150584 7868 150590 7880
rect 150805 7871 150863 7877
rect 150805 7868 150817 7871
rect 150584 7840 150817 7868
rect 150584 7828 150590 7840
rect 150805 7837 150817 7840
rect 150851 7837 150863 7871
rect 150805 7831 150863 7837
rect 151081 7871 151139 7877
rect 151081 7837 151093 7871
rect 151127 7868 151139 7871
rect 151170 7868 151176 7880
rect 151127 7840 151176 7868
rect 151127 7837 151139 7840
rect 151081 7831 151139 7837
rect 151170 7828 151176 7840
rect 151228 7828 151234 7880
rect 152274 7868 152280 7880
rect 152235 7840 152280 7868
rect 152274 7828 152280 7840
rect 152332 7828 152338 7880
rect 152366 7828 152372 7880
rect 152424 7868 152430 7880
rect 152568 7868 152596 7908
rect 152918 7896 152924 7948
rect 152976 7936 152982 7948
rect 152976 7908 154620 7936
rect 152976 7896 152982 7908
rect 153565 7871 153623 7877
rect 153565 7868 153577 7871
rect 152424 7840 152469 7868
rect 152568 7840 153577 7868
rect 152424 7828 152430 7840
rect 153565 7837 153577 7840
rect 153611 7837 153623 7871
rect 153746 7868 153752 7880
rect 153707 7840 153752 7868
rect 153565 7831 153623 7837
rect 153746 7828 153752 7840
rect 153804 7828 153810 7880
rect 154022 7828 154028 7880
rect 154080 7868 154086 7880
rect 154485 7871 154543 7877
rect 154485 7868 154497 7871
rect 154080 7840 154497 7868
rect 154080 7828 154086 7840
rect 154485 7837 154497 7840
rect 154531 7837 154543 7871
rect 154592 7868 154620 7908
rect 155770 7896 155776 7948
rect 155828 7936 155834 7948
rect 156785 7939 156843 7945
rect 156785 7936 156797 7939
rect 155828 7908 156797 7936
rect 155828 7896 155834 7908
rect 156785 7905 156797 7908
rect 156831 7905 156843 7939
rect 156785 7899 156843 7905
rect 154741 7871 154799 7877
rect 154741 7868 154753 7871
rect 154592 7840 154753 7868
rect 154485 7831 154543 7837
rect 154741 7837 154753 7840
rect 154787 7868 154799 7871
rect 156046 7868 156052 7880
rect 154787 7840 156052 7868
rect 154787 7837 154799 7840
rect 154741 7831 154799 7837
rect 156046 7828 156052 7840
rect 156104 7828 156110 7880
rect 156598 7868 156604 7880
rect 156559 7840 156604 7868
rect 156598 7828 156604 7840
rect 156656 7828 156662 7880
rect 157429 7871 157487 7877
rect 157429 7837 157441 7871
rect 157475 7837 157487 7871
rect 157429 7831 157487 7837
rect 155494 7800 155500 7812
rect 150268 7772 155500 7800
rect 155494 7760 155500 7772
rect 155552 7760 155558 7812
rect 157444 7800 157472 7831
rect 155604 7772 157472 7800
rect 148192 7704 149100 7732
rect 149609 7735 149667 7741
rect 148192 7692 148198 7704
rect 149609 7701 149621 7735
rect 149655 7732 149667 7735
rect 151538 7732 151544 7744
rect 149655 7704 151544 7732
rect 149655 7701 149667 7704
rect 149609 7695 149667 7701
rect 151538 7692 151544 7704
rect 151596 7692 151602 7744
rect 151814 7692 151820 7744
rect 151872 7732 151878 7744
rect 152182 7732 152188 7744
rect 151872 7704 152188 7732
rect 151872 7692 151878 7704
rect 152182 7692 152188 7704
rect 152240 7692 152246 7744
rect 153378 7732 153384 7744
rect 153339 7704 153384 7732
rect 153378 7692 153384 7704
rect 153436 7692 153442 7744
rect 154022 7692 154028 7744
rect 154080 7732 154086 7744
rect 155604 7732 155632 7772
rect 155862 7732 155868 7744
rect 154080 7704 155632 7732
rect 155823 7704 155868 7732
rect 154080 7692 154086 7704
rect 155862 7692 155868 7704
rect 155920 7692 155926 7744
rect 156138 7692 156144 7744
rect 156196 7732 156202 7744
rect 156417 7735 156475 7741
rect 156417 7732 156429 7735
rect 156196 7704 156429 7732
rect 156196 7692 156202 7704
rect 156417 7701 156429 7704
rect 156463 7701 156475 7735
rect 156417 7695 156475 7701
rect 157518 7692 157524 7744
rect 157576 7732 157582 7744
rect 157981 7735 158039 7741
rect 157981 7732 157993 7735
rect 157576 7704 157993 7732
rect 157576 7692 157582 7704
rect 157981 7701 157993 7704
rect 158027 7732 158039 7735
rect 158254 7732 158260 7744
rect 158027 7704 158260 7732
rect 158027 7701 158039 7704
rect 157981 7695 158039 7701
rect 158254 7692 158260 7704
rect 158312 7692 158318 7744
rect 1104 7642 159043 7664
rect 1104 7590 40394 7642
rect 40446 7590 40458 7642
rect 40510 7590 40522 7642
rect 40574 7590 40586 7642
rect 40638 7590 40650 7642
rect 40702 7590 79839 7642
rect 79891 7590 79903 7642
rect 79955 7590 79967 7642
rect 80019 7590 80031 7642
rect 80083 7590 80095 7642
rect 80147 7590 119284 7642
rect 119336 7590 119348 7642
rect 119400 7590 119412 7642
rect 119464 7590 119476 7642
rect 119528 7590 119540 7642
rect 119592 7590 158729 7642
rect 158781 7590 158793 7642
rect 158845 7590 158857 7642
rect 158909 7590 158921 7642
rect 158973 7590 158985 7642
rect 159037 7590 159043 7642
rect 1104 7568 159043 7590
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5994 7528 6000 7540
rect 5907 7500 6000 7528
rect 5994 7488 6000 7500
rect 6052 7528 6058 7540
rect 6730 7528 6736 7540
rect 6052 7500 6736 7528
rect 6052 7488 6058 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 14090 7528 14096 7540
rect 14051 7500 14096 7528
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 15102 7528 15108 7540
rect 15063 7500 15108 7528
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 15160 7500 16865 7528
rect 15160 7488 15166 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 21082 7528 21088 7540
rect 21043 7500 21088 7528
rect 16853 7491 16911 7497
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 23290 7488 23296 7540
rect 23348 7528 23354 7540
rect 32858 7528 32864 7540
rect 23348 7500 31754 7528
rect 32819 7500 32864 7528
rect 23348 7488 23354 7500
rect 15749 7463 15807 7469
rect 15749 7429 15761 7463
rect 15795 7460 15807 7463
rect 16390 7460 16396 7472
rect 15795 7432 16396 7460
rect 15795 7429 15807 7432
rect 15749 7423 15807 7429
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 18598 7460 18604 7472
rect 18064 7432 18604 7460
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5132 7364 5457 7392
rect 5132 7352 5138 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 5445 7355 5503 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13679 7364 14289 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16850 7392 16856 7404
rect 16347 7364 16856 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 17862 7392 17868 7404
rect 17451 7364 17868 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 11204 7296 12817 7324
rect 11204 7284 11210 7296
rect 12805 7293 12817 7296
rect 12851 7324 12863 7327
rect 13265 7327 13323 7333
rect 13265 7324 13277 7327
rect 12851 7296 13277 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13265 7293 13277 7296
rect 13311 7293 13323 7327
rect 13265 7287 13323 7293
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 18064 7333 18092 7432
rect 18598 7420 18604 7432
rect 18656 7420 18662 7472
rect 30101 7463 30159 7469
rect 30101 7460 30113 7463
rect 29288 7432 30113 7460
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21634 7392 21640 7404
rect 21315 7364 21640 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17828 7296 18061 7324
rect 17828 7284 17834 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 15838 7256 15844 7268
rect 12768 7228 15844 7256
rect 12768 7216 12774 7228
rect 15838 7216 15844 7228
rect 15896 7216 15902 7268
rect 18248 7256 18276 7355
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21818 7352 21824 7404
rect 21876 7392 21882 7404
rect 26062 7395 26120 7401
rect 26062 7392 26074 7395
rect 21876 7364 26074 7392
rect 21876 7352 21882 7364
rect 26062 7361 26074 7364
rect 26108 7361 26120 7395
rect 26062 7355 26120 7361
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 29288 7401 29316 7432
rect 30101 7429 30113 7432
rect 30147 7460 30159 7463
rect 30558 7460 30564 7472
rect 30147 7432 30564 7460
rect 30147 7429 30159 7432
rect 30101 7423 30159 7429
rect 30558 7420 30564 7432
rect 30616 7460 30622 7472
rect 31018 7460 31024 7472
rect 30616 7432 31024 7460
rect 30616 7420 30622 7432
rect 31018 7420 31024 7432
rect 31076 7460 31082 7472
rect 31113 7463 31171 7469
rect 31113 7460 31125 7463
rect 31076 7432 31125 7460
rect 31076 7420 31082 7432
rect 31113 7429 31125 7432
rect 31159 7429 31171 7463
rect 31726 7460 31754 7500
rect 32858 7488 32864 7500
rect 32916 7488 32922 7540
rect 34701 7531 34759 7537
rect 34701 7497 34713 7531
rect 34747 7497 34759 7531
rect 34701 7491 34759 7497
rect 36725 7531 36783 7537
rect 36725 7497 36737 7531
rect 36771 7497 36783 7531
rect 38562 7528 38568 7540
rect 38523 7500 38568 7528
rect 36725 7491 36783 7497
rect 32401 7463 32459 7469
rect 31726 7432 32352 7460
rect 31113 7423 31171 7429
rect 29273 7395 29331 7401
rect 29273 7392 29285 7395
rect 26660 7364 29285 7392
rect 26660 7352 26666 7364
rect 29273 7361 29285 7364
rect 29319 7361 29331 7395
rect 29273 7355 29331 7361
rect 29457 7395 29515 7401
rect 29457 7361 29469 7395
rect 29503 7361 29515 7395
rect 32324 7392 32352 7432
rect 32401 7429 32413 7463
rect 32447 7460 32459 7463
rect 33778 7460 33784 7472
rect 32447 7432 33784 7460
rect 32447 7429 32459 7432
rect 32401 7423 32459 7429
rect 33778 7420 33784 7432
rect 33836 7420 33842 7472
rect 34716 7460 34744 7491
rect 33888 7432 34744 7460
rect 36740 7460 36768 7491
rect 38562 7488 38568 7500
rect 38620 7488 38626 7540
rect 40310 7488 40316 7540
rect 40368 7528 40374 7540
rect 40497 7531 40555 7537
rect 40497 7528 40509 7531
rect 40368 7500 40509 7528
rect 40368 7488 40374 7500
rect 40497 7497 40509 7500
rect 40543 7497 40555 7531
rect 40497 7491 40555 7497
rect 41417 7531 41475 7537
rect 41417 7497 41429 7531
rect 41463 7497 41475 7531
rect 41417 7491 41475 7497
rect 41969 7531 42027 7537
rect 41969 7497 41981 7531
rect 42015 7528 42027 7531
rect 42058 7528 42064 7540
rect 42015 7500 42064 7528
rect 42015 7497 42027 7500
rect 41969 7491 42027 7497
rect 39362 7463 39420 7469
rect 39362 7460 39374 7463
rect 36740 7432 39374 7460
rect 33888 7392 33916 7432
rect 39362 7429 39374 7432
rect 39408 7429 39420 7463
rect 41432 7460 41460 7491
rect 42058 7488 42064 7500
rect 42116 7488 42122 7540
rect 43073 7531 43131 7537
rect 43073 7497 43085 7531
rect 43119 7528 43131 7531
rect 43162 7528 43168 7540
rect 43119 7500 43168 7528
rect 43119 7497 43131 7500
rect 43073 7491 43131 7497
rect 43162 7488 43168 7500
rect 43220 7488 43226 7540
rect 45189 7531 45247 7537
rect 45189 7497 45201 7531
rect 45235 7528 45247 7531
rect 45370 7528 45376 7540
rect 45235 7500 45376 7528
rect 45235 7497 45247 7500
rect 45189 7491 45247 7497
rect 45370 7488 45376 7500
rect 45428 7488 45434 7540
rect 49329 7531 49387 7537
rect 49329 7497 49341 7531
rect 49375 7528 49387 7531
rect 49602 7528 49608 7540
rect 49375 7500 49608 7528
rect 49375 7497 49387 7500
rect 49329 7491 49387 7497
rect 49602 7488 49608 7500
rect 49660 7488 49666 7540
rect 49786 7488 49792 7540
rect 49844 7528 49850 7540
rect 50433 7531 50491 7537
rect 50433 7528 50445 7531
rect 49844 7500 50445 7528
rect 49844 7488 49850 7500
rect 50433 7497 50445 7500
rect 50479 7528 50491 7531
rect 57425 7531 57483 7537
rect 57425 7528 57437 7531
rect 50479 7500 57437 7528
rect 50479 7497 50491 7500
rect 50433 7491 50491 7497
rect 57425 7497 57437 7500
rect 57471 7528 57483 7531
rect 57698 7528 57704 7540
rect 57471 7500 57704 7528
rect 57471 7497 57483 7500
rect 57425 7491 57483 7497
rect 57698 7488 57704 7500
rect 57756 7488 57762 7540
rect 57790 7488 57796 7540
rect 57848 7528 57854 7540
rect 58069 7531 58127 7537
rect 58069 7528 58081 7531
rect 57848 7500 58081 7528
rect 57848 7488 57854 7500
rect 58069 7497 58081 7500
rect 58115 7497 58127 7531
rect 58069 7491 58127 7497
rect 58526 7488 58532 7540
rect 58584 7528 58590 7540
rect 58713 7531 58771 7537
rect 58713 7528 58725 7531
rect 58584 7500 58725 7528
rect 58584 7488 58590 7500
rect 58713 7497 58725 7500
rect 58759 7528 58771 7531
rect 59170 7528 59176 7540
rect 58759 7500 59176 7528
rect 58759 7497 58771 7500
rect 58713 7491 58771 7497
rect 59170 7488 59176 7500
rect 59228 7488 59234 7540
rect 59722 7528 59728 7540
rect 59683 7500 59728 7528
rect 59722 7488 59728 7500
rect 59780 7488 59786 7540
rect 63218 7528 63224 7540
rect 63179 7500 63224 7528
rect 63218 7488 63224 7500
rect 63276 7488 63282 7540
rect 64782 7528 64788 7540
rect 64743 7500 64788 7528
rect 64782 7488 64788 7500
rect 64840 7488 64846 7540
rect 65242 7528 65248 7540
rect 65203 7500 65248 7528
rect 65242 7488 65248 7500
rect 65300 7488 65306 7540
rect 67082 7528 67088 7540
rect 67043 7500 67088 7528
rect 67082 7488 67088 7500
rect 67140 7488 67146 7540
rect 71593 7531 71651 7537
rect 71593 7528 71605 7531
rect 70366 7500 71605 7528
rect 45554 7460 45560 7472
rect 41432 7432 45560 7460
rect 39362 7423 39420 7429
rect 45554 7420 45560 7432
rect 45612 7420 45618 7472
rect 45830 7420 45836 7472
rect 45888 7460 45894 7472
rect 46477 7463 46535 7469
rect 46477 7460 46489 7463
rect 45888 7432 46489 7460
rect 45888 7420 45894 7432
rect 46477 7429 46489 7432
rect 46523 7460 46535 7463
rect 49510 7460 49516 7472
rect 46523 7432 49516 7460
rect 46523 7429 46535 7432
rect 46477 7423 46535 7429
rect 49510 7420 49516 7432
rect 49568 7420 49574 7472
rect 52120 7463 52178 7469
rect 52120 7429 52132 7463
rect 52166 7460 52178 7463
rect 54754 7460 54760 7472
rect 52166 7432 54760 7460
rect 52166 7429 52178 7432
rect 52120 7423 52178 7429
rect 54754 7420 54760 7432
rect 54812 7420 54818 7472
rect 64230 7420 64236 7472
rect 64288 7460 64294 7472
rect 66073 7463 66131 7469
rect 66073 7460 66085 7463
rect 64288 7432 66085 7460
rect 64288 7420 64294 7432
rect 66073 7429 66085 7432
rect 66119 7429 66131 7463
rect 66073 7423 66131 7429
rect 32324 7364 33916 7392
rect 29457 7355 29515 7361
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 23934 7324 23940 7336
rect 18463 7296 23940 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 26326 7324 26332 7336
rect 26287 7296 26332 7324
rect 26326 7284 26332 7296
rect 26384 7284 26390 7336
rect 18874 7256 18880 7268
rect 18248 7228 18880 7256
rect 18874 7216 18880 7228
rect 18932 7256 18938 7268
rect 18932 7228 19012 7256
rect 18932 7216 18938 7228
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 17589 7191 17647 7197
rect 17589 7157 17601 7191
rect 17635 7188 17647 7191
rect 18322 7188 18328 7200
rect 17635 7160 18328 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 18984 7197 19012 7228
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 24949 7259 25007 7265
rect 24949 7256 24961 7259
rect 19208 7228 24961 7256
rect 19208 7216 19214 7228
rect 24949 7225 24961 7228
rect 24995 7225 25007 7259
rect 29472 7256 29500 7355
rect 33962 7352 33968 7404
rect 34020 7401 34026 7404
rect 34020 7392 34032 7401
rect 34238 7392 34244 7404
rect 34020 7364 34065 7392
rect 34199 7364 34244 7392
rect 34020 7355 34032 7364
rect 34020 7352 34026 7355
rect 34238 7352 34244 7364
rect 34296 7352 34302 7404
rect 34882 7352 34888 7404
rect 34940 7392 34946 7404
rect 35814 7395 35872 7401
rect 35814 7392 35826 7395
rect 34940 7364 35826 7392
rect 34940 7352 34946 7364
rect 35814 7361 35826 7364
rect 35860 7361 35872 7395
rect 35814 7355 35872 7361
rect 36446 7352 36452 7404
rect 36504 7392 36510 7404
rect 36541 7395 36599 7401
rect 36541 7392 36553 7395
rect 36504 7364 36553 7392
rect 36504 7352 36510 7364
rect 36541 7361 36553 7364
rect 36587 7361 36599 7395
rect 36541 7355 36599 7361
rect 37826 7352 37832 7404
rect 37884 7392 37890 7404
rect 40770 7392 40776 7404
rect 37884 7364 40776 7392
rect 37884 7352 37890 7364
rect 40770 7352 40776 7364
rect 40828 7392 40834 7404
rect 41230 7392 41236 7404
rect 40828 7364 41000 7392
rect 41191 7364 41236 7392
rect 40828 7352 40834 7364
rect 29641 7327 29699 7333
rect 29641 7293 29653 7327
rect 29687 7324 29699 7327
rect 33134 7324 33140 7336
rect 29687 7296 33140 7324
rect 29687 7293 29699 7296
rect 29641 7287 29699 7293
rect 33134 7284 33140 7296
rect 33192 7284 33198 7336
rect 36081 7327 36139 7333
rect 36081 7293 36093 7327
rect 36127 7324 36139 7327
rect 37182 7324 37188 7336
rect 36127 7296 37188 7324
rect 36127 7293 36139 7296
rect 36081 7287 36139 7293
rect 37182 7284 37188 7296
rect 37240 7284 37246 7336
rect 38013 7327 38071 7333
rect 38013 7293 38025 7327
rect 38059 7324 38071 7327
rect 38470 7324 38476 7336
rect 38059 7296 38476 7324
rect 38059 7293 38071 7296
rect 38013 7287 38071 7293
rect 38470 7284 38476 7296
rect 38528 7324 38534 7336
rect 39117 7327 39175 7333
rect 39117 7324 39129 7327
rect 38528 7296 39129 7324
rect 38528 7284 38534 7296
rect 39117 7293 39129 7296
rect 39163 7293 39175 7327
rect 40972 7324 41000 7364
rect 41230 7352 41236 7364
rect 41288 7352 41294 7404
rect 42426 7352 42432 7404
rect 42484 7392 42490 7404
rect 49694 7392 49700 7404
rect 42484 7364 49700 7392
rect 42484 7352 42490 7364
rect 49694 7352 49700 7364
rect 49752 7352 49758 7404
rect 53098 7352 53104 7404
rect 53156 7392 53162 7404
rect 53193 7395 53251 7401
rect 53193 7392 53205 7395
rect 53156 7364 53205 7392
rect 53156 7352 53162 7364
rect 53193 7361 53205 7364
rect 53239 7361 53251 7395
rect 53834 7392 53840 7404
rect 53795 7364 53840 7392
rect 53193 7355 53251 7361
rect 53834 7352 53840 7364
rect 53892 7352 53898 7404
rect 54294 7352 54300 7404
rect 54352 7392 54358 7404
rect 54849 7395 54907 7401
rect 54849 7392 54861 7395
rect 54352 7364 54861 7392
rect 54352 7352 54358 7364
rect 54849 7361 54861 7364
rect 54895 7361 54907 7395
rect 54849 7355 54907 7361
rect 58253 7395 58311 7401
rect 58253 7361 58265 7395
rect 58299 7392 58311 7395
rect 59998 7392 60004 7404
rect 58299 7364 60004 7392
rect 58299 7361 58311 7364
rect 58253 7355 58311 7361
rect 59998 7352 60004 7364
rect 60056 7352 60062 7404
rect 60550 7392 60556 7404
rect 60511 7364 60556 7392
rect 60550 7352 60556 7364
rect 60608 7352 60614 7404
rect 61562 7352 61568 7404
rect 61620 7392 61626 7404
rect 63402 7392 63408 7404
rect 61620 7364 62804 7392
rect 63363 7364 63408 7392
rect 61620 7352 61626 7364
rect 45830 7324 45836 7336
rect 40972 7296 45836 7324
rect 39117 7287 39175 7293
rect 45830 7284 45836 7296
rect 45888 7284 45894 7336
rect 52362 7284 52368 7336
rect 52420 7324 52426 7336
rect 62577 7327 62635 7333
rect 62577 7324 62589 7327
rect 52420 7296 62589 7324
rect 52420 7284 52426 7296
rect 62577 7293 62589 7296
rect 62623 7324 62635 7327
rect 62666 7324 62672 7336
rect 62623 7296 62672 7324
rect 62623 7293 62635 7296
rect 62577 7287 62635 7293
rect 62666 7284 62672 7296
rect 62724 7284 62730 7336
rect 62776 7324 62804 7364
rect 63402 7352 63408 7364
rect 63460 7352 63466 7404
rect 64598 7392 64604 7404
rect 64559 7364 64604 7392
rect 64598 7352 64604 7364
rect 64656 7352 64662 7404
rect 66901 7395 66959 7401
rect 66901 7361 66913 7395
rect 66947 7392 66959 7395
rect 66990 7392 66996 7404
rect 66947 7364 66996 7392
rect 66947 7361 66959 7364
rect 66901 7355 66959 7361
rect 66990 7352 66996 7364
rect 67048 7352 67054 7404
rect 70366 7324 70394 7500
rect 71593 7497 71605 7500
rect 71639 7528 71651 7531
rect 73614 7528 73620 7540
rect 71639 7500 73620 7528
rect 71639 7497 71651 7500
rect 71593 7491 71651 7497
rect 73614 7488 73620 7500
rect 73672 7488 73678 7540
rect 74077 7531 74135 7537
rect 74077 7497 74089 7531
rect 74123 7528 74135 7531
rect 74718 7528 74724 7540
rect 74123 7500 74724 7528
rect 74123 7497 74135 7500
rect 74077 7491 74135 7497
rect 74718 7488 74724 7500
rect 74776 7488 74782 7540
rect 76561 7531 76619 7537
rect 76561 7528 76573 7531
rect 76484 7500 76573 7528
rect 72717 7395 72775 7401
rect 72717 7361 72729 7395
rect 72763 7392 72775 7395
rect 72878 7392 72884 7404
rect 72763 7364 72884 7392
rect 72763 7361 72775 7364
rect 72717 7355 72775 7361
rect 72878 7352 72884 7364
rect 72936 7352 72942 7404
rect 75201 7395 75259 7401
rect 75201 7361 75213 7395
rect 75247 7392 75259 7395
rect 76484 7392 76512 7500
rect 76561 7497 76573 7500
rect 76607 7528 76619 7531
rect 76607 7500 84884 7528
rect 76607 7497 76619 7500
rect 76561 7491 76619 7497
rect 79312 7463 79370 7469
rect 79312 7429 79324 7463
rect 79358 7460 79370 7463
rect 83458 7460 83464 7472
rect 79358 7432 83464 7460
rect 79358 7429 79370 7432
rect 79312 7423 79370 7429
rect 83458 7420 83464 7432
rect 83516 7420 83522 7472
rect 84856 7460 84884 7500
rect 85298 7488 85304 7540
rect 85356 7528 85362 7540
rect 86218 7528 86224 7540
rect 85356 7500 86224 7528
rect 85356 7488 85362 7500
rect 86218 7488 86224 7500
rect 86276 7488 86282 7540
rect 93486 7488 93492 7540
rect 93544 7528 93550 7540
rect 96890 7528 96896 7540
rect 93544 7500 96896 7528
rect 93544 7488 93550 7500
rect 96890 7488 96896 7500
rect 96948 7488 96954 7540
rect 97350 7528 97356 7540
rect 97311 7500 97356 7528
rect 97350 7488 97356 7500
rect 97408 7488 97414 7540
rect 97442 7488 97448 7540
rect 97500 7528 97506 7540
rect 108850 7528 108856 7540
rect 97500 7500 108856 7528
rect 97500 7488 97506 7500
rect 108850 7488 108856 7500
rect 108908 7488 108914 7540
rect 116762 7528 116768 7540
rect 109006 7500 116768 7528
rect 89346 7460 89352 7472
rect 84856 7432 89352 7460
rect 89346 7420 89352 7432
rect 89404 7420 89410 7472
rect 89806 7420 89812 7472
rect 89864 7460 89870 7472
rect 109006 7460 109034 7500
rect 116762 7488 116768 7500
rect 116820 7488 116826 7540
rect 127161 7531 127219 7537
rect 127161 7528 127173 7531
rect 117424 7500 127173 7528
rect 110598 7460 110604 7472
rect 89864 7432 109034 7460
rect 110524 7432 110604 7460
rect 89864 7420 89870 7432
rect 75247 7364 76512 7392
rect 81428 7395 81486 7401
rect 75247 7361 75259 7364
rect 75201 7355 75259 7361
rect 81428 7361 81440 7395
rect 81474 7392 81486 7395
rect 83090 7392 83096 7404
rect 81474 7364 83096 7392
rect 81474 7361 81486 7364
rect 81428 7355 81486 7361
rect 83090 7352 83096 7364
rect 83148 7352 83154 7404
rect 84654 7392 84660 7404
rect 84615 7364 84660 7392
rect 84654 7352 84660 7364
rect 84712 7352 84718 7404
rect 90818 7392 90824 7404
rect 84764 7364 90824 7392
rect 62776 7296 70394 7324
rect 72973 7327 73031 7333
rect 72973 7293 72985 7327
rect 73019 7324 73031 7327
rect 73154 7324 73160 7336
rect 73019 7296 73160 7324
rect 73019 7293 73031 7296
rect 72973 7287 73031 7293
rect 73154 7284 73160 7296
rect 73212 7284 73218 7336
rect 75457 7327 75515 7333
rect 75457 7293 75469 7327
rect 75503 7324 75515 7327
rect 75914 7324 75920 7336
rect 75503 7296 75920 7324
rect 75503 7293 75515 7296
rect 75457 7287 75515 7293
rect 75914 7284 75920 7296
rect 75972 7284 75978 7336
rect 79042 7324 79048 7336
rect 79003 7296 79048 7324
rect 79042 7284 79048 7296
rect 79100 7284 79106 7336
rect 81066 7284 81072 7336
rect 81124 7324 81130 7336
rect 81161 7327 81219 7333
rect 81161 7324 81173 7327
rect 81124 7296 81173 7324
rect 81124 7284 81130 7296
rect 81161 7293 81173 7296
rect 81207 7293 81219 7327
rect 84764 7324 84792 7364
rect 90818 7352 90824 7364
rect 90876 7352 90882 7404
rect 90910 7352 90916 7404
rect 90968 7392 90974 7404
rect 91557 7395 91615 7401
rect 91557 7392 91569 7395
rect 90968 7364 91569 7392
rect 90968 7352 90974 7364
rect 91557 7361 91569 7364
rect 91603 7361 91615 7395
rect 91557 7355 91615 7361
rect 91824 7395 91882 7401
rect 91824 7361 91836 7395
rect 91870 7392 91882 7395
rect 93486 7392 93492 7404
rect 91870 7364 93492 7392
rect 91870 7361 91882 7364
rect 91824 7355 91882 7361
rect 93486 7352 93492 7364
rect 93544 7352 93550 7404
rect 96522 7352 96528 7404
rect 96580 7401 96586 7404
rect 96580 7392 96592 7401
rect 96798 7392 96804 7404
rect 96580 7364 96625 7392
rect 96711 7364 96804 7392
rect 96580 7355 96592 7364
rect 96580 7352 96586 7355
rect 96798 7352 96804 7364
rect 96856 7392 96862 7404
rect 97350 7392 97356 7404
rect 96856 7364 97356 7392
rect 96856 7352 96862 7364
rect 97350 7352 97356 7364
rect 97408 7352 97414 7404
rect 110524 7401 110552 7432
rect 110598 7420 110604 7432
rect 110656 7420 110662 7472
rect 111610 7469 111616 7472
rect 111604 7423 111616 7469
rect 111668 7460 111674 7472
rect 111668 7432 111704 7460
rect 111610 7420 111616 7423
rect 111668 7420 111674 7432
rect 110509 7395 110567 7401
rect 110509 7361 110521 7395
rect 110555 7361 110567 7395
rect 110690 7392 110696 7404
rect 110651 7364 110696 7392
rect 110509 7355 110567 7361
rect 110690 7352 110696 7364
rect 110748 7352 110754 7404
rect 114094 7392 114100 7404
rect 114055 7364 114100 7392
rect 114094 7352 114100 7364
rect 114152 7352 114158 7404
rect 116765 7395 116823 7401
rect 116765 7361 116777 7395
rect 116811 7392 116823 7395
rect 116946 7392 116952 7404
rect 116811 7364 116952 7392
rect 116811 7361 116823 7364
rect 116765 7355 116823 7361
rect 116946 7352 116952 7364
rect 117004 7392 117010 7404
rect 117225 7395 117283 7401
rect 117225 7392 117237 7395
rect 117004 7364 117237 7392
rect 117004 7352 117010 7364
rect 117225 7361 117237 7364
rect 117271 7361 117283 7395
rect 117225 7355 117283 7361
rect 81161 7287 81219 7293
rect 82464 7296 84792 7324
rect 42886 7256 42892 7268
rect 29472 7228 33364 7256
rect 24949 7219 25007 7225
rect 18969 7191 19027 7197
rect 18969 7157 18981 7191
rect 19015 7188 19027 7191
rect 19242 7188 19248 7200
rect 19015 7160 19248 7188
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 22097 7191 22155 7197
rect 22097 7157 22109 7191
rect 22143 7188 22155 7191
rect 22554 7188 22560 7200
rect 22143 7160 22560 7188
rect 22143 7157 22155 7160
rect 22097 7151 22155 7157
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 33336 7188 33364 7228
rect 41386 7228 42892 7256
rect 35342 7188 35348 7200
rect 33336 7160 35348 7188
rect 35342 7148 35348 7160
rect 35400 7188 35406 7200
rect 41386 7188 41414 7228
rect 42886 7216 42892 7228
rect 42944 7216 42950 7268
rect 50798 7216 50804 7268
rect 50856 7256 50862 7268
rect 50985 7259 51043 7265
rect 50985 7256 50997 7259
rect 50856 7228 50997 7256
rect 50856 7216 50862 7228
rect 50985 7225 50997 7228
rect 51031 7225 51043 7259
rect 50985 7219 51043 7225
rect 60826 7216 60832 7268
rect 60884 7256 60890 7268
rect 82464 7256 82492 7296
rect 86218 7284 86224 7336
rect 86276 7324 86282 7336
rect 86276 7296 91600 7324
rect 86276 7284 86282 7296
rect 82541 7259 82599 7265
rect 82541 7256 82553 7259
rect 60884 7228 70394 7256
rect 60884 7216 60890 7228
rect 35400 7160 41414 7188
rect 35400 7148 35406 7160
rect 44358 7148 44364 7200
rect 44416 7188 44422 7200
rect 45738 7188 45744 7200
rect 44416 7160 45744 7188
rect 44416 7148 44422 7160
rect 45738 7148 45744 7160
rect 45796 7188 45802 7200
rect 45833 7191 45891 7197
rect 45833 7188 45845 7191
rect 45796 7160 45845 7188
rect 45796 7148 45802 7160
rect 45833 7157 45845 7160
rect 45879 7188 45891 7191
rect 47026 7188 47032 7200
rect 45879 7160 47032 7188
rect 45879 7157 45891 7160
rect 45833 7151 45891 7157
rect 47026 7148 47032 7160
rect 47084 7148 47090 7200
rect 60737 7191 60795 7197
rect 60737 7157 60749 7191
rect 60783 7188 60795 7191
rect 61102 7188 61108 7200
rect 60783 7160 61108 7188
rect 60783 7157 60795 7160
rect 60737 7151 60795 7157
rect 61102 7148 61108 7160
rect 61160 7148 61166 7200
rect 68370 7188 68376 7200
rect 68331 7160 68376 7188
rect 68370 7148 68376 7160
rect 68428 7148 68434 7200
rect 70366 7188 70394 7228
rect 80256 7228 80560 7256
rect 82464 7228 82553 7256
rect 80256 7188 80284 7228
rect 80422 7188 80428 7200
rect 70366 7160 80284 7188
rect 80383 7160 80428 7188
rect 80422 7148 80428 7160
rect 80480 7148 80486 7200
rect 80532 7188 80560 7228
rect 82541 7225 82553 7228
rect 82587 7225 82599 7259
rect 82541 7219 82599 7225
rect 82630 7216 82636 7268
rect 82688 7256 82694 7268
rect 82688 7228 89714 7256
rect 82688 7216 82694 7228
rect 82446 7188 82452 7200
rect 80532 7160 82452 7188
rect 82446 7148 82452 7160
rect 82504 7148 82510 7200
rect 83090 7188 83096 7200
rect 83051 7160 83096 7188
rect 83090 7148 83096 7160
rect 83148 7148 83154 7200
rect 83642 7148 83648 7200
rect 83700 7188 83706 7200
rect 84473 7191 84531 7197
rect 84473 7188 84485 7191
rect 83700 7160 84485 7188
rect 83700 7148 83706 7160
rect 84473 7157 84485 7160
rect 84519 7157 84531 7191
rect 84473 7151 84531 7157
rect 85574 7148 85580 7200
rect 85632 7188 85638 7200
rect 86037 7191 86095 7197
rect 86037 7188 86049 7191
rect 85632 7160 86049 7188
rect 85632 7148 85638 7160
rect 86037 7157 86049 7160
rect 86083 7188 86095 7191
rect 86402 7188 86408 7200
rect 86083 7160 86408 7188
rect 86083 7157 86095 7160
rect 86037 7151 86095 7157
rect 86402 7148 86408 7160
rect 86460 7148 86466 7200
rect 86770 7148 86776 7200
rect 86828 7188 86834 7200
rect 87233 7191 87291 7197
rect 87233 7188 87245 7191
rect 86828 7160 87245 7188
rect 86828 7148 86834 7160
rect 87233 7157 87245 7160
rect 87279 7188 87291 7191
rect 87690 7188 87696 7200
rect 87279 7160 87696 7188
rect 87279 7157 87291 7160
rect 87233 7151 87291 7157
rect 87690 7148 87696 7160
rect 87748 7148 87754 7200
rect 89686 7188 89714 7228
rect 91370 7188 91376 7200
rect 89686 7160 91376 7188
rect 91370 7148 91376 7160
rect 91428 7148 91434 7200
rect 91572 7188 91600 7296
rect 92584 7296 95556 7324
rect 92584 7188 92612 7296
rect 91572 7160 92612 7188
rect 92934 7148 92940 7200
rect 92992 7188 92998 7200
rect 93486 7188 93492 7200
rect 92992 7160 93037 7188
rect 93447 7160 93492 7188
rect 92992 7148 92998 7160
rect 93486 7148 93492 7160
rect 93544 7148 93550 7200
rect 93578 7148 93584 7200
rect 93636 7188 93642 7200
rect 95421 7191 95479 7197
rect 95421 7188 95433 7191
rect 93636 7160 95433 7188
rect 93636 7148 93642 7160
rect 95421 7157 95433 7160
rect 95467 7157 95479 7191
rect 95528 7188 95556 7296
rect 96890 7284 96896 7336
rect 96948 7324 96954 7336
rect 99190 7324 99196 7336
rect 96948 7296 99196 7324
rect 96948 7284 96954 7296
rect 99190 7284 99196 7296
rect 99248 7284 99254 7336
rect 107010 7284 107016 7336
rect 107068 7324 107074 7336
rect 110877 7327 110935 7333
rect 107068 7296 110460 7324
rect 107068 7284 107074 7296
rect 96982 7216 96988 7268
rect 97040 7256 97046 7268
rect 110322 7256 110328 7268
rect 97040 7228 110328 7256
rect 97040 7216 97046 7228
rect 110322 7216 110328 7228
rect 110380 7216 110386 7268
rect 97442 7188 97448 7200
rect 95528 7160 97448 7188
rect 95421 7151 95479 7157
rect 97442 7148 97448 7160
rect 97500 7148 97506 7200
rect 97534 7148 97540 7200
rect 97592 7188 97598 7200
rect 109862 7188 109868 7200
rect 97592 7160 109868 7188
rect 97592 7148 97598 7160
rect 109862 7148 109868 7160
rect 109920 7148 109926 7200
rect 110046 7188 110052 7200
rect 110007 7160 110052 7188
rect 110046 7148 110052 7160
rect 110104 7148 110110 7200
rect 110432 7188 110460 7296
rect 110877 7293 110889 7327
rect 110923 7324 110935 7327
rect 110966 7324 110972 7336
rect 110923 7296 110972 7324
rect 110923 7293 110935 7296
rect 110877 7287 110935 7293
rect 110966 7284 110972 7296
rect 111024 7284 111030 7336
rect 111334 7324 111340 7336
rect 111295 7296 111340 7324
rect 111334 7284 111340 7296
rect 111392 7284 111398 7336
rect 112438 7284 112444 7336
rect 112496 7324 112502 7336
rect 112898 7324 112904 7336
rect 112496 7296 112904 7324
rect 112496 7284 112502 7296
rect 112898 7284 112904 7296
rect 112956 7324 112962 7336
rect 113177 7327 113235 7333
rect 113177 7324 113189 7327
rect 112956 7296 113189 7324
rect 112956 7284 112962 7296
rect 113177 7293 113189 7296
rect 113223 7293 113235 7327
rect 113177 7287 113235 7293
rect 113266 7284 113272 7336
rect 113324 7324 113330 7336
rect 117424 7324 117452 7500
rect 118418 7420 118424 7472
rect 118476 7460 118482 7472
rect 122938 7463 122996 7469
rect 122938 7460 122950 7463
rect 118476 7432 122950 7460
rect 118476 7420 118482 7432
rect 122938 7429 122950 7432
rect 122984 7429 122996 7463
rect 122938 7423 122996 7429
rect 123110 7420 123116 7472
rect 123168 7460 123174 7472
rect 124398 7460 124404 7472
rect 123168 7432 124404 7460
rect 123168 7420 123174 7432
rect 124398 7420 124404 7432
rect 124456 7420 124462 7472
rect 125410 7420 125416 7472
rect 125468 7460 125474 7472
rect 126330 7460 126336 7472
rect 125468 7432 126336 7460
rect 125468 7420 125474 7432
rect 126330 7420 126336 7432
rect 126388 7420 126394 7472
rect 119062 7392 119068 7404
rect 119120 7401 119126 7404
rect 119120 7395 119143 7401
rect 118995 7364 119068 7392
rect 119062 7352 119068 7364
rect 119131 7392 119143 7395
rect 121109 7395 121167 7401
rect 119131 7364 120396 7392
rect 119131 7361 119143 7364
rect 119120 7355 119143 7361
rect 119120 7352 119126 7355
rect 113324 7296 117452 7324
rect 119341 7327 119399 7333
rect 113324 7284 113330 7296
rect 119341 7293 119353 7327
rect 119387 7293 119399 7327
rect 119341 7287 119399 7293
rect 117961 7259 118019 7265
rect 117961 7256 117973 7259
rect 112272 7228 117973 7256
rect 112272 7188 112300 7228
rect 117961 7225 117973 7228
rect 118007 7225 118019 7259
rect 117961 7219 118019 7225
rect 112714 7188 112720 7200
rect 110432 7160 112300 7188
rect 112675 7160 112720 7188
rect 112714 7148 112720 7160
rect 112772 7148 112778 7200
rect 112898 7148 112904 7200
rect 112956 7188 112962 7200
rect 113913 7191 113971 7197
rect 113913 7188 113925 7191
rect 112956 7160 113925 7188
rect 112956 7148 112962 7160
rect 113913 7157 113925 7160
rect 113959 7157 113971 7191
rect 113913 7151 113971 7157
rect 114922 7148 114928 7200
rect 114980 7188 114986 7200
rect 117406 7188 117412 7200
rect 114980 7160 117412 7188
rect 114980 7148 114986 7160
rect 117406 7148 117412 7160
rect 117464 7148 117470 7200
rect 118970 7148 118976 7200
rect 119028 7188 119034 7200
rect 119356 7188 119384 7287
rect 119982 7188 119988 7200
rect 119028 7160 119384 7188
rect 119943 7160 119988 7188
rect 119028 7148 119034 7160
rect 119982 7148 119988 7160
rect 120040 7148 120046 7200
rect 120368 7188 120396 7364
rect 121109 7361 121121 7395
rect 121155 7392 121167 7395
rect 124306 7392 124312 7404
rect 121155 7364 124312 7392
rect 121155 7361 121167 7364
rect 121109 7355 121167 7361
rect 124306 7352 124312 7364
rect 124364 7352 124370 7404
rect 126992 7392 127020 7500
rect 127161 7497 127173 7500
rect 127207 7497 127219 7531
rect 127161 7491 127219 7497
rect 127713 7531 127771 7537
rect 127713 7497 127725 7531
rect 127759 7528 127771 7531
rect 127802 7528 127808 7540
rect 127759 7500 127808 7528
rect 127759 7497 127771 7500
rect 127713 7491 127771 7497
rect 127802 7488 127808 7500
rect 127860 7488 127866 7540
rect 128725 7531 128783 7537
rect 128725 7497 128737 7531
rect 128771 7497 128783 7531
rect 128725 7491 128783 7497
rect 127066 7420 127072 7472
rect 127124 7460 127130 7472
rect 128740 7460 128768 7491
rect 128906 7488 128912 7540
rect 128964 7528 128970 7540
rect 129366 7528 129372 7540
rect 128964 7500 129372 7528
rect 128964 7488 128970 7500
rect 129366 7488 129372 7500
rect 129424 7488 129430 7540
rect 130194 7528 130200 7540
rect 130155 7500 130200 7528
rect 130194 7488 130200 7500
rect 130252 7488 130258 7540
rect 130838 7528 130844 7540
rect 130799 7500 130844 7528
rect 130838 7488 130844 7500
rect 130896 7488 130902 7540
rect 131206 7488 131212 7540
rect 131264 7528 131270 7540
rect 131761 7531 131819 7537
rect 131761 7528 131773 7531
rect 131264 7500 131773 7528
rect 131264 7488 131270 7500
rect 131761 7497 131773 7500
rect 131807 7497 131819 7531
rect 131761 7491 131819 7497
rect 132034 7488 132040 7540
rect 132092 7528 132098 7540
rect 133417 7531 133475 7537
rect 133417 7528 133429 7531
rect 132092 7500 133429 7528
rect 132092 7488 132098 7500
rect 133417 7497 133429 7500
rect 133463 7497 133475 7531
rect 136085 7531 136143 7537
rect 133417 7491 133475 7497
rect 134545 7500 135944 7528
rect 127124 7432 128354 7460
rect 128740 7432 129228 7460
rect 127124 7420 127130 7432
rect 127897 7395 127955 7401
rect 127897 7392 127909 7395
rect 126992 7364 127909 7392
rect 127897 7361 127909 7364
rect 127943 7361 127955 7395
rect 127897 7355 127955 7361
rect 121365 7327 121423 7333
rect 121365 7293 121377 7327
rect 121411 7324 121423 7327
rect 121638 7324 121644 7336
rect 121411 7296 121644 7324
rect 121411 7293 121423 7296
rect 121365 7287 121423 7293
rect 121638 7284 121644 7296
rect 121696 7324 121702 7336
rect 123205 7327 123263 7333
rect 121696 7296 122144 7324
rect 121696 7284 121702 7296
rect 121730 7216 121736 7268
rect 121788 7256 121794 7268
rect 121825 7259 121883 7265
rect 121825 7256 121837 7259
rect 121788 7228 121837 7256
rect 121788 7216 121794 7228
rect 121825 7225 121837 7228
rect 121871 7225 121883 7259
rect 121825 7219 121883 7225
rect 122006 7188 122012 7200
rect 120368 7160 122012 7188
rect 122006 7148 122012 7160
rect 122064 7148 122070 7200
rect 122116 7188 122144 7296
rect 123205 7293 123217 7327
rect 123251 7324 123263 7327
rect 123294 7324 123300 7336
rect 123251 7296 123300 7324
rect 123251 7293 123263 7296
rect 123205 7287 123263 7293
rect 123294 7284 123300 7296
rect 123352 7284 123358 7336
rect 123662 7284 123668 7336
rect 123720 7324 123726 7336
rect 125410 7324 125416 7336
rect 123720 7296 125416 7324
rect 123720 7284 123726 7296
rect 125410 7284 125416 7296
rect 125468 7284 125474 7336
rect 125597 7327 125655 7333
rect 125597 7293 125609 7327
rect 125643 7324 125655 7327
rect 126422 7324 126428 7336
rect 125643 7296 126428 7324
rect 125643 7293 125655 7296
rect 125597 7287 125655 7293
rect 126422 7284 126428 7296
rect 126480 7284 126486 7336
rect 126606 7324 126612 7336
rect 126567 7296 126612 7324
rect 126606 7284 126612 7296
rect 126664 7284 126670 7336
rect 127250 7284 127256 7336
rect 127308 7324 127314 7336
rect 127802 7324 127808 7336
rect 127308 7296 127808 7324
rect 127308 7284 127314 7296
rect 127802 7284 127808 7296
rect 127860 7324 127866 7336
rect 128081 7327 128139 7333
rect 128081 7324 128093 7327
rect 127860 7296 128093 7324
rect 127860 7284 127866 7296
rect 128081 7293 128093 7296
rect 128127 7293 128139 7327
rect 128326 7324 128354 7432
rect 128541 7395 128599 7401
rect 128541 7361 128553 7395
rect 128587 7392 128599 7395
rect 128906 7392 128912 7404
rect 128587 7364 128912 7392
rect 128587 7361 128599 7364
rect 128541 7355 128599 7361
rect 128906 7352 128912 7364
rect 128964 7352 128970 7404
rect 129200 7392 129228 7432
rect 129274 7420 129280 7472
rect 129332 7460 129338 7472
rect 130856 7460 130884 7488
rect 129332 7432 130884 7460
rect 129332 7420 129338 7432
rect 131942 7420 131948 7472
rect 132000 7460 132006 7472
rect 134545 7469 134573 7500
rect 132865 7463 132923 7469
rect 132865 7460 132877 7463
rect 132000 7432 132877 7460
rect 132000 7420 132006 7432
rect 132865 7429 132877 7432
rect 132911 7460 132923 7463
rect 134530 7463 134588 7469
rect 134530 7460 134542 7463
rect 132911 7432 134542 7460
rect 132911 7429 132923 7432
rect 132865 7423 132923 7429
rect 134530 7429 134542 7432
rect 134576 7429 134588 7463
rect 135916 7460 135944 7500
rect 136085 7497 136097 7531
rect 136131 7528 136143 7531
rect 137554 7528 137560 7540
rect 136131 7500 137560 7528
rect 136131 7497 136143 7500
rect 136085 7491 136143 7497
rect 137554 7488 137560 7500
rect 137612 7488 137618 7540
rect 139210 7488 139216 7540
rect 139268 7528 139274 7540
rect 141786 7528 141792 7540
rect 139268 7500 141792 7528
rect 139268 7488 139274 7500
rect 141786 7488 141792 7500
rect 141844 7488 141850 7540
rect 141881 7531 141939 7537
rect 141881 7497 141893 7531
rect 141927 7528 141939 7531
rect 141970 7528 141976 7540
rect 141927 7500 141976 7528
rect 141927 7497 141939 7500
rect 141881 7491 141939 7497
rect 141970 7488 141976 7500
rect 142028 7488 142034 7540
rect 142430 7488 142436 7540
rect 142488 7528 142494 7540
rect 146202 7528 146208 7540
rect 142488 7500 146208 7528
rect 142488 7488 142494 7500
rect 146202 7488 146208 7500
rect 146260 7488 146266 7540
rect 146956 7500 148272 7528
rect 137278 7460 137284 7472
rect 134530 7423 134588 7429
rect 134628 7432 135484 7460
rect 135916 7432 137284 7460
rect 129826 7392 129832 7404
rect 129200 7364 129832 7392
rect 129826 7352 129832 7364
rect 129884 7352 129890 7404
rect 130381 7395 130439 7401
rect 130381 7361 130393 7395
rect 130427 7392 130439 7395
rect 130838 7392 130844 7404
rect 130427 7364 130844 7392
rect 130427 7361 130439 7364
rect 130381 7355 130439 7361
rect 130838 7352 130844 7364
rect 130896 7352 130902 7404
rect 134628 7392 134656 7432
rect 134794 7392 134800 7404
rect 130948 7364 134656 7392
rect 134755 7364 134800 7392
rect 129550 7324 129556 7336
rect 128326 7296 129556 7324
rect 128081 7287 128139 7293
rect 129550 7284 129556 7296
rect 129608 7324 129614 7336
rect 130948 7324 130976 7364
rect 134794 7352 134800 7364
rect 134852 7352 134858 7404
rect 135346 7392 135352 7404
rect 135307 7364 135352 7392
rect 135346 7352 135352 7364
rect 135404 7352 135410 7404
rect 135456 7392 135484 7432
rect 137278 7420 137284 7432
rect 137336 7420 137342 7472
rect 138308 7432 141096 7460
rect 138014 7392 138020 7404
rect 135456 7364 138020 7392
rect 138014 7352 138020 7364
rect 138072 7352 138078 7404
rect 129608 7296 130976 7324
rect 129608 7284 129614 7296
rect 131298 7284 131304 7336
rect 131356 7324 131362 7336
rect 132494 7324 132500 7336
rect 131356 7296 132500 7324
rect 131356 7284 131362 7296
rect 132494 7284 132500 7296
rect 132552 7284 132558 7336
rect 137741 7327 137799 7333
rect 137741 7324 137753 7327
rect 135548 7296 137753 7324
rect 123757 7259 123815 7265
rect 123757 7225 123769 7259
rect 123803 7256 123815 7259
rect 133782 7256 133788 7268
rect 123803 7228 133788 7256
rect 123803 7225 123815 7228
rect 123757 7219 123815 7225
rect 122466 7188 122472 7200
rect 122116 7160 122472 7188
rect 122466 7148 122472 7160
rect 122524 7188 122530 7200
rect 123772 7188 123800 7219
rect 133782 7216 133788 7228
rect 133840 7216 133846 7268
rect 135548 7256 135576 7296
rect 137741 7293 137753 7296
rect 137787 7324 137799 7327
rect 138308 7324 138336 7432
rect 138385 7395 138443 7401
rect 138385 7361 138397 7395
rect 138431 7392 138443 7395
rect 138431 7364 139164 7392
rect 138431 7361 138443 7364
rect 138385 7355 138443 7361
rect 137787 7296 138336 7324
rect 138569 7327 138627 7333
rect 137787 7293 137799 7296
rect 137741 7287 137799 7293
rect 138569 7293 138581 7327
rect 138615 7324 138627 7327
rect 139029 7327 139087 7333
rect 139029 7324 139041 7327
rect 138615 7296 139041 7324
rect 138615 7293 138627 7296
rect 138569 7287 138627 7293
rect 139029 7293 139041 7296
rect 139075 7293 139087 7327
rect 139136 7324 139164 7364
rect 139210 7352 139216 7404
rect 139268 7392 139274 7404
rect 140866 7392 140872 7404
rect 139268 7364 139313 7392
rect 140827 7364 140872 7392
rect 139268 7352 139274 7364
rect 140866 7352 140872 7364
rect 140924 7352 140930 7404
rect 141068 7401 141096 7432
rect 141053 7395 141111 7401
rect 141053 7361 141065 7395
rect 141099 7392 141111 7395
rect 142448 7392 142476 7488
rect 146956 7472 146984 7500
rect 143994 7469 144000 7472
rect 143988 7423 144000 7469
rect 144052 7460 144058 7472
rect 145282 7460 145288 7472
rect 144052 7432 144088 7460
rect 144196 7432 145288 7460
rect 143994 7420 144000 7423
rect 144052 7420 144058 7432
rect 141099 7364 142476 7392
rect 143005 7395 143063 7401
rect 141099 7361 141111 7364
rect 141053 7355 141111 7361
rect 143005 7361 143017 7395
rect 143051 7392 143063 7395
rect 144196 7392 144224 7432
rect 145282 7420 145288 7432
rect 145340 7420 145346 7472
rect 146938 7460 146944 7472
rect 146312 7432 146944 7460
rect 143051 7390 143948 7392
rect 144012 7390 144224 7392
rect 143051 7364 144224 7390
rect 143051 7361 143063 7364
rect 143920 7362 144040 7364
rect 143005 7355 143063 7361
rect 144362 7352 144368 7404
rect 144420 7392 144426 7404
rect 146312 7392 146340 7432
rect 146938 7420 146944 7432
rect 146996 7420 147002 7472
rect 147340 7463 147398 7469
rect 147340 7429 147352 7463
rect 147386 7460 147398 7463
rect 148134 7460 148140 7472
rect 147386 7432 148140 7460
rect 147386 7429 147398 7432
rect 147340 7423 147398 7429
rect 148134 7420 148140 7432
rect 148192 7420 148198 7472
rect 148244 7460 148272 7500
rect 148318 7488 148324 7540
rect 148376 7528 148382 7540
rect 150434 7528 150440 7540
rect 148376 7500 150440 7528
rect 148376 7488 148382 7500
rect 150434 7488 150440 7500
rect 150492 7488 150498 7540
rect 150802 7528 150808 7540
rect 150763 7500 150808 7528
rect 150802 7488 150808 7500
rect 150860 7488 150866 7540
rect 151078 7488 151084 7540
rect 151136 7528 151142 7540
rect 154574 7528 154580 7540
rect 151136 7500 154580 7528
rect 151136 7488 151142 7500
rect 154574 7488 154580 7500
rect 154632 7488 154638 7540
rect 155313 7531 155371 7537
rect 155313 7497 155325 7531
rect 155359 7528 155371 7531
rect 155586 7528 155592 7540
rect 155359 7500 155592 7528
rect 155359 7497 155371 7500
rect 155313 7491 155371 7497
rect 155586 7488 155592 7500
rect 155644 7488 155650 7540
rect 155862 7488 155868 7540
rect 155920 7528 155926 7540
rect 156322 7528 156328 7540
rect 155920 7500 156328 7528
rect 155920 7488 155926 7500
rect 156322 7488 156328 7500
rect 156380 7488 156386 7540
rect 157610 7528 157616 7540
rect 157571 7500 157616 7528
rect 157610 7488 157616 7500
rect 157668 7488 157674 7540
rect 148496 7463 148554 7469
rect 148244 7432 148456 7460
rect 144420 7364 146340 7392
rect 144420 7352 144426 7364
rect 146386 7352 146392 7404
rect 146444 7392 146450 7404
rect 147585 7395 147643 7401
rect 147585 7392 147597 7395
rect 146444 7364 147597 7392
rect 146444 7352 146450 7364
rect 147333 7362 147383 7364
rect 147585 7361 147597 7364
rect 147631 7392 147643 7395
rect 148229 7395 148287 7401
rect 148229 7392 148241 7395
rect 147631 7364 148241 7392
rect 147631 7361 147643 7364
rect 147585 7355 147643 7361
rect 148229 7361 148241 7364
rect 148275 7361 148287 7395
rect 148428 7392 148456 7432
rect 148496 7429 148508 7463
rect 148542 7460 148554 7463
rect 148594 7460 148600 7472
rect 148542 7432 148600 7460
rect 148542 7429 148554 7432
rect 148496 7423 148554 7429
rect 148594 7420 148600 7432
rect 148652 7420 148658 7472
rect 149330 7460 149336 7472
rect 148888 7432 149336 7460
rect 148888 7392 148916 7432
rect 149330 7420 149336 7432
rect 149388 7420 149394 7472
rect 149514 7420 149520 7472
rect 149572 7460 149578 7472
rect 151918 7463 151976 7469
rect 151918 7460 151930 7463
rect 149572 7432 151930 7460
rect 149572 7420 149578 7432
rect 151918 7429 151930 7432
rect 151964 7429 151976 7463
rect 155678 7460 155684 7472
rect 151918 7423 151976 7429
rect 152016 7432 155684 7460
rect 148428 7364 148916 7392
rect 148229 7355 148287 7361
rect 148962 7352 148968 7404
rect 149020 7392 149026 7404
rect 150069 7395 150127 7401
rect 150069 7392 150081 7395
rect 149020 7364 150081 7392
rect 149020 7352 149026 7364
rect 150069 7361 150081 7364
rect 150115 7361 150127 7395
rect 152016 7392 152044 7432
rect 155678 7420 155684 7432
rect 155736 7420 155742 7472
rect 155770 7420 155776 7472
rect 155828 7460 155834 7472
rect 158257 7463 158315 7469
rect 158257 7460 158269 7463
rect 155828 7432 158269 7460
rect 155828 7420 155834 7432
rect 158257 7429 158269 7432
rect 158303 7429 158315 7463
rect 158257 7423 158315 7429
rect 150069 7355 150127 7361
rect 151208 7364 152044 7392
rect 153473 7395 153531 7401
rect 143258 7324 143264 7336
rect 139136 7296 142292 7324
rect 143219 7296 143264 7324
rect 139029 7287 139087 7293
rect 134812 7228 135576 7256
rect 122524 7160 123800 7188
rect 122524 7148 122530 7160
rect 124214 7148 124220 7200
rect 124272 7188 124278 7200
rect 124401 7191 124459 7197
rect 124401 7188 124413 7191
rect 124272 7160 124413 7188
rect 124272 7148 124278 7160
rect 124401 7157 124413 7160
rect 124447 7157 124459 7191
rect 126146 7188 126152 7200
rect 126107 7160 126152 7188
rect 124401 7151 124459 7157
rect 126146 7148 126152 7160
rect 126204 7148 126210 7200
rect 126330 7148 126336 7200
rect 126388 7188 126394 7200
rect 132034 7188 132040 7200
rect 126388 7160 132040 7188
rect 126388 7148 126394 7160
rect 132034 7148 132040 7160
rect 132092 7188 132098 7200
rect 132313 7191 132371 7197
rect 132313 7188 132325 7191
rect 132092 7160 132325 7188
rect 132092 7148 132098 7160
rect 132313 7157 132325 7160
rect 132359 7157 132371 7191
rect 132313 7151 132371 7157
rect 132494 7148 132500 7200
rect 132552 7188 132558 7200
rect 134812 7188 134840 7228
rect 136818 7216 136824 7268
rect 136876 7256 136882 7268
rect 138201 7259 138259 7265
rect 138201 7256 138213 7259
rect 136876 7228 138213 7256
rect 136876 7216 136882 7228
rect 138201 7225 138213 7228
rect 138247 7225 138259 7259
rect 138201 7219 138259 7225
rect 132552 7160 134840 7188
rect 135533 7191 135591 7197
rect 132552 7148 132558 7160
rect 135533 7157 135545 7191
rect 135579 7188 135591 7191
rect 135622 7188 135628 7200
rect 135579 7160 135628 7188
rect 135579 7157 135591 7160
rect 135533 7151 135591 7157
rect 135622 7148 135628 7160
rect 135680 7148 135686 7200
rect 136634 7188 136640 7200
rect 136595 7160 136640 7188
rect 136634 7148 136640 7160
rect 136692 7188 136698 7200
rect 137097 7191 137155 7197
rect 137097 7188 137109 7191
rect 136692 7160 137109 7188
rect 136692 7148 136698 7160
rect 137097 7157 137109 7160
rect 137143 7157 137155 7191
rect 137097 7151 137155 7157
rect 138474 7148 138480 7200
rect 138532 7188 138538 7200
rect 138934 7188 138940 7200
rect 138532 7160 138940 7188
rect 138532 7148 138538 7160
rect 138934 7148 138940 7160
rect 138992 7148 138998 7200
rect 139044 7188 139072 7287
rect 139397 7259 139455 7265
rect 139397 7225 139409 7259
rect 139443 7256 139455 7259
rect 140498 7256 140504 7268
rect 139443 7228 140504 7256
rect 139443 7225 139455 7228
rect 139397 7219 139455 7225
rect 140498 7216 140504 7228
rect 140556 7216 140562 7268
rect 139486 7188 139492 7200
rect 139044 7160 139492 7188
rect 139486 7148 139492 7160
rect 139544 7188 139550 7200
rect 139949 7191 140007 7197
rect 139949 7188 139961 7191
rect 139544 7160 139961 7188
rect 139544 7148 139550 7160
rect 139949 7157 139961 7160
rect 139995 7188 140007 7191
rect 140038 7188 140044 7200
rect 139995 7160 140044 7188
rect 139995 7157 140007 7160
rect 139949 7151 140007 7157
rect 140038 7148 140044 7160
rect 140096 7148 140102 7200
rect 140130 7148 140136 7200
rect 140188 7188 140194 7200
rect 140685 7191 140743 7197
rect 140685 7188 140697 7191
rect 140188 7160 140697 7188
rect 140188 7148 140194 7160
rect 140685 7157 140697 7160
rect 140731 7157 140743 7191
rect 142264 7188 142292 7296
rect 143258 7284 143264 7296
rect 143316 7284 143322 7336
rect 143442 7284 143448 7336
rect 143500 7324 143506 7336
rect 143721 7327 143779 7333
rect 143721 7324 143733 7327
rect 143500 7296 143733 7324
rect 143500 7284 143506 7296
rect 143721 7293 143733 7296
rect 143767 7293 143779 7327
rect 143721 7287 143779 7293
rect 145006 7284 145012 7336
rect 145064 7324 145070 7336
rect 146570 7324 146576 7336
rect 145064 7296 146576 7324
rect 145064 7284 145070 7296
rect 146570 7284 146576 7296
rect 146628 7284 146634 7336
rect 149238 7284 149244 7336
rect 149296 7324 149302 7336
rect 151208 7324 151236 7364
rect 153473 7361 153485 7395
rect 153519 7392 153531 7395
rect 153654 7392 153660 7404
rect 153519 7364 153660 7392
rect 153519 7361 153531 7364
rect 153473 7355 153531 7361
rect 153654 7352 153660 7364
rect 153712 7352 153718 7404
rect 154298 7392 154304 7404
rect 154259 7364 154304 7392
rect 154298 7352 154304 7364
rect 154356 7352 154362 7404
rect 155129 7395 155187 7401
rect 154592 7364 155080 7392
rect 152182 7324 152188 7336
rect 149296 7296 151236 7324
rect 152143 7296 152188 7324
rect 149296 7284 149302 7296
rect 152182 7284 152188 7296
rect 152240 7284 152246 7336
rect 153197 7327 153255 7333
rect 153197 7293 153209 7327
rect 153243 7324 153255 7327
rect 153286 7324 153292 7336
rect 153243 7296 153292 7324
rect 153243 7293 153255 7296
rect 153197 7287 153255 7293
rect 153286 7284 153292 7296
rect 153344 7284 153350 7336
rect 153562 7284 153568 7336
rect 153620 7324 153626 7336
rect 153930 7324 153936 7336
rect 153620 7296 153936 7324
rect 153620 7284 153626 7296
rect 153930 7284 153936 7296
rect 153988 7324 153994 7336
rect 154117 7327 154175 7333
rect 154117 7324 154129 7327
rect 153988 7296 154129 7324
rect 153988 7284 153994 7296
rect 154117 7293 154129 7296
rect 154163 7293 154175 7327
rect 154592 7324 154620 7364
rect 154117 7287 154175 7293
rect 154224 7296 154620 7324
rect 145101 7259 145159 7265
rect 145101 7225 145113 7259
rect 145147 7256 145159 7259
rect 145374 7256 145380 7268
rect 145147 7228 145380 7256
rect 145147 7225 145159 7228
rect 145101 7219 145159 7225
rect 145374 7216 145380 7228
rect 145432 7216 145438 7268
rect 145926 7216 145932 7268
rect 145984 7256 145990 7268
rect 145984 7228 146708 7256
rect 145984 7216 145990 7228
rect 146018 7188 146024 7200
rect 142264 7160 146024 7188
rect 140685 7151 140743 7157
rect 146018 7148 146024 7160
rect 146076 7148 146082 7200
rect 146110 7148 146116 7200
rect 146168 7188 146174 7200
rect 146205 7191 146263 7197
rect 146205 7188 146217 7191
rect 146168 7160 146217 7188
rect 146168 7148 146174 7160
rect 146205 7157 146217 7160
rect 146251 7157 146263 7191
rect 146680 7188 146708 7228
rect 147858 7216 147864 7268
rect 147916 7256 147922 7268
rect 147916 7228 148272 7256
rect 147916 7216 147922 7228
rect 148134 7188 148140 7200
rect 146680 7160 148140 7188
rect 146205 7151 146263 7157
rect 148134 7148 148140 7160
rect 148192 7148 148198 7200
rect 148244 7188 148272 7228
rect 149535 7228 151308 7256
rect 149535 7188 149563 7228
rect 148244 7160 149563 7188
rect 149609 7191 149667 7197
rect 149609 7157 149621 7191
rect 149655 7188 149667 7191
rect 149790 7188 149796 7200
rect 149655 7160 149796 7188
rect 149655 7157 149667 7160
rect 149609 7151 149667 7157
rect 149790 7148 149796 7160
rect 149848 7148 149854 7200
rect 151280 7188 151308 7228
rect 153470 7216 153476 7268
rect 153528 7256 153534 7268
rect 154224 7256 154252 7296
rect 154758 7284 154764 7336
rect 154816 7324 154822 7336
rect 154945 7327 155003 7333
rect 154945 7324 154957 7327
rect 154816 7296 154957 7324
rect 154816 7284 154822 7296
rect 154945 7293 154957 7296
rect 154991 7293 155003 7327
rect 155052 7324 155080 7364
rect 155129 7361 155141 7395
rect 155175 7392 155187 7395
rect 155586 7392 155592 7404
rect 155175 7364 155592 7392
rect 155175 7361 155187 7364
rect 155129 7355 155187 7361
rect 155586 7352 155592 7364
rect 155644 7352 155650 7404
rect 156046 7352 156052 7404
rect 156104 7392 156110 7404
rect 156141 7395 156199 7401
rect 156141 7392 156153 7395
rect 156104 7364 156153 7392
rect 156104 7352 156110 7364
rect 156141 7361 156153 7364
rect 156187 7361 156199 7395
rect 156966 7392 156972 7404
rect 156927 7364 156972 7392
rect 156141 7355 156199 7361
rect 156966 7352 156972 7364
rect 157024 7352 157030 7404
rect 157794 7392 157800 7404
rect 157755 7364 157800 7392
rect 157794 7352 157800 7364
rect 157852 7352 157858 7404
rect 155957 7327 156015 7333
rect 155957 7324 155969 7327
rect 155052 7296 155969 7324
rect 154945 7287 155003 7293
rect 155957 7293 155969 7296
rect 156003 7324 156015 7327
rect 156230 7324 156236 7336
rect 156003 7296 156236 7324
rect 156003 7293 156015 7296
rect 155957 7287 156015 7293
rect 156230 7284 156236 7296
rect 156288 7324 156294 7336
rect 156690 7324 156696 7336
rect 156288 7296 156696 7324
rect 156288 7284 156294 7296
rect 156690 7284 156696 7296
rect 156748 7324 156754 7336
rect 156785 7327 156843 7333
rect 156785 7324 156797 7327
rect 156748 7296 156797 7324
rect 156748 7284 156754 7296
rect 156785 7293 156797 7296
rect 156831 7293 156843 7327
rect 156785 7287 156843 7293
rect 155678 7256 155684 7268
rect 153528 7228 154252 7256
rect 154316 7228 155684 7256
rect 153528 7216 153534 7228
rect 154316 7188 154344 7228
rect 155678 7216 155684 7228
rect 155736 7216 155742 7268
rect 157153 7259 157211 7265
rect 157153 7225 157165 7259
rect 157199 7256 157211 7259
rect 157518 7256 157524 7268
rect 157199 7228 157524 7256
rect 157199 7225 157211 7228
rect 157153 7219 157211 7225
rect 157518 7216 157524 7228
rect 157576 7216 157582 7268
rect 151280 7160 154344 7188
rect 154390 7148 154396 7200
rect 154448 7188 154454 7200
rect 154485 7191 154543 7197
rect 154485 7188 154497 7191
rect 154448 7160 154497 7188
rect 154448 7148 154454 7160
rect 154485 7157 154497 7160
rect 154531 7157 154543 7191
rect 154485 7151 154543 7157
rect 154758 7148 154764 7200
rect 154816 7188 154822 7200
rect 155770 7188 155776 7200
rect 154816 7160 155776 7188
rect 154816 7148 154822 7160
rect 155770 7148 155776 7160
rect 155828 7148 155834 7200
rect 156325 7191 156383 7197
rect 156325 7157 156337 7191
rect 156371 7188 156383 7191
rect 156966 7188 156972 7200
rect 156371 7160 156972 7188
rect 156371 7157 156383 7160
rect 156325 7151 156383 7157
rect 156966 7148 156972 7160
rect 157024 7148 157030 7200
rect 1104 7098 158884 7120
rect 1104 7046 20672 7098
rect 20724 7046 20736 7098
rect 20788 7046 20800 7098
rect 20852 7046 20864 7098
rect 20916 7046 20928 7098
rect 20980 7046 60117 7098
rect 60169 7046 60181 7098
rect 60233 7046 60245 7098
rect 60297 7046 60309 7098
rect 60361 7046 60373 7098
rect 60425 7046 99562 7098
rect 99614 7046 99626 7098
rect 99678 7046 99690 7098
rect 99742 7046 99754 7098
rect 99806 7046 99818 7098
rect 99870 7046 139007 7098
rect 139059 7046 139071 7098
rect 139123 7046 139135 7098
rect 139187 7046 139199 7098
rect 139251 7046 139263 7098
rect 139315 7046 158884 7098
rect 1104 7024 158884 7046
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13446 6984 13452 6996
rect 13035 6956 13452 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 14826 6944 14832 6996
rect 14884 6984 14890 6996
rect 20254 6984 20260 6996
rect 14884 6956 18460 6984
rect 14884 6944 14890 6956
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 18325 6919 18383 6925
rect 18325 6916 18337 6919
rect 17920 6888 18337 6916
rect 17920 6876 17926 6888
rect 18325 6885 18337 6888
rect 18371 6885 18383 6919
rect 18325 6879 18383 6885
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 15160 6820 16221 6848
rect 15160 6808 15166 6820
rect 16209 6817 16221 6820
rect 16255 6817 16267 6851
rect 18432 6848 18460 6956
rect 19904 6956 20260 6984
rect 19904 6860 19932 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 30374 6944 30380 6996
rect 30432 6984 30438 6996
rect 34882 6984 34888 6996
rect 30432 6956 34888 6984
rect 30432 6944 30438 6956
rect 34882 6944 34888 6956
rect 34940 6944 34946 6996
rect 37642 6984 37648 6996
rect 37603 6956 37648 6984
rect 37642 6944 37648 6956
rect 37700 6984 37706 6996
rect 40218 6984 40224 6996
rect 37700 6956 40224 6984
rect 37700 6944 37706 6956
rect 40218 6944 40224 6956
rect 40276 6944 40282 6996
rect 51629 6987 51687 6993
rect 44928 6956 45508 6984
rect 24857 6919 24915 6925
rect 24857 6885 24869 6919
rect 24903 6885 24915 6919
rect 33962 6916 33968 6928
rect 24857 6879 24915 6885
rect 33152 6888 33968 6916
rect 18693 6851 18751 6857
rect 18693 6848 18705 6851
rect 18432 6820 18705 6848
rect 16209 6811 16267 6817
rect 18693 6817 18705 6820
rect 18739 6848 18751 6851
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 18739 6820 19441 6848
rect 18739 6817 18751 6820
rect 18693 6811 18751 6817
rect 19429 6817 19441 6820
rect 19475 6848 19487 6851
rect 19886 6848 19892 6860
rect 19475 6820 19892 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 20070 6848 20076 6860
rect 20031 6820 20076 6848
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 21726 6808 21732 6860
rect 21784 6848 21790 6860
rect 24872 6848 24900 6879
rect 21784 6820 24900 6848
rect 26237 6851 26295 6857
rect 21784 6808 21790 6820
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26326 6848 26332 6860
rect 26283 6820 26332 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26326 6808 26332 6820
rect 26384 6848 26390 6860
rect 30190 6848 30196 6860
rect 26384 6820 30196 6848
rect 26384 6808 26390 6820
rect 30190 6808 30196 6820
rect 30248 6808 30254 6860
rect 32030 6808 32036 6860
rect 32088 6848 32094 6860
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 32088 6820 32781 6848
rect 32088 6808 32094 6820
rect 32769 6817 32781 6820
rect 32815 6848 32827 6851
rect 33152 6848 33180 6888
rect 33962 6876 33968 6888
rect 34020 6876 34026 6928
rect 37182 6876 37188 6928
rect 37240 6916 37246 6928
rect 37240 6888 37964 6916
rect 37240 6876 37246 6888
rect 32815 6820 33180 6848
rect 32815 6817 32827 6820
rect 32769 6811 32827 6817
rect 33226 6808 33232 6860
rect 33284 6848 33290 6860
rect 33502 6848 33508 6860
rect 33284 6820 33508 6848
rect 33284 6808 33290 6820
rect 33502 6808 33508 6820
rect 33560 6808 33566 6860
rect 33873 6851 33931 6857
rect 33873 6817 33885 6851
rect 33919 6848 33931 6851
rect 37826 6848 37832 6860
rect 33919 6820 37832 6848
rect 33919 6817 33931 6820
rect 33873 6811 33931 6817
rect 37826 6808 37832 6820
rect 37884 6808 37890 6860
rect 37936 6848 37964 6888
rect 38105 6851 38163 6857
rect 38105 6848 38117 6851
rect 37936 6820 38117 6848
rect 38105 6817 38117 6820
rect 38151 6817 38163 6851
rect 44928 6848 44956 6956
rect 38105 6811 38163 6817
rect 41386 6820 44956 6848
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 13262 6780 13268 6792
rect 11931 6752 13268 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6780 15255 6783
rect 15286 6780 15292 6792
rect 15243 6752 15292 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16482 6789 16488 6792
rect 16476 6780 16488 6789
rect 16443 6752 16488 6780
rect 16476 6743 16488 6752
rect 16482 6740 16488 6743
rect 16540 6740 16546 6792
rect 18506 6780 18512 6792
rect 18467 6752 18512 6780
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18800 6752 20484 6780
rect 13722 6712 13728 6724
rect 13635 6684 13728 6712
rect 13722 6672 13728 6684
rect 13780 6712 13786 6724
rect 13780 6684 17724 6712
rect 13780 6672 13786 6684
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4525 6647 4583 6653
rect 4525 6644 4537 6647
rect 4120 6616 4537 6644
rect 4120 6604 4126 6616
rect 4525 6613 4537 6616
rect 4571 6613 4583 6647
rect 11698 6644 11704 6656
rect 11659 6616 11704 6644
rect 4525 6607 4583 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15381 6647 15439 6653
rect 15381 6613 15393 6647
rect 15427 6644 15439 6647
rect 16850 6644 16856 6656
rect 15427 6616 16856 6644
rect 15427 6613 15439 6616
rect 15381 6607 15439 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17276 6616 17601 6644
rect 17276 6604 17282 6616
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 17696 6644 17724 6684
rect 18800 6644 18828 6752
rect 19886 6672 19892 6724
rect 19944 6712 19950 6724
rect 20318 6715 20376 6721
rect 20318 6712 20330 6715
rect 19944 6684 20330 6712
rect 19944 6672 19950 6684
rect 20318 6681 20330 6684
rect 20364 6681 20376 6715
rect 20456 6712 20484 6752
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 22097 6783 22155 6789
rect 22097 6780 22109 6783
rect 21232 6752 22109 6780
rect 21232 6740 21238 6752
rect 22097 6749 22109 6752
rect 22143 6749 22155 6783
rect 27062 6780 27068 6792
rect 22097 6743 22155 6749
rect 22204 6752 26096 6780
rect 27023 6752 27068 6780
rect 22204 6712 22232 6752
rect 23566 6712 23572 6724
rect 20456 6684 22232 6712
rect 22296 6684 23572 6712
rect 20318 6675 20376 6681
rect 17696 6616 18828 6644
rect 17589 6607 17647 6613
rect 18874 6604 18880 6656
rect 18932 6644 18938 6656
rect 21450 6644 21456 6656
rect 18932 6616 21456 6644
rect 18932 6604 18938 6616
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 22296 6653 22324 6684
rect 23566 6672 23572 6684
rect 23624 6672 23630 6724
rect 25970 6715 26028 6721
rect 25970 6712 25982 6715
rect 23952 6684 25982 6712
rect 22281 6647 22339 6653
rect 22281 6613 22293 6647
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 22741 6647 22799 6653
rect 22741 6644 22753 6647
rect 22612 6616 22753 6644
rect 22612 6604 22618 6616
rect 22741 6613 22753 6616
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 23842 6604 23848 6656
rect 23900 6644 23906 6656
rect 23952 6653 23980 6684
rect 25970 6681 25982 6684
rect 26016 6681 26028 6715
rect 26068 6712 26096 6752
rect 27062 6740 27068 6752
rect 27120 6740 27126 6792
rect 33689 6783 33747 6789
rect 33689 6749 33701 6783
rect 33735 6780 33747 6783
rect 33962 6780 33968 6792
rect 33735 6752 33968 6780
rect 33735 6749 33747 6752
rect 33689 6743 33747 6749
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 36538 6780 36544 6792
rect 36499 6752 36544 6780
rect 36538 6740 36544 6752
rect 36596 6740 36602 6792
rect 36998 6780 37004 6792
rect 36959 6752 37004 6780
rect 36998 6740 37004 6752
rect 37056 6740 37062 6792
rect 41386 6780 41414 6820
rect 45002 6808 45008 6860
rect 45060 6848 45066 6860
rect 45480 6848 45508 6956
rect 51629 6953 51641 6987
rect 51675 6984 51687 6987
rect 52362 6984 52368 6996
rect 51675 6956 52368 6984
rect 51675 6953 51687 6956
rect 51629 6947 51687 6953
rect 52362 6944 52368 6956
rect 52420 6944 52426 6996
rect 54202 6944 54208 6996
rect 54260 6984 54266 6996
rect 54481 6987 54539 6993
rect 54481 6984 54493 6987
rect 54260 6956 54493 6984
rect 54260 6944 54266 6956
rect 54481 6953 54493 6956
rect 54527 6953 54539 6987
rect 63678 6984 63684 6996
rect 63639 6956 63684 6984
rect 54481 6947 54539 6953
rect 63678 6944 63684 6956
rect 63736 6944 63742 6996
rect 119982 6984 119988 6996
rect 63788 6956 119988 6984
rect 50522 6876 50528 6928
rect 50580 6916 50586 6928
rect 50709 6919 50767 6925
rect 50709 6916 50721 6919
rect 50580 6888 50721 6916
rect 50580 6876 50586 6888
rect 50709 6885 50721 6888
rect 50755 6916 50767 6919
rect 55766 6916 55772 6928
rect 50755 6888 55772 6916
rect 50755 6885 50767 6888
rect 50709 6879 50767 6885
rect 55766 6876 55772 6888
rect 55824 6876 55830 6928
rect 61654 6876 61660 6928
rect 61712 6916 61718 6928
rect 63788 6916 63816 6956
rect 119982 6944 119988 6956
rect 120040 6944 120046 6996
rect 120626 6984 120632 6996
rect 120276 6956 120632 6984
rect 61712 6888 63816 6916
rect 61712 6876 61718 6888
rect 82998 6876 83004 6928
rect 83056 6916 83062 6928
rect 86770 6916 86776 6928
rect 83056 6888 86776 6916
rect 83056 6876 83062 6888
rect 86770 6876 86776 6888
rect 86828 6876 86834 6928
rect 108942 6876 108948 6928
rect 109000 6916 109006 6928
rect 110598 6916 110604 6928
rect 109000 6888 109172 6916
rect 110559 6888 110604 6916
rect 109000 6876 109006 6888
rect 50430 6848 50436 6860
rect 45060 6820 45324 6848
rect 45480 6820 50436 6848
rect 45060 6808 45066 6820
rect 43530 6780 43536 6792
rect 37108 6752 41414 6780
rect 43491 6752 43536 6780
rect 30558 6712 30564 6724
rect 26068 6684 30564 6712
rect 25970 6675 26028 6681
rect 30558 6672 30564 6684
rect 30616 6672 30622 6724
rect 30650 6672 30656 6724
rect 30708 6712 30714 6724
rect 37108 6712 37136 6752
rect 43530 6740 43536 6752
rect 43588 6740 43594 6792
rect 43717 6783 43775 6789
rect 43717 6749 43729 6783
rect 43763 6780 43775 6783
rect 44174 6780 44180 6792
rect 43763 6752 44180 6780
rect 43763 6749 43775 6752
rect 43717 6743 43775 6749
rect 44174 6740 44180 6752
rect 44232 6780 44238 6792
rect 45094 6780 45100 6792
rect 44232 6752 45100 6780
rect 44232 6740 44238 6752
rect 45094 6740 45100 6752
rect 45152 6740 45158 6792
rect 45296 6780 45324 6820
rect 50430 6808 50436 6820
rect 50488 6808 50494 6860
rect 52086 6848 52092 6860
rect 52047 6820 52092 6848
rect 52086 6808 52092 6820
rect 52144 6808 52150 6860
rect 56318 6848 56324 6860
rect 53852 6820 56324 6848
rect 45296 6752 45600 6780
rect 38378 6721 38384 6724
rect 38372 6712 38384 6721
rect 30708 6684 37136 6712
rect 38339 6684 38384 6712
rect 30708 6672 30714 6684
rect 38372 6675 38384 6684
rect 38378 6672 38384 6675
rect 38436 6672 38442 6724
rect 43901 6715 43959 6721
rect 43901 6681 43913 6715
rect 43947 6712 43959 6715
rect 45462 6712 45468 6724
rect 43947 6684 45468 6712
rect 43947 6681 43959 6684
rect 43901 6675 43959 6681
rect 45462 6672 45468 6684
rect 45520 6672 45526 6724
rect 45572 6712 45600 6752
rect 46198 6740 46204 6792
rect 46256 6780 46262 6792
rect 52270 6780 52276 6792
rect 46256 6752 52276 6780
rect 46256 6740 46262 6752
rect 52270 6740 52276 6752
rect 52328 6740 52334 6792
rect 53852 6789 53880 6820
rect 56318 6808 56324 6820
rect 56376 6808 56382 6860
rect 58986 6808 58992 6860
rect 59044 6848 59050 6860
rect 68465 6851 68523 6857
rect 59044 6820 59676 6848
rect 59044 6808 59050 6820
rect 53837 6783 53895 6789
rect 53837 6749 53849 6783
rect 53883 6749 53895 6783
rect 53837 6743 53895 6749
rect 54021 6783 54079 6789
rect 54021 6749 54033 6783
rect 54067 6780 54079 6783
rect 54294 6780 54300 6792
rect 54067 6752 54300 6780
rect 54067 6749 54079 6752
rect 54021 6743 54079 6749
rect 54294 6740 54300 6752
rect 54352 6780 54358 6792
rect 55493 6783 55551 6789
rect 55493 6780 55505 6783
rect 54352 6752 55505 6780
rect 54352 6740 54358 6752
rect 55493 6749 55505 6752
rect 55539 6780 55551 6783
rect 57514 6780 57520 6792
rect 55539 6752 57520 6780
rect 55539 6749 55551 6752
rect 55493 6743 55551 6749
rect 57514 6740 57520 6752
rect 57572 6780 57578 6792
rect 59648 6789 59676 6820
rect 68465 6817 68477 6851
rect 68511 6848 68523 6851
rect 69106 6848 69112 6860
rect 68511 6820 69112 6848
rect 68511 6817 68523 6820
rect 68465 6811 68523 6817
rect 69106 6808 69112 6820
rect 69164 6808 69170 6860
rect 81158 6848 81164 6860
rect 80026 6820 81164 6848
rect 57609 6783 57667 6789
rect 57609 6780 57621 6783
rect 57572 6752 57621 6780
rect 57572 6740 57578 6752
rect 57609 6749 57621 6752
rect 57655 6749 57667 6783
rect 57609 6743 57667 6749
rect 59449 6783 59507 6789
rect 59449 6749 59461 6783
rect 59495 6749 59507 6783
rect 59449 6743 59507 6749
rect 59633 6783 59691 6789
rect 59633 6749 59645 6783
rect 59679 6780 59691 6783
rect 59722 6780 59728 6792
rect 59679 6752 59728 6780
rect 59679 6749 59691 6752
rect 59633 6743 59691 6749
rect 46566 6712 46572 6724
rect 45572 6684 46572 6712
rect 46566 6672 46572 6684
rect 46624 6672 46630 6724
rect 47026 6672 47032 6724
rect 47084 6712 47090 6724
rect 50706 6712 50712 6724
rect 47084 6684 50712 6712
rect 47084 6672 47090 6684
rect 50706 6672 50712 6684
rect 50764 6672 50770 6724
rect 52178 6672 52184 6724
rect 52236 6712 52242 6724
rect 52733 6715 52791 6721
rect 52733 6712 52745 6715
rect 52236 6684 52745 6712
rect 52236 6672 52242 6684
rect 52733 6681 52745 6684
rect 52779 6712 52791 6715
rect 57146 6712 57152 6724
rect 52779 6684 57152 6712
rect 52779 6681 52791 6684
rect 52733 6675 52791 6681
rect 57146 6672 57152 6684
rect 57204 6672 57210 6724
rect 59464 6712 59492 6743
rect 59722 6740 59728 6752
rect 59780 6780 59786 6792
rect 64414 6780 64420 6792
rect 59780 6752 64420 6780
rect 59780 6740 59786 6752
rect 64414 6740 64420 6752
rect 64472 6740 64478 6792
rect 64506 6740 64512 6792
rect 64564 6780 64570 6792
rect 64794 6783 64852 6789
rect 64794 6780 64806 6783
rect 64564 6752 64806 6780
rect 64564 6740 64570 6752
rect 64794 6749 64806 6752
rect 64840 6749 64852 6783
rect 64794 6743 64852 6749
rect 65061 6783 65119 6789
rect 65061 6749 65073 6783
rect 65107 6749 65119 6783
rect 66530 6780 66536 6792
rect 66491 6752 66536 6780
rect 65061 6743 65119 6749
rect 60458 6712 60464 6724
rect 59464 6684 60464 6712
rect 60458 6672 60464 6684
rect 60516 6712 60522 6724
rect 65076 6712 65104 6743
rect 66530 6740 66536 6752
rect 66588 6740 66594 6792
rect 73154 6780 73160 6792
rect 66640 6752 73160 6780
rect 66640 6724 66668 6752
rect 73154 6740 73160 6752
rect 73212 6780 73218 6792
rect 73709 6783 73767 6789
rect 73709 6780 73721 6783
rect 73212 6752 73721 6780
rect 73212 6740 73218 6752
rect 73709 6749 73721 6752
rect 73755 6780 73767 6783
rect 73798 6780 73804 6792
rect 73755 6752 73804 6780
rect 73755 6749 73767 6752
rect 73709 6743 73767 6749
rect 73798 6740 73804 6752
rect 73856 6780 73862 6792
rect 75549 6783 75607 6789
rect 75549 6780 75561 6783
rect 73856 6752 75561 6780
rect 73856 6740 73862 6752
rect 75549 6749 75561 6752
rect 75595 6780 75607 6783
rect 75914 6780 75920 6792
rect 75595 6752 75920 6780
rect 75595 6749 75607 6752
rect 75549 6743 75607 6749
rect 75914 6740 75920 6752
rect 75972 6780 75978 6792
rect 76101 6783 76159 6789
rect 76101 6780 76113 6783
rect 75972 6752 76113 6780
rect 75972 6740 75978 6752
rect 76101 6749 76113 6752
rect 76147 6780 76159 6783
rect 78861 6783 78919 6789
rect 78861 6780 78873 6783
rect 76147 6752 78873 6780
rect 76147 6749 76159 6752
rect 76101 6743 76159 6749
rect 78861 6749 78873 6752
rect 78907 6780 78919 6783
rect 79042 6780 79048 6792
rect 78907 6752 79048 6780
rect 78907 6749 78919 6752
rect 78861 6743 78919 6749
rect 79042 6740 79048 6752
rect 79100 6740 79106 6792
rect 79134 6740 79140 6792
rect 79192 6780 79198 6792
rect 80026 6780 80054 6820
rect 81158 6808 81164 6820
rect 81216 6808 81222 6860
rect 88245 6851 88303 6857
rect 88245 6817 88257 6851
rect 88291 6848 88303 6851
rect 88291 6820 92336 6848
rect 88291 6817 88303 6820
rect 88245 6811 88303 6817
rect 79192 6752 80054 6780
rect 81176 6752 82584 6780
rect 79192 6740 79198 6752
rect 65889 6715 65947 6721
rect 65889 6712 65901 6715
rect 60516 6684 65012 6712
rect 65076 6684 65901 6712
rect 60516 6672 60522 6684
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 23900 6616 23949 6644
rect 23900 6604 23906 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 26234 6644 26240 6656
rect 25648 6616 26240 6644
rect 25648 6604 25654 6616
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 26878 6644 26884 6656
rect 26839 6616 26884 6644
rect 26878 6604 26884 6616
rect 26936 6604 26942 6656
rect 36354 6644 36360 6656
rect 36315 6616 36360 6644
rect 36354 6604 36360 6616
rect 36412 6604 36418 6656
rect 36446 6604 36452 6656
rect 36504 6644 36510 6656
rect 39485 6647 39543 6653
rect 39485 6644 39497 6647
rect 36504 6616 39497 6644
rect 36504 6604 36510 6616
rect 39485 6613 39497 6616
rect 39531 6613 39543 6647
rect 39485 6607 39543 6613
rect 43530 6604 43536 6656
rect 43588 6644 43594 6656
rect 44358 6644 44364 6656
rect 43588 6616 44364 6644
rect 43588 6604 43594 6616
rect 44358 6604 44364 6616
rect 44416 6604 44422 6656
rect 53374 6604 53380 6656
rect 53432 6644 53438 6656
rect 53653 6647 53711 6653
rect 53653 6644 53665 6647
rect 53432 6616 53665 6644
rect 53432 6604 53438 6616
rect 53653 6613 53665 6616
rect 53699 6613 53711 6647
rect 53653 6607 53711 6613
rect 58618 6604 58624 6656
rect 58676 6644 58682 6656
rect 59265 6647 59323 6653
rect 59265 6644 59277 6647
rect 58676 6616 59277 6644
rect 58676 6604 58682 6616
rect 59265 6613 59277 6616
rect 59311 6613 59323 6647
rect 64984 6644 65012 6684
rect 65889 6681 65901 6684
rect 65935 6712 65947 6715
rect 66622 6712 66628 6724
rect 65935 6684 66628 6712
rect 65935 6681 65947 6684
rect 65889 6675 65947 6681
rect 66622 6672 66628 6684
rect 66680 6672 66686 6724
rect 66800 6715 66858 6721
rect 66800 6681 66812 6715
rect 66846 6712 66858 6715
rect 66846 6684 73292 6712
rect 66846 6681 66858 6684
rect 66800 6675 66858 6681
rect 66254 6644 66260 6656
rect 64984 6616 66260 6644
rect 59265 6607 59323 6613
rect 66254 6604 66260 6616
rect 66312 6604 66318 6656
rect 67910 6644 67916 6656
rect 67871 6616 67916 6644
rect 67910 6604 67916 6616
rect 67968 6604 67974 6656
rect 72326 6644 72332 6656
rect 72287 6616 72332 6644
rect 72326 6604 72332 6616
rect 72384 6604 72390 6656
rect 73264 6644 73292 6684
rect 73338 6672 73344 6724
rect 73396 6712 73402 6724
rect 73442 6715 73500 6721
rect 73442 6712 73454 6715
rect 73396 6684 73454 6712
rect 73396 6672 73402 6684
rect 73442 6681 73454 6684
rect 73488 6681 73500 6715
rect 75178 6712 75184 6724
rect 73442 6675 73500 6681
rect 73540 6684 75184 6712
rect 73540 6644 73568 6684
rect 75178 6672 75184 6684
rect 75236 6672 75242 6724
rect 75304 6715 75362 6721
rect 75304 6681 75316 6715
rect 75350 6712 75362 6715
rect 76006 6712 76012 6724
rect 75350 6684 76012 6712
rect 75350 6681 75362 6684
rect 75304 6675 75362 6681
rect 76006 6672 76012 6684
rect 76064 6672 76070 6724
rect 79060 6712 79088 6740
rect 81176 6724 81204 6752
rect 81158 6712 81164 6724
rect 79060 6684 81164 6712
rect 81158 6672 81164 6684
rect 81216 6672 81222 6724
rect 82377 6715 82435 6721
rect 82377 6681 82389 6715
rect 82423 6712 82435 6715
rect 82556 6712 82584 6752
rect 82630 6740 82636 6792
rect 82688 6780 82694 6792
rect 87785 6783 87843 6789
rect 87785 6780 87797 6783
rect 82688 6752 82733 6780
rect 85776 6752 87797 6780
rect 82688 6740 82694 6752
rect 85776 6721 85804 6752
rect 87785 6749 87797 6752
rect 87831 6780 87843 6783
rect 88334 6780 88340 6792
rect 87831 6752 88340 6780
rect 87831 6749 87843 6752
rect 87785 6743 87843 6749
rect 88334 6740 88340 6752
rect 88392 6740 88398 6792
rect 85761 6715 85819 6721
rect 85761 6712 85773 6715
rect 82423 6684 82492 6712
rect 82556 6684 85773 6712
rect 82423 6681 82435 6684
rect 82377 6675 82435 6681
rect 73264 6616 73568 6644
rect 74169 6647 74227 6653
rect 74169 6613 74181 6647
rect 74215 6644 74227 6647
rect 74626 6644 74632 6656
rect 74215 6616 74632 6644
rect 74215 6613 74227 6616
rect 74169 6607 74227 6613
rect 74626 6604 74632 6616
rect 74684 6604 74690 6656
rect 75086 6604 75092 6656
rect 75144 6644 75150 6656
rect 79318 6644 79324 6656
rect 75144 6616 79324 6644
rect 75144 6604 75150 6616
rect 79318 6604 79324 6616
rect 79376 6604 79382 6656
rect 80606 6604 80612 6656
rect 80664 6644 80670 6656
rect 81253 6647 81311 6653
rect 81253 6644 81265 6647
rect 80664 6616 81265 6644
rect 80664 6604 80670 6616
rect 81253 6613 81265 6616
rect 81299 6613 81311 6647
rect 82464 6644 82492 6684
rect 85761 6681 85773 6684
rect 85807 6681 85819 6715
rect 87540 6715 87598 6721
rect 85761 6675 85819 6681
rect 85868 6684 86540 6712
rect 83185 6647 83243 6653
rect 83185 6644 83197 6647
rect 82464 6616 83197 6644
rect 81253 6607 81311 6613
rect 83185 6613 83197 6616
rect 83231 6644 83243 6647
rect 85868 6644 85896 6684
rect 86402 6644 86408 6656
rect 83231 6616 85896 6644
rect 86363 6616 86408 6644
rect 83231 6613 83243 6616
rect 83185 6607 83243 6613
rect 86402 6604 86408 6616
rect 86460 6604 86466 6656
rect 86512 6644 86540 6684
rect 87540 6681 87552 6715
rect 87586 6712 87598 6715
rect 88444 6712 88472 6820
rect 92198 6780 92204 6792
rect 87586 6684 88472 6712
rect 89686 6752 92204 6780
rect 87586 6681 87598 6684
rect 87540 6675 87598 6681
rect 89686 6644 89714 6752
rect 92198 6740 92204 6752
rect 92256 6740 92262 6792
rect 92308 6780 92336 6820
rect 93302 6808 93308 6860
rect 93360 6848 93366 6860
rect 93857 6851 93915 6857
rect 93857 6848 93869 6851
rect 93360 6820 93869 6848
rect 93360 6808 93366 6820
rect 93857 6817 93869 6820
rect 93903 6848 93915 6851
rect 96798 6848 96804 6860
rect 93903 6820 96804 6848
rect 93903 6817 93915 6820
rect 93857 6811 93915 6817
rect 96798 6808 96804 6820
rect 96856 6808 96862 6860
rect 96890 6808 96896 6860
rect 96948 6848 96954 6860
rect 101582 6848 101588 6860
rect 96948 6820 101588 6848
rect 96948 6808 96954 6820
rect 101582 6808 101588 6820
rect 101640 6808 101646 6860
rect 103606 6808 103612 6860
rect 103664 6848 103670 6860
rect 106918 6848 106924 6860
rect 103664 6820 106924 6848
rect 103664 6808 103670 6820
rect 106918 6808 106924 6820
rect 106976 6808 106982 6860
rect 108390 6848 108396 6860
rect 108351 6820 108396 6848
rect 108390 6808 108396 6820
rect 108448 6848 108454 6860
rect 108850 6848 108856 6860
rect 108448 6820 108856 6848
rect 108448 6808 108454 6820
rect 108850 6808 108856 6820
rect 108908 6808 108914 6860
rect 109144 6848 109172 6888
rect 110598 6876 110604 6888
rect 110656 6876 110662 6928
rect 111058 6916 111064 6928
rect 111019 6888 111064 6916
rect 111058 6876 111064 6888
rect 111116 6876 111122 6928
rect 111334 6876 111340 6928
rect 111392 6916 111398 6928
rect 111392 6888 111472 6916
rect 111392 6876 111398 6888
rect 111444 6848 111472 6888
rect 111518 6876 111524 6928
rect 111576 6916 111582 6928
rect 112898 6916 112904 6928
rect 111576 6888 112904 6916
rect 111576 6876 111582 6888
rect 112898 6876 112904 6888
rect 112956 6876 112962 6928
rect 114462 6876 114468 6928
rect 114520 6916 114526 6928
rect 115385 6919 115443 6925
rect 115385 6916 115397 6919
rect 114520 6888 115397 6916
rect 114520 6876 114526 6888
rect 112809 6851 112867 6857
rect 112809 6848 112821 6851
rect 109144 6820 111380 6848
rect 111444 6820 112821 6848
rect 105446 6780 105452 6792
rect 92308 6752 105452 6780
rect 105446 6740 105452 6752
rect 105504 6740 105510 6792
rect 105722 6740 105728 6792
rect 105780 6780 105786 6792
rect 108137 6783 108195 6789
rect 105780 6752 108068 6780
rect 105780 6740 105786 6752
rect 92474 6672 92480 6724
rect 92532 6712 92538 6724
rect 93038 6715 93096 6721
rect 93038 6712 93050 6715
rect 92532 6684 93050 6712
rect 92532 6672 92538 6684
rect 93038 6681 93050 6684
rect 93084 6681 93096 6715
rect 93038 6675 93096 6681
rect 93210 6672 93216 6724
rect 93268 6712 93274 6724
rect 99374 6712 99380 6724
rect 93268 6684 99380 6712
rect 93268 6672 93274 6684
rect 99374 6672 99380 6684
rect 99432 6672 99438 6724
rect 101582 6672 101588 6724
rect 101640 6712 101646 6724
rect 107378 6712 107384 6724
rect 101640 6684 107384 6712
rect 101640 6672 101646 6684
rect 107378 6672 107384 6684
rect 107436 6672 107442 6724
rect 108040 6712 108068 6752
rect 108137 6749 108149 6783
rect 108183 6780 108195 6783
rect 110598 6780 110604 6792
rect 108183 6752 110604 6780
rect 108183 6749 108195 6752
rect 108137 6743 108195 6749
rect 110598 6740 110604 6752
rect 110656 6740 110662 6792
rect 110690 6740 110696 6792
rect 110748 6780 110754 6792
rect 111225 6785 111283 6791
rect 111225 6782 111237 6785
rect 111168 6780 111237 6782
rect 110748 6754 111237 6780
rect 110748 6752 111196 6754
rect 110748 6740 110754 6752
rect 111225 6751 111237 6754
rect 111271 6751 111283 6785
rect 111352 6780 111380 6820
rect 112809 6817 112821 6820
rect 112855 6848 112867 6851
rect 113082 6848 113088 6860
rect 112855 6820 113088 6848
rect 112855 6817 112867 6820
rect 112809 6811 112867 6817
rect 113082 6808 113088 6820
rect 113140 6808 113146 6860
rect 114554 6848 114560 6860
rect 114515 6820 114560 6848
rect 114554 6808 114560 6820
rect 114612 6808 114618 6860
rect 114940 6857 114968 6888
rect 115385 6885 115397 6888
rect 115431 6885 115443 6919
rect 115385 6879 115443 6885
rect 116670 6876 116676 6928
rect 116728 6916 116734 6928
rect 120276 6916 120304 6956
rect 120626 6944 120632 6956
rect 120684 6984 120690 6996
rect 124214 6984 124220 6996
rect 120684 6956 124220 6984
rect 120684 6944 120690 6956
rect 124214 6944 124220 6956
rect 124272 6944 124278 6996
rect 125152 6956 125732 6984
rect 116728 6888 120304 6916
rect 116728 6876 116734 6888
rect 122006 6876 122012 6928
rect 122064 6916 122070 6928
rect 123110 6916 123116 6928
rect 122064 6888 123116 6916
rect 122064 6876 122070 6888
rect 123110 6876 123116 6888
rect 123168 6876 123174 6928
rect 114925 6851 114983 6857
rect 114925 6817 114937 6851
rect 114971 6817 114983 6851
rect 114925 6811 114983 6817
rect 115474 6808 115480 6860
rect 115532 6848 115538 6860
rect 116302 6848 116308 6860
rect 115532 6820 116308 6848
rect 115532 6808 115538 6820
rect 116302 6808 116308 6820
rect 116360 6808 116366 6860
rect 116765 6851 116823 6857
rect 116765 6817 116777 6851
rect 116811 6848 116823 6851
rect 116854 6848 116860 6860
rect 116811 6820 116860 6848
rect 116811 6817 116823 6820
rect 116765 6811 116823 6817
rect 116854 6808 116860 6820
rect 116912 6808 116918 6860
rect 118602 6808 118608 6860
rect 118660 6848 118666 6860
rect 118789 6851 118847 6857
rect 118789 6848 118801 6851
rect 118660 6820 118801 6848
rect 118660 6808 118666 6820
rect 118789 6817 118801 6820
rect 118835 6817 118847 6851
rect 121638 6848 121644 6860
rect 121599 6820 121644 6848
rect 118789 6811 118847 6817
rect 121638 6808 121644 6820
rect 121696 6808 121702 6860
rect 122469 6851 122527 6857
rect 122469 6817 122481 6851
rect 122515 6848 122527 6851
rect 122558 6848 122564 6860
rect 122515 6820 122564 6848
rect 122515 6817 122527 6820
rect 122469 6811 122527 6817
rect 122558 6808 122564 6820
rect 122616 6808 122622 6860
rect 124950 6808 124956 6860
rect 125008 6848 125014 6860
rect 125152 6848 125180 6956
rect 125008 6820 125180 6848
rect 125008 6808 125014 6820
rect 125226 6808 125232 6860
rect 125284 6848 125290 6860
rect 125704 6848 125732 6956
rect 126422 6944 126428 6996
rect 126480 6984 126486 6996
rect 126480 6956 129872 6984
rect 126480 6944 126486 6956
rect 126330 6876 126336 6928
rect 126388 6916 126394 6928
rect 127069 6919 127127 6925
rect 127069 6916 127081 6919
rect 126388 6888 127081 6916
rect 126388 6876 126394 6888
rect 127069 6885 127081 6888
rect 127115 6916 127127 6919
rect 128538 6916 128544 6928
rect 127115 6888 128544 6916
rect 127115 6885 127127 6888
rect 127069 6879 127127 6885
rect 128538 6876 128544 6888
rect 128596 6876 128602 6928
rect 129844 6916 129872 6956
rect 129918 6944 129924 6996
rect 129976 6984 129982 6996
rect 130197 6987 130255 6993
rect 130197 6984 130209 6987
rect 129976 6956 130209 6984
rect 129976 6944 129982 6956
rect 130197 6953 130209 6956
rect 130243 6953 130255 6987
rect 130838 6984 130844 6996
rect 130799 6956 130844 6984
rect 130197 6947 130255 6953
rect 130838 6944 130844 6956
rect 130896 6944 130902 6996
rect 130930 6944 130936 6996
rect 130988 6984 130994 6996
rect 133598 6984 133604 6996
rect 130988 6956 133604 6984
rect 130988 6944 130994 6956
rect 133598 6944 133604 6956
rect 133656 6944 133662 6996
rect 133782 6944 133788 6996
rect 133840 6984 133846 6996
rect 134245 6987 134303 6993
rect 134245 6984 134257 6987
rect 133840 6956 134257 6984
rect 133840 6944 133846 6956
rect 134245 6953 134257 6956
rect 134291 6953 134303 6987
rect 134245 6947 134303 6953
rect 134334 6944 134340 6996
rect 134392 6984 134398 6996
rect 137922 6984 137928 6996
rect 134392 6956 137928 6984
rect 134392 6944 134398 6956
rect 137922 6944 137928 6956
rect 137980 6944 137986 6996
rect 138201 6987 138259 6993
rect 138201 6953 138213 6987
rect 138247 6984 138259 6987
rect 138566 6984 138572 6996
rect 138247 6956 138572 6984
rect 138247 6953 138259 6956
rect 138201 6947 138259 6953
rect 138566 6944 138572 6956
rect 138624 6944 138630 6996
rect 138753 6987 138811 6993
rect 138753 6953 138765 6987
rect 138799 6984 138811 6987
rect 139486 6984 139492 6996
rect 138799 6956 139492 6984
rect 138799 6953 138811 6956
rect 138753 6947 138811 6953
rect 139486 6944 139492 6956
rect 139544 6944 139550 6996
rect 139854 6944 139860 6996
rect 139912 6984 139918 6996
rect 146757 6987 146815 6993
rect 139912 6956 146432 6984
rect 139912 6944 139918 6956
rect 132862 6916 132868 6928
rect 129844 6888 132868 6916
rect 132862 6876 132868 6888
rect 132920 6916 132926 6928
rect 135530 6916 135536 6928
rect 132920 6888 135536 6916
rect 132920 6876 132926 6888
rect 135530 6876 135536 6888
rect 135588 6876 135594 6928
rect 140317 6919 140375 6925
rect 140317 6885 140329 6919
rect 140363 6916 140375 6919
rect 141142 6916 141148 6928
rect 140363 6888 141148 6916
rect 140363 6885 140375 6888
rect 140317 6879 140375 6885
rect 141142 6876 141148 6888
rect 141200 6876 141206 6928
rect 143077 6919 143135 6925
rect 143077 6885 143089 6919
rect 143123 6885 143135 6919
rect 143077 6879 143135 6885
rect 128722 6848 128728 6860
rect 125284 6820 125594 6848
rect 125704 6820 128728 6848
rect 125284 6808 125290 6820
rect 111426 6780 111432 6792
rect 111352 6752 111432 6780
rect 111225 6745 111283 6751
rect 111426 6740 111432 6752
rect 111484 6780 111490 6792
rect 114741 6783 114799 6789
rect 111484 6752 111577 6780
rect 111484 6740 111490 6752
rect 114741 6749 114753 6783
rect 114787 6780 114799 6783
rect 114830 6780 114836 6792
rect 114787 6752 114836 6780
rect 114787 6749 114799 6752
rect 114741 6743 114799 6749
rect 114830 6740 114836 6752
rect 114888 6740 114894 6792
rect 115014 6740 115020 6792
rect 115072 6780 115078 6792
rect 118237 6783 118295 6789
rect 118237 6780 118249 6783
rect 115072 6752 118249 6780
rect 115072 6740 115078 6752
rect 118237 6749 118249 6752
rect 118283 6780 118295 6783
rect 118694 6780 118700 6792
rect 118283 6752 118700 6780
rect 118283 6749 118295 6752
rect 118237 6743 118295 6749
rect 118694 6740 118700 6752
rect 118752 6740 118758 6792
rect 119525 6783 119583 6789
rect 119525 6749 119537 6783
rect 119571 6780 119583 6783
rect 120810 6780 120816 6792
rect 119571 6752 120816 6780
rect 119571 6749 119583 6752
rect 119525 6743 119583 6749
rect 120810 6740 120816 6752
rect 120868 6740 120874 6792
rect 122650 6780 122656 6792
rect 121104 6752 121500 6780
rect 122611 6752 122656 6780
rect 111610 6712 111616 6724
rect 108040 6684 111616 6712
rect 111610 6672 111616 6684
rect 111668 6672 111674 6724
rect 115382 6672 115388 6724
rect 115440 6712 115446 6724
rect 121104 6712 121132 6752
rect 115440 6684 121132 6712
rect 121374 6715 121432 6721
rect 115440 6672 115446 6684
rect 121374 6681 121386 6715
rect 121420 6681 121432 6715
rect 121472 6712 121500 6752
rect 122650 6740 122656 6752
rect 122708 6740 122714 6792
rect 122837 6783 122895 6789
rect 122837 6749 122849 6783
rect 122883 6780 122895 6783
rect 123018 6780 123024 6792
rect 122883 6752 123024 6780
rect 122883 6749 122895 6752
rect 122837 6743 122895 6749
rect 123018 6740 123024 6752
rect 123076 6740 123082 6792
rect 124858 6740 124864 6792
rect 124916 6780 124922 6792
rect 124916 6752 124961 6780
rect 124916 6740 124922 6752
rect 125410 6740 125416 6792
rect 125468 6740 125474 6792
rect 125566 6780 125594 6820
rect 128722 6808 128728 6820
rect 128780 6808 128786 6860
rect 129737 6851 129795 6857
rect 129737 6817 129749 6851
rect 129783 6848 129795 6851
rect 129826 6848 129832 6860
rect 129783 6820 129832 6848
rect 129783 6817 129795 6820
rect 129737 6811 129795 6817
rect 129826 6808 129832 6820
rect 129884 6848 129890 6860
rect 130930 6848 130936 6860
rect 129884 6820 130936 6848
rect 129884 6808 129890 6820
rect 130930 6808 130936 6820
rect 130988 6808 130994 6860
rect 132770 6808 132776 6860
rect 132828 6848 132834 6860
rect 133693 6851 133751 6857
rect 133693 6848 133705 6851
rect 132828 6820 133705 6848
rect 132828 6808 132834 6820
rect 133693 6817 133705 6820
rect 133739 6817 133751 6851
rect 133693 6811 133751 6817
rect 138198 6808 138204 6860
rect 138256 6848 138262 6860
rect 142157 6851 142215 6857
rect 138256 6820 139808 6848
rect 138256 6808 138262 6820
rect 128170 6780 128176 6792
rect 125566 6752 128176 6780
rect 128170 6740 128176 6752
rect 128228 6740 128234 6792
rect 129090 6740 129096 6792
rect 129148 6780 129154 6792
rect 129470 6783 129528 6789
rect 129470 6780 129482 6783
rect 129148 6752 129482 6780
rect 129148 6740 129154 6752
rect 129470 6749 129482 6752
rect 129516 6780 129528 6783
rect 130194 6780 130200 6792
rect 129516 6752 130200 6780
rect 129516 6749 129528 6752
rect 129470 6743 129528 6749
rect 130194 6740 130200 6752
rect 130252 6740 130258 6792
rect 132221 6783 132279 6789
rect 132221 6749 132233 6783
rect 132267 6780 132279 6783
rect 133046 6780 133052 6792
rect 132267 6752 133052 6780
rect 132267 6749 132279 6752
rect 132221 6743 132279 6749
rect 133046 6740 133052 6752
rect 133104 6780 133110 6792
rect 133782 6780 133788 6792
rect 133104 6752 133788 6780
rect 133104 6740 133110 6752
rect 133782 6740 133788 6752
rect 133840 6740 133846 6792
rect 135806 6780 135812 6792
rect 134996 6752 135812 6780
rect 124616 6715 124674 6721
rect 121472 6684 123524 6712
rect 121374 6675 121432 6681
rect 91922 6644 91928 6656
rect 86512 6616 89714 6644
rect 91883 6616 91928 6644
rect 91922 6604 91928 6616
rect 91980 6644 91986 6656
rect 92566 6644 92572 6656
rect 91980 6616 92572 6644
rect 91980 6604 91986 6616
rect 92566 6604 92572 6616
rect 92624 6604 92630 6656
rect 93394 6604 93400 6656
rect 93452 6644 93458 6656
rect 96890 6644 96896 6656
rect 93452 6616 96896 6644
rect 93452 6604 93458 6616
rect 96890 6604 96896 6616
rect 96948 6604 96954 6656
rect 97350 6604 97356 6656
rect 97408 6644 97414 6656
rect 106366 6644 106372 6656
rect 97408 6616 106372 6644
rect 97408 6604 97414 6616
rect 106366 6604 106372 6616
rect 106424 6604 106430 6656
rect 107010 6644 107016 6656
rect 106923 6616 107016 6644
rect 107010 6604 107016 6616
rect 107068 6644 107074 6656
rect 115014 6644 115020 6656
rect 107068 6616 115020 6644
rect 107068 6604 107074 6616
rect 115014 6604 115020 6616
rect 115072 6604 115078 6656
rect 117777 6647 117835 6653
rect 117777 6613 117789 6647
rect 117823 6644 117835 6647
rect 118142 6644 118148 6656
rect 117823 6616 118148 6644
rect 117823 6613 117835 6616
rect 117777 6607 117835 6613
rect 118142 6604 118148 6616
rect 118200 6604 118206 6656
rect 119709 6647 119767 6653
rect 119709 6613 119721 6647
rect 119755 6644 119767 6647
rect 120166 6644 120172 6656
rect 119755 6616 120172 6644
rect 119755 6613 119767 6616
rect 119709 6607 119767 6613
rect 120166 6604 120172 6616
rect 120224 6604 120230 6656
rect 120261 6647 120319 6653
rect 120261 6613 120273 6647
rect 120307 6644 120319 6647
rect 121086 6644 121092 6656
rect 120307 6616 121092 6644
rect 120307 6613 120319 6616
rect 120261 6607 120319 6613
rect 121086 6604 121092 6616
rect 121144 6604 121150 6656
rect 121380 6644 121408 6675
rect 121546 6644 121552 6656
rect 121380 6616 121552 6644
rect 121546 6604 121552 6616
rect 121604 6604 121610 6656
rect 121638 6604 121644 6656
rect 121696 6644 121702 6656
rect 123294 6644 123300 6656
rect 121696 6616 123300 6644
rect 121696 6604 121702 6616
rect 123294 6604 123300 6616
rect 123352 6604 123358 6656
rect 123496 6653 123524 6684
rect 124616 6681 124628 6715
rect 124662 6712 124674 6715
rect 125428 6712 125456 6740
rect 129366 6712 129372 6724
rect 124662 6684 124996 6712
rect 125428 6684 129372 6712
rect 124662 6681 124674 6684
rect 124616 6675 124674 6681
rect 123481 6647 123539 6653
rect 123481 6613 123493 6647
rect 123527 6613 123539 6647
rect 124968 6644 124996 6684
rect 129366 6672 129372 6684
rect 129424 6672 129430 6724
rect 131669 6715 131727 6721
rect 131669 6681 131681 6715
rect 131715 6712 131727 6715
rect 133230 6712 133236 6724
rect 131715 6684 133236 6712
rect 131715 6681 131727 6684
rect 131669 6675 131727 6681
rect 125410 6644 125416 6656
rect 124968 6616 125416 6644
rect 123481 6607 123539 6613
rect 125410 6604 125416 6616
rect 125468 6604 125474 6656
rect 125962 6644 125968 6656
rect 125923 6616 125968 6644
rect 125962 6604 125968 6616
rect 126020 6604 126026 6656
rect 126146 6604 126152 6656
rect 126204 6644 126210 6656
rect 126514 6644 126520 6656
rect 126204 6616 126520 6644
rect 126204 6604 126210 6616
rect 126514 6604 126520 6616
rect 126572 6604 126578 6656
rect 127713 6647 127771 6653
rect 127713 6613 127725 6647
rect 127759 6644 127771 6647
rect 127802 6644 127808 6656
rect 127759 6616 127808 6644
rect 127759 6613 127771 6616
rect 127713 6607 127771 6613
rect 127802 6604 127808 6616
rect 127860 6604 127866 6656
rect 128354 6604 128360 6656
rect 128412 6644 128418 6656
rect 128412 6616 128457 6644
rect 128412 6604 128418 6616
rect 129274 6604 129280 6656
rect 129332 6644 129338 6656
rect 131684 6644 131712 6675
rect 133230 6672 133236 6684
rect 133288 6672 133294 6724
rect 133322 6672 133328 6724
rect 133380 6712 133386 6724
rect 134150 6712 134156 6724
rect 133380 6684 134156 6712
rect 133380 6672 133386 6684
rect 134150 6672 134156 6684
rect 134208 6672 134214 6724
rect 129332 6616 131712 6644
rect 133141 6647 133199 6653
rect 129332 6604 129338 6616
rect 133141 6613 133153 6647
rect 133187 6644 133199 6647
rect 133414 6644 133420 6656
rect 133187 6616 133420 6644
rect 133187 6613 133199 6616
rect 133141 6607 133199 6613
rect 133414 6604 133420 6616
rect 133472 6604 133478 6656
rect 133690 6604 133696 6656
rect 133748 6644 133754 6656
rect 134996 6644 135024 6752
rect 135806 6740 135812 6752
rect 135864 6740 135870 6792
rect 136545 6783 136603 6789
rect 136545 6749 136557 6783
rect 136591 6780 136603 6783
rect 136634 6780 136640 6792
rect 136591 6752 136640 6780
rect 136591 6749 136603 6752
rect 136545 6743 136603 6749
rect 136634 6740 136640 6752
rect 136692 6740 136698 6792
rect 139489 6783 139547 6789
rect 139489 6749 139501 6783
rect 139535 6780 139547 6783
rect 139670 6780 139676 6792
rect 139535 6752 139676 6780
rect 139535 6749 139547 6752
rect 139489 6743 139547 6749
rect 139670 6740 139676 6752
rect 139728 6740 139734 6792
rect 135070 6672 135076 6724
rect 135128 6712 135134 6724
rect 136300 6715 136358 6721
rect 135128 6684 135300 6712
rect 135128 6672 135134 6684
rect 135162 6644 135168 6656
rect 133748 6616 135024 6644
rect 135123 6616 135168 6644
rect 133748 6604 133754 6616
rect 135162 6604 135168 6616
rect 135220 6604 135226 6656
rect 135272 6644 135300 6684
rect 136300 6681 136312 6715
rect 136346 6712 136358 6715
rect 137097 6715 137155 6721
rect 137097 6712 137109 6715
rect 136346 6684 137109 6712
rect 136346 6681 136358 6684
rect 136300 6675 136358 6681
rect 137097 6681 137109 6684
rect 137143 6712 137155 6715
rect 139578 6712 139584 6724
rect 137143 6684 139584 6712
rect 137143 6681 137155 6684
rect 137097 6675 137155 6681
rect 139578 6672 139584 6684
rect 139636 6672 139642 6724
rect 139780 6712 139808 6820
rect 142157 6817 142169 6851
rect 142203 6848 142215 6851
rect 142338 6848 142344 6860
rect 142203 6820 142344 6848
rect 142203 6817 142215 6820
rect 142157 6811 142215 6817
rect 142338 6808 142344 6820
rect 142396 6808 142402 6860
rect 142614 6808 142620 6860
rect 142672 6848 142678 6860
rect 143092 6848 143120 6879
rect 142672 6820 143120 6848
rect 146404 6848 146432 6956
rect 146757 6953 146769 6987
rect 146803 6984 146815 6987
rect 147030 6984 147036 6996
rect 146803 6956 147036 6984
rect 146803 6953 146815 6956
rect 146757 6947 146815 6953
rect 147030 6944 147036 6956
rect 147088 6944 147094 6996
rect 148229 6987 148287 6993
rect 148229 6984 148241 6987
rect 147263 6956 148241 6984
rect 146478 6876 146484 6928
rect 146536 6916 146542 6928
rect 147263 6916 147291 6956
rect 148229 6953 148241 6956
rect 148275 6953 148287 6987
rect 148229 6947 148287 6953
rect 148428 6956 149652 6984
rect 146536 6888 147291 6916
rect 146536 6876 146542 6888
rect 148134 6876 148140 6928
rect 148192 6916 148198 6928
rect 148428 6916 148456 6956
rect 148192 6888 148456 6916
rect 148192 6876 148198 6888
rect 148502 6848 148508 6860
rect 146404 6820 148508 6848
rect 142672 6808 142678 6820
rect 148502 6808 148508 6820
rect 148560 6808 148566 6860
rect 149624 6848 149652 6956
rect 150066 6944 150072 6996
rect 150124 6984 150130 6996
rect 156969 6987 157027 6993
rect 156969 6984 156981 6987
rect 150124 6956 156981 6984
rect 150124 6944 150130 6956
rect 156969 6953 156981 6956
rect 157015 6953 157027 6987
rect 156969 6947 157027 6953
rect 149698 6876 149704 6928
rect 149756 6916 149762 6928
rect 150253 6919 150311 6925
rect 150253 6916 150265 6919
rect 149756 6888 150265 6916
rect 149756 6876 149762 6888
rect 150253 6885 150265 6888
rect 150299 6916 150311 6919
rect 151446 6916 151452 6928
rect 150299 6888 150756 6916
rect 151407 6888 151452 6916
rect 150299 6885 150311 6888
rect 150253 6879 150311 6885
rect 150434 6848 150440 6860
rect 149624 6820 150440 6848
rect 150434 6808 150440 6820
rect 150492 6808 150498 6860
rect 150728 6848 150756 6888
rect 151446 6876 151452 6888
rect 151504 6876 151510 6928
rect 152826 6876 152832 6928
rect 152884 6916 152890 6928
rect 153746 6916 153752 6928
rect 152884 6888 153752 6916
rect 152884 6876 152890 6888
rect 153746 6876 153752 6888
rect 153804 6876 153810 6928
rect 152182 6848 152188 6860
rect 150728 6820 152188 6848
rect 152182 6808 152188 6820
rect 152240 6808 152246 6860
rect 155218 6848 155224 6860
rect 154776 6820 155224 6848
rect 140130 6740 140136 6792
rect 140188 6780 140194 6792
rect 140188 6752 140233 6780
rect 140516 6752 142016 6780
rect 140188 6740 140194 6752
rect 140516 6712 140544 6752
rect 139780 6684 140544 6712
rect 141890 6715 141948 6721
rect 141890 6681 141902 6715
rect 141936 6681 141948 6715
rect 141988 6712 142016 6752
rect 142798 6740 142804 6792
rect 142856 6780 142862 6792
rect 143074 6780 143080 6792
rect 142856 6752 143080 6780
rect 142856 6740 142862 6752
rect 143074 6740 143080 6752
rect 143132 6780 143138 6792
rect 143442 6780 143448 6792
rect 143132 6752 143448 6780
rect 143132 6740 143138 6752
rect 143442 6740 143448 6752
rect 143500 6780 143506 6792
rect 144457 6783 144515 6789
rect 144457 6780 144469 6783
rect 143500 6752 144469 6780
rect 143500 6740 143506 6752
rect 144457 6749 144469 6752
rect 144503 6780 144515 6783
rect 145377 6783 145435 6789
rect 145377 6780 145389 6783
rect 144503 6752 145389 6780
rect 144503 6749 144515 6752
rect 144457 6743 144515 6749
rect 145377 6749 145389 6752
rect 145423 6780 145435 6783
rect 146386 6780 146392 6792
rect 145423 6752 146392 6780
rect 145423 6749 145435 6752
rect 145377 6743 145435 6749
rect 146386 6740 146392 6752
rect 146444 6740 146450 6792
rect 146570 6740 146576 6792
rect 146628 6780 146634 6792
rect 147217 6783 147275 6789
rect 147493 6783 147551 6789
rect 147217 6780 147229 6783
rect 146628 6752 147229 6780
rect 146628 6740 146634 6752
rect 147217 6749 147229 6752
rect 147263 6749 147275 6783
rect 147401 6780 147459 6783
rect 147217 6743 147275 6749
rect 147324 6777 147459 6780
rect 147324 6752 147413 6777
rect 144212 6715 144270 6721
rect 141988 6684 143212 6712
rect 141890 6675 141948 6681
rect 139486 6644 139492 6656
rect 135272 6616 139492 6644
rect 139486 6604 139492 6616
rect 139544 6604 139550 6656
rect 139673 6647 139731 6653
rect 139673 6613 139685 6647
rect 139719 6644 139731 6647
rect 139854 6644 139860 6656
rect 139719 6616 139860 6644
rect 139719 6613 139731 6616
rect 139673 6607 139731 6613
rect 139854 6604 139860 6616
rect 139912 6604 139918 6656
rect 140774 6644 140780 6656
rect 140735 6616 140780 6644
rect 140774 6604 140780 6616
rect 140832 6604 140838 6656
rect 141896 6644 141924 6675
rect 143074 6644 143080 6656
rect 141896 6616 143080 6644
rect 143074 6604 143080 6616
rect 143132 6604 143138 6656
rect 143184 6644 143212 6684
rect 144212 6681 144224 6715
rect 144258 6712 144270 6715
rect 145282 6712 145288 6724
rect 144258 6684 145288 6712
rect 144258 6681 144270 6684
rect 144212 6675 144270 6681
rect 145282 6672 145288 6684
rect 145340 6672 145346 6724
rect 145644 6715 145702 6721
rect 145644 6681 145656 6715
rect 145690 6712 145702 6715
rect 146294 6712 146300 6724
rect 145690 6684 146300 6712
rect 145690 6681 145702 6684
rect 145644 6675 145702 6681
rect 146294 6672 146300 6684
rect 146352 6672 146358 6724
rect 147324 6712 147352 6752
rect 147401 6743 147413 6752
rect 147447 6743 147459 6777
rect 147493 6749 147505 6783
rect 147539 6749 147551 6783
rect 147493 6743 147551 6749
rect 147401 6737 147459 6743
rect 146588 6684 147352 6712
rect 146588 6644 146616 6684
rect 143184 6616 146616 6644
rect 147306 6604 147312 6656
rect 147364 6644 147370 6656
rect 147508 6644 147536 6743
rect 147674 6740 147680 6792
rect 147732 6780 147738 6792
rect 149342 6783 149400 6789
rect 149342 6780 149354 6783
rect 147732 6752 149354 6780
rect 147732 6740 147738 6752
rect 149342 6749 149354 6752
rect 149388 6749 149400 6783
rect 149342 6743 149400 6749
rect 149609 6783 149667 6789
rect 149609 6749 149621 6783
rect 149655 6780 149667 6783
rect 149698 6780 149704 6792
rect 149655 6752 149704 6780
rect 149655 6749 149667 6752
rect 149609 6743 149667 6749
rect 149698 6740 149704 6752
rect 149756 6740 149762 6792
rect 150069 6783 150127 6789
rect 150069 6749 150081 6783
rect 150115 6780 150127 6783
rect 150250 6780 150256 6792
rect 150115 6752 150256 6780
rect 150115 6749 150127 6752
rect 150069 6743 150127 6749
rect 150250 6740 150256 6752
rect 150308 6740 150314 6792
rect 150989 6783 151047 6789
rect 150989 6749 151001 6783
rect 151035 6776 151047 6783
rect 151262 6780 151268 6792
rect 151096 6776 151268 6780
rect 151035 6752 151268 6776
rect 151035 6749 151124 6752
rect 150989 6748 151124 6749
rect 150989 6743 151047 6748
rect 151262 6740 151268 6752
rect 151320 6740 151326 6792
rect 151633 6783 151691 6789
rect 151633 6749 151645 6783
rect 151679 6780 151691 6783
rect 151722 6780 151728 6792
rect 151679 6752 151728 6780
rect 151679 6749 151691 6752
rect 151633 6743 151691 6749
rect 151722 6740 151728 6752
rect 151780 6740 151786 6792
rect 152090 6740 152096 6792
rect 152148 6780 152154 6792
rect 152277 6783 152335 6789
rect 152277 6780 152289 6783
rect 152148 6752 152289 6780
rect 152148 6740 152154 6752
rect 152277 6749 152289 6752
rect 152323 6749 152335 6783
rect 152277 6743 152335 6749
rect 152826 6740 152832 6792
rect 152884 6780 152890 6792
rect 154776 6780 154804 6820
rect 155218 6808 155224 6820
rect 155276 6808 155282 6860
rect 155313 6851 155371 6857
rect 155313 6817 155325 6851
rect 155359 6848 155371 6851
rect 155402 6848 155408 6860
rect 155359 6820 155408 6848
rect 155359 6817 155371 6820
rect 155313 6811 155371 6817
rect 155402 6808 155408 6820
rect 155460 6808 155466 6860
rect 156509 6851 156567 6857
rect 156509 6817 156521 6851
rect 156555 6848 156567 6851
rect 156782 6848 156788 6860
rect 156555 6820 156788 6848
rect 156555 6817 156567 6820
rect 156509 6811 156567 6817
rect 156782 6808 156788 6820
rect 156840 6808 156846 6860
rect 152884 6752 154804 6780
rect 154853 6783 154911 6789
rect 152884 6740 152890 6752
rect 154853 6749 154865 6783
rect 154899 6749 154911 6783
rect 155494 6780 155500 6792
rect 155455 6752 155500 6780
rect 154853 6743 154911 6749
rect 147600 6684 150940 6712
rect 147600 6656 147628 6684
rect 147364 6616 147536 6644
rect 147364 6604 147370 6616
rect 147582 6604 147588 6656
rect 147640 6604 147646 6656
rect 147766 6604 147772 6656
rect 147824 6644 147830 6656
rect 150158 6644 150164 6656
rect 147824 6616 150164 6644
rect 147824 6604 147830 6616
rect 150158 6604 150164 6616
rect 150216 6604 150222 6656
rect 150434 6604 150440 6656
rect 150492 6644 150498 6656
rect 150805 6647 150863 6653
rect 150805 6644 150817 6647
rect 150492 6616 150817 6644
rect 150492 6604 150498 6616
rect 150805 6613 150817 6616
rect 150851 6613 150863 6647
rect 150912 6644 150940 6684
rect 152182 6672 152188 6724
rect 152240 6712 152246 6724
rect 152240 6684 154068 6712
rect 152240 6672 152246 6684
rect 152093 6647 152151 6653
rect 152093 6644 152105 6647
rect 150912 6616 152105 6644
rect 150805 6607 150863 6613
rect 152093 6613 152105 6616
rect 152139 6613 152151 6647
rect 152826 6644 152832 6656
rect 152787 6616 152832 6644
rect 152093 6607 152151 6613
rect 152826 6604 152832 6616
rect 152884 6604 152890 6656
rect 153470 6644 153476 6656
rect 153431 6616 153476 6644
rect 153470 6604 153476 6616
rect 153528 6604 153534 6656
rect 154040 6644 154068 6684
rect 154574 6672 154580 6724
rect 154632 6721 154638 6724
rect 154632 6715 154666 6721
rect 154654 6681 154666 6715
rect 154632 6675 154666 6681
rect 154632 6672 154638 6675
rect 154868 6644 154896 6743
rect 155494 6740 155500 6752
rect 155552 6740 155558 6792
rect 156046 6740 156052 6792
rect 156104 6780 156110 6792
rect 156325 6783 156383 6789
rect 156325 6780 156337 6783
rect 156104 6752 156337 6780
rect 156104 6740 156110 6752
rect 156325 6749 156337 6752
rect 156371 6749 156383 6783
rect 156325 6743 156383 6749
rect 157058 6740 157064 6792
rect 157116 6780 157122 6792
rect 157153 6783 157211 6789
rect 157153 6780 157165 6783
rect 157116 6752 157165 6780
rect 157116 6740 157122 6752
rect 157153 6749 157165 6752
rect 157199 6749 157211 6783
rect 157153 6743 157211 6749
rect 157797 6783 157855 6789
rect 157797 6749 157809 6783
rect 157843 6780 157855 6783
rect 157886 6780 157892 6792
rect 157843 6752 157892 6780
rect 157843 6749 157855 6752
rect 157797 6743 157855 6749
rect 157886 6740 157892 6752
rect 157944 6740 157950 6792
rect 155681 6715 155739 6721
rect 155681 6681 155693 6715
rect 155727 6712 155739 6715
rect 157702 6712 157708 6724
rect 155727 6684 157708 6712
rect 155727 6681 155739 6684
rect 155681 6675 155739 6681
rect 157702 6672 157708 6684
rect 157760 6672 157766 6724
rect 154040 6616 154896 6644
rect 155954 6604 155960 6656
rect 156012 6644 156018 6656
rect 156141 6647 156199 6653
rect 156141 6644 156153 6647
rect 156012 6616 156153 6644
rect 156012 6604 156018 6616
rect 156141 6613 156153 6616
rect 156187 6613 156199 6647
rect 157610 6644 157616 6656
rect 157571 6616 157616 6644
rect 156141 6607 156199 6613
rect 157610 6604 157616 6616
rect 157668 6604 157674 6656
rect 1104 6554 159043 6576
rect 1104 6502 40394 6554
rect 40446 6502 40458 6554
rect 40510 6502 40522 6554
rect 40574 6502 40586 6554
rect 40638 6502 40650 6554
rect 40702 6502 79839 6554
rect 79891 6502 79903 6554
rect 79955 6502 79967 6554
rect 80019 6502 80031 6554
rect 80083 6502 80095 6554
rect 80147 6502 119284 6554
rect 119336 6502 119348 6554
rect 119400 6502 119412 6554
rect 119464 6502 119476 6554
rect 119528 6502 119540 6554
rect 119592 6502 158729 6554
rect 158781 6502 158793 6554
rect 158845 6502 158857 6554
rect 158909 6502 158921 6554
rect 158973 6502 158985 6554
rect 159037 6502 159043 6554
rect 1104 6480 159043 6502
rect 8018 6440 8024 6452
rect 7979 6412 8024 6440
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 14918 6400 14924 6452
rect 14976 6440 14982 6452
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 14976 6412 15025 6440
rect 14976 6400 14982 6412
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15654 6440 15660 6452
rect 15615 6412 15660 6440
rect 15013 6403 15071 6409
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 18874 6440 18880 6452
rect 18064 6412 18880 6440
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6304 1642 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 1636 6276 2237 6304
rect 1636 6264 1642 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 8036 6304 8064 6400
rect 17494 6372 17500 6384
rect 16960 6344 17500 6372
rect 16960 6316 16988 6344
rect 17494 6332 17500 6344
rect 17552 6332 17558 6384
rect 18064 6372 18092 6412
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 20070 6440 20076 6452
rect 19383 6412 20076 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 20312 6412 20361 6440
rect 20312 6400 20318 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 21266 6440 21272 6452
rect 21227 6412 21272 6440
rect 20349 6403 20407 6409
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 23750 6440 23756 6452
rect 21508 6412 23756 6440
rect 21508 6400 21514 6412
rect 23750 6400 23756 6412
rect 23808 6400 23814 6452
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6409 23903 6443
rect 37458 6440 37464 6452
rect 23845 6403 23903 6409
rect 25976 6412 37464 6440
rect 17972 6344 18092 6372
rect 18141 6375 18199 6381
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 8036 6276 9321 6304
rect 2225 6267 2283 6273
rect 9309 6273 9321 6276
rect 9355 6304 9367 6307
rect 13998 6304 14004 6316
rect 9355 6276 12434 6304
rect 13911 6276 14004 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 8662 6236 8668 6248
rect 8575 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 8720 6208 9505 6236
rect 8720 6196 8726 6208
rect 9493 6205 9505 6208
rect 9539 6236 9551 6239
rect 11146 6236 11152 6248
rect 9539 6208 11152 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 12406 6236 12434 6276
rect 13998 6264 14004 6276
rect 14056 6304 14062 6316
rect 15010 6304 15016 6316
rect 14056 6276 15016 6304
rect 14056 6264 14062 6276
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15194 6304 15200 6316
rect 15155 6276 15200 6304
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15712 6276 15853 6304
rect 15712 6264 15718 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 16942 6304 16948 6316
rect 16903 6276 16948 6304
rect 15841 6267 15899 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17972 6313 18000 6344
rect 18141 6341 18153 6375
rect 18187 6372 18199 6375
rect 20990 6372 20996 6384
rect 18187 6344 20996 6372
rect 18187 6341 18199 6344
rect 18141 6335 18199 6341
rect 20990 6332 20996 6344
rect 21048 6332 21054 6384
rect 23860 6372 23888 6403
rect 21744 6344 23888 6372
rect 17773 6307 17831 6313
rect 17773 6304 17785 6307
rect 17092 6276 17785 6304
rect 17092 6264 17098 6276
rect 17773 6273 17785 6276
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18104 6276 18613 6304
rect 18104 6264 18110 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 21085 6307 21143 6313
rect 18840 6276 21036 6304
rect 18840 6264 18846 6276
rect 17494 6236 17500 6248
rect 12406 6208 17500 6236
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18564 6208 20300 6236
rect 18564 6196 18570 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 9306 6168 9312 6180
rect 1811 6140 9312 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 14553 6171 14611 6177
rect 14553 6137 14565 6171
rect 14599 6168 14611 6171
rect 15286 6168 15292 6180
rect 14599 6140 15292 6168
rect 14599 6137 14611 6140
rect 14553 6131 14611 6137
rect 15286 6128 15292 6140
rect 15344 6168 15350 6180
rect 18785 6171 18843 6177
rect 15344 6140 17816 6168
rect 15344 6128 15350 6140
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 5994 6100 6000 6112
rect 5583 6072 6000 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 17034 6100 17040 6112
rect 12308 6072 17040 6100
rect 12308 6060 12314 6072
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 17221 6103 17279 6109
rect 17221 6069 17233 6103
rect 17267 6100 17279 6103
rect 17678 6100 17684 6112
rect 17267 6072 17684 6100
rect 17267 6069 17279 6072
rect 17221 6063 17279 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17788 6100 17816 6140
rect 18785 6137 18797 6171
rect 18831 6168 18843 6171
rect 19334 6168 19340 6180
rect 18831 6140 19340 6168
rect 18831 6137 18843 6140
rect 18785 6131 18843 6137
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 20272 6168 20300 6208
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 20404 6208 20913 6236
rect 20404 6196 20410 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 21008 6236 21036 6276
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21634 6304 21640 6316
rect 21131 6276 21640 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 21744 6236 21772 6344
rect 23934 6332 23940 6384
rect 23992 6372 23998 6384
rect 23992 6344 25728 6372
rect 23992 6332 23998 6344
rect 22186 6304 22192 6316
rect 22147 6276 22192 6304
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 25700 6313 25728 6344
rect 25976 6313 26004 6412
rect 37458 6400 37464 6412
rect 37516 6400 37522 6452
rect 37550 6400 37556 6452
rect 37608 6440 37614 6452
rect 37829 6443 37887 6449
rect 37829 6440 37841 6443
rect 37608 6412 37841 6440
rect 37608 6400 37614 6412
rect 37829 6409 37841 6412
rect 37875 6440 37887 6443
rect 38378 6440 38384 6452
rect 37875 6412 38384 6440
rect 37875 6409 37887 6412
rect 37829 6403 37887 6409
rect 38378 6400 38384 6412
rect 38436 6400 38442 6452
rect 40589 6443 40647 6449
rect 40589 6409 40601 6443
rect 40635 6440 40647 6443
rect 41230 6440 41236 6452
rect 40635 6412 41236 6440
rect 40635 6409 40647 6412
rect 40589 6403 40647 6409
rect 41230 6400 41236 6412
rect 41288 6400 41294 6452
rect 44637 6443 44695 6449
rect 44637 6440 44649 6443
rect 41386 6412 44649 6440
rect 27614 6332 27620 6384
rect 27672 6372 27678 6384
rect 28813 6375 28871 6381
rect 28813 6372 28825 6375
rect 27672 6344 28825 6372
rect 27672 6332 27678 6344
rect 28813 6341 28825 6344
rect 28859 6372 28871 6375
rect 30478 6375 30536 6381
rect 30478 6372 30490 6375
rect 28859 6344 30490 6372
rect 28859 6341 28871 6344
rect 28813 6335 28871 6341
rect 30478 6341 30490 6344
rect 30524 6341 30536 6375
rect 30478 6335 30536 6341
rect 33536 6375 33594 6381
rect 33536 6341 33548 6375
rect 33582 6372 33594 6375
rect 36354 6372 36360 6384
rect 33582 6344 36360 6372
rect 33582 6341 33594 6344
rect 33536 6335 33594 6341
rect 36354 6332 36360 6344
rect 36412 6332 36418 6384
rect 36464 6344 40448 6372
rect 24958 6307 25016 6313
rect 24958 6304 24970 6307
rect 23492 6276 24970 6304
rect 22002 6236 22008 6248
rect 21008 6208 21772 6236
rect 21963 6208 22008 6236
rect 20901 6199 20959 6205
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 23290 6168 23296 6180
rect 20272 6140 23296 6168
rect 23290 6128 23296 6140
rect 23348 6168 23354 6180
rect 23492 6168 23520 6276
rect 24958 6273 24970 6276
rect 25004 6273 25016 6307
rect 24958 6267 25016 6273
rect 25685 6307 25743 6313
rect 25685 6273 25697 6307
rect 25731 6273 25743 6307
rect 25685 6267 25743 6273
rect 25961 6307 26019 6313
rect 25961 6273 25973 6307
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 30190 6264 30196 6316
rect 30248 6304 30254 6316
rect 30745 6307 30803 6313
rect 30745 6304 30757 6307
rect 30248 6276 30757 6304
rect 30248 6264 30254 6276
rect 30745 6273 30757 6276
rect 30791 6273 30803 6307
rect 32398 6304 32404 6316
rect 32311 6276 32404 6304
rect 30745 6267 30803 6273
rect 32398 6264 32404 6276
rect 32456 6304 32462 6316
rect 36464 6304 36492 6344
rect 32456 6276 36492 6304
rect 38381 6307 38439 6313
rect 32456 6264 32462 6276
rect 38381 6273 38393 6307
rect 38427 6304 38439 6307
rect 38470 6304 38476 6316
rect 38427 6276 38476 6304
rect 38427 6273 38439 6276
rect 38381 6267 38439 6273
rect 38470 6264 38476 6276
rect 38528 6264 38534 6316
rect 38654 6313 38660 6316
rect 38648 6267 38660 6313
rect 38712 6304 38718 6316
rect 40218 6304 40224 6316
rect 38712 6276 38748 6304
rect 40179 6276 40224 6304
rect 38654 6264 38660 6267
rect 38712 6264 38718 6276
rect 40218 6264 40224 6276
rect 40276 6264 40282 6316
rect 40420 6313 40448 6344
rect 40862 6332 40868 6384
rect 40920 6372 40926 6384
rect 41386 6372 41414 6412
rect 44637 6409 44649 6412
rect 44683 6409 44695 6443
rect 44637 6403 44695 6409
rect 44726 6400 44732 6452
rect 44784 6440 44790 6452
rect 46014 6440 46020 6452
rect 44784 6412 46020 6440
rect 44784 6400 44790 6412
rect 46014 6400 46020 6412
rect 46072 6400 46078 6452
rect 46477 6443 46535 6449
rect 46477 6409 46489 6443
rect 46523 6409 46535 6443
rect 46477 6403 46535 6409
rect 46492 6372 46520 6403
rect 46566 6400 46572 6452
rect 46624 6440 46630 6452
rect 52362 6440 52368 6452
rect 46624 6412 52368 6440
rect 46624 6400 46630 6412
rect 52362 6400 52368 6412
rect 52420 6400 52426 6452
rect 53190 6440 53196 6452
rect 53151 6412 53196 6440
rect 53190 6400 53196 6412
rect 53248 6400 53254 6452
rect 54113 6443 54171 6449
rect 54113 6440 54125 6443
rect 53300 6412 54125 6440
rect 40920 6344 41414 6372
rect 43824 6344 46520 6372
rect 40920 6332 40926 6344
rect 40405 6307 40463 6313
rect 40405 6273 40417 6307
rect 40451 6273 40463 6307
rect 41049 6307 41107 6313
rect 41049 6304 41061 6307
rect 40405 6267 40463 6273
rect 40880 6276 41061 6304
rect 25225 6239 25283 6245
rect 25225 6205 25237 6239
rect 25271 6236 25283 6239
rect 26326 6236 26332 6248
rect 25271 6208 26332 6236
rect 25271 6205 25283 6208
rect 25225 6199 25283 6205
rect 26326 6196 26332 6208
rect 26384 6196 26390 6248
rect 29362 6168 29368 6180
rect 23348 6140 23520 6168
rect 29323 6140 29368 6168
rect 23348 6128 23354 6140
rect 29362 6128 29368 6140
rect 29420 6128 29426 6180
rect 32416 6177 32444 6264
rect 33778 6236 33784 6248
rect 33739 6208 33784 6236
rect 33778 6196 33784 6208
rect 33836 6196 33842 6248
rect 40236 6236 40264 6264
rect 40880 6236 40908 6276
rect 41049 6273 41061 6276
rect 41095 6304 41107 6307
rect 43530 6304 43536 6316
rect 41095 6276 43536 6304
rect 41095 6273 41107 6276
rect 41049 6267 41107 6273
rect 43530 6264 43536 6276
rect 43588 6264 43594 6316
rect 40236 6208 40908 6236
rect 40954 6196 40960 6248
rect 41012 6236 41018 6248
rect 43824 6236 43852 6344
rect 50706 6332 50712 6384
rect 50764 6372 50770 6384
rect 50764 6344 51764 6372
rect 50764 6332 50770 6344
rect 45750 6307 45808 6313
rect 45750 6304 45762 6307
rect 41012 6208 43852 6236
rect 44192 6276 45762 6304
rect 41012 6196 41018 6208
rect 32401 6171 32459 6177
rect 32401 6137 32413 6171
rect 32447 6137 32459 6171
rect 32401 6131 32459 6137
rect 33962 6128 33968 6180
rect 34020 6168 34026 6180
rect 38010 6168 38016 6180
rect 34020 6140 38016 6168
rect 34020 6128 34026 6140
rect 38010 6128 38016 6140
rect 38068 6128 38074 6180
rect 39761 6171 39819 6177
rect 39761 6137 39773 6171
rect 39807 6168 39819 6171
rect 39807 6140 41184 6168
rect 39807 6137 39819 6140
rect 39761 6131 39819 6137
rect 19978 6100 19984 6112
rect 17788 6072 19984 6100
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 22186 6100 22192 6112
rect 20312 6072 22192 6100
rect 20312 6060 20318 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22370 6100 22376 6112
rect 22331 6072 22376 6100
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 30834 6100 30840 6112
rect 23808 6072 30840 6100
rect 23808 6060 23814 6072
rect 30834 6060 30840 6072
rect 30892 6060 30898 6112
rect 33502 6060 33508 6112
rect 33560 6100 33566 6112
rect 34241 6103 34299 6109
rect 34241 6100 34253 6103
rect 33560 6072 34253 6100
rect 33560 6060 33566 6072
rect 34241 6069 34253 6072
rect 34287 6069 34299 6103
rect 34241 6063 34299 6069
rect 34974 6060 34980 6112
rect 35032 6100 35038 6112
rect 39776 6100 39804 6131
rect 35032 6072 39804 6100
rect 41156 6100 41184 6140
rect 41230 6128 41236 6180
rect 41288 6168 41294 6180
rect 44192 6177 44220 6276
rect 45750 6273 45762 6276
rect 45796 6273 45808 6307
rect 45750 6267 45808 6273
rect 45922 6264 45928 6316
rect 45980 6304 45986 6316
rect 46658 6304 46664 6316
rect 45980 6276 46152 6304
rect 46619 6276 46664 6304
rect 45980 6264 45986 6276
rect 46014 6236 46020 6248
rect 45975 6208 46020 6236
rect 46014 6196 46020 6208
rect 46072 6196 46078 6248
rect 46124 6236 46152 6276
rect 46658 6264 46664 6276
rect 46716 6264 46722 6316
rect 50798 6264 50804 6316
rect 50856 6304 50862 6316
rect 51629 6307 51687 6313
rect 51629 6304 51641 6307
rect 50856 6276 51641 6304
rect 50856 6264 50862 6276
rect 51629 6273 51641 6276
rect 51675 6273 51687 6307
rect 51629 6267 51687 6273
rect 48590 6236 48596 6248
rect 46124 6208 48596 6236
rect 48590 6196 48596 6208
rect 48648 6196 48654 6248
rect 51445 6239 51503 6245
rect 51445 6205 51457 6239
rect 51491 6236 51503 6239
rect 51736 6236 51764 6344
rect 51810 6332 51816 6384
rect 51868 6372 51874 6384
rect 53300 6372 53328 6412
rect 54113 6409 54125 6412
rect 54159 6409 54171 6443
rect 59722 6440 59728 6452
rect 59683 6412 59728 6440
rect 54113 6403 54171 6409
rect 59722 6400 59728 6412
rect 59780 6400 59786 6452
rect 63494 6400 63500 6452
rect 63552 6440 63558 6452
rect 63589 6443 63647 6449
rect 63589 6440 63601 6443
rect 63552 6412 63601 6440
rect 63552 6400 63558 6412
rect 63589 6409 63601 6412
rect 63635 6409 63647 6443
rect 63589 6403 63647 6409
rect 64046 6400 64052 6452
rect 64104 6440 64110 6452
rect 64141 6443 64199 6449
rect 64141 6440 64153 6443
rect 64104 6412 64153 6440
rect 64104 6400 64110 6412
rect 64141 6409 64153 6412
rect 64187 6409 64199 6443
rect 64141 6403 64199 6409
rect 64414 6400 64420 6452
rect 64472 6440 64478 6452
rect 65886 6440 65892 6452
rect 64472 6412 65892 6440
rect 64472 6400 64478 6412
rect 65886 6400 65892 6412
rect 65944 6400 65950 6452
rect 66070 6440 66076 6452
rect 66031 6412 66076 6440
rect 66070 6400 66076 6412
rect 66128 6400 66134 6452
rect 66530 6400 66536 6452
rect 66588 6440 66594 6452
rect 66625 6443 66683 6449
rect 66625 6440 66637 6443
rect 66588 6412 66637 6440
rect 66588 6400 66594 6412
rect 66625 6409 66637 6412
rect 66671 6440 66683 6443
rect 69106 6440 69112 6452
rect 66671 6412 69112 6440
rect 66671 6409 66683 6412
rect 66625 6403 66683 6409
rect 69106 6400 69112 6412
rect 69164 6440 69170 6452
rect 69293 6443 69351 6449
rect 69293 6440 69305 6443
rect 69164 6412 69305 6440
rect 69164 6400 69170 6412
rect 69293 6409 69305 6412
rect 69339 6409 69351 6443
rect 72878 6440 72884 6452
rect 72839 6412 72884 6440
rect 69293 6403 69351 6409
rect 68922 6372 68928 6384
rect 51868 6344 53328 6372
rect 54036 6344 68928 6372
rect 51868 6332 51874 6344
rect 53374 6304 53380 6316
rect 53335 6276 53380 6304
rect 53374 6264 53380 6276
rect 53432 6264 53438 6316
rect 52273 6239 52331 6245
rect 52273 6236 52285 6239
rect 51491 6208 52285 6236
rect 51491 6205 51503 6208
rect 51445 6199 51503 6205
rect 52273 6205 52285 6208
rect 52319 6205 52331 6239
rect 54036 6236 54064 6344
rect 68922 6332 68928 6344
rect 68980 6332 68986 6384
rect 54110 6264 54116 6316
rect 54168 6304 54174 6316
rect 55226 6307 55284 6313
rect 55226 6304 55238 6307
rect 54168 6276 55238 6304
rect 54168 6264 54174 6276
rect 55226 6273 55238 6276
rect 55272 6273 55284 6307
rect 55226 6267 55284 6273
rect 55398 6264 55404 6316
rect 55456 6304 55462 6316
rect 55493 6307 55551 6313
rect 55493 6304 55505 6307
rect 55456 6276 55505 6304
rect 55456 6264 55462 6276
rect 55493 6273 55505 6276
rect 55539 6273 55551 6307
rect 55493 6267 55551 6273
rect 56505 6307 56563 6313
rect 56505 6273 56517 6307
rect 56551 6273 56563 6307
rect 56505 6267 56563 6273
rect 65265 6307 65323 6313
rect 65265 6273 65277 6307
rect 65311 6304 65323 6307
rect 66809 6307 66867 6313
rect 65311 6276 66760 6304
rect 65311 6273 65323 6276
rect 65265 6267 65323 6273
rect 54036 6208 54331 6236
rect 52273 6199 52331 6205
rect 44177 6171 44235 6177
rect 44177 6168 44189 6171
rect 41288 6140 44189 6168
rect 41288 6128 41294 6140
rect 44177 6137 44189 6140
rect 44223 6137 44235 6171
rect 44177 6131 44235 6137
rect 50246 6128 50252 6180
rect 50304 6168 50310 6180
rect 51813 6171 51871 6177
rect 50304 6140 51074 6168
rect 50304 6128 50310 6140
rect 46198 6100 46204 6112
rect 41156 6072 46204 6100
rect 35032 6060 35038 6072
rect 46198 6060 46204 6072
rect 46256 6060 46262 6112
rect 50798 6060 50804 6112
rect 50856 6100 50862 6112
rect 50893 6103 50951 6109
rect 50893 6100 50905 6103
rect 50856 6072 50905 6100
rect 50856 6060 50862 6072
rect 50893 6069 50905 6072
rect 50939 6069 50951 6103
rect 51046 6100 51074 6140
rect 51813 6137 51825 6171
rect 51859 6168 51871 6171
rect 54202 6168 54208 6180
rect 51859 6140 54208 6168
rect 51859 6137 51871 6140
rect 51813 6131 51871 6137
rect 54202 6128 54208 6140
rect 54260 6128 54266 6180
rect 54303 6100 54331 6208
rect 51046 6072 54331 6100
rect 50893 6063 50951 6069
rect 54846 6060 54852 6112
rect 54904 6100 54910 6112
rect 56520 6100 56548 6267
rect 65521 6239 65579 6245
rect 65521 6205 65533 6239
rect 65567 6205 65579 6239
rect 65521 6199 65579 6205
rect 56689 6171 56747 6177
rect 56689 6137 56701 6171
rect 56735 6168 56747 6171
rect 63954 6168 63960 6180
rect 56735 6140 63960 6168
rect 56735 6137 56747 6140
rect 56689 6131 56747 6137
rect 63954 6128 63960 6140
rect 64012 6128 64018 6180
rect 54904 6072 56548 6100
rect 54904 6060 54910 6072
rect 63494 6060 63500 6112
rect 63552 6100 63558 6112
rect 65536 6100 65564 6199
rect 66732 6168 66760 6276
rect 66809 6273 66821 6307
rect 66855 6304 66867 6307
rect 67269 6307 67327 6313
rect 67269 6304 67281 6307
rect 66855 6276 67281 6304
rect 66855 6273 66867 6276
rect 66809 6267 66867 6273
rect 67269 6273 67281 6276
rect 67315 6304 67327 6307
rect 68370 6304 68376 6316
rect 67315 6276 68376 6304
rect 67315 6273 67327 6276
rect 67269 6267 67327 6273
rect 68370 6264 68376 6276
rect 68428 6264 68434 6316
rect 69308 6304 69336 6403
rect 72878 6400 72884 6412
rect 72936 6400 72942 6452
rect 73798 6440 73804 6452
rect 73759 6412 73804 6440
rect 73798 6400 73804 6412
rect 73856 6400 73862 6452
rect 74994 6440 75000 6452
rect 74955 6412 75000 6440
rect 74994 6400 75000 6412
rect 75052 6400 75058 6452
rect 78858 6440 78864 6452
rect 78819 6412 78864 6440
rect 78858 6400 78864 6412
rect 78916 6400 78922 6452
rect 79318 6400 79324 6452
rect 79376 6440 79382 6452
rect 80606 6440 80612 6452
rect 79376 6412 80612 6440
rect 79376 6400 79382 6412
rect 80606 6400 80612 6412
rect 80664 6400 80670 6452
rect 81066 6400 81072 6452
rect 81124 6440 81130 6452
rect 82630 6440 82636 6452
rect 81124 6412 82636 6440
rect 81124 6400 81130 6412
rect 82630 6400 82636 6412
rect 82688 6400 82694 6452
rect 85574 6400 85580 6452
rect 85632 6440 85638 6452
rect 85669 6443 85727 6449
rect 85669 6440 85681 6443
rect 85632 6412 85681 6440
rect 85632 6400 85638 6412
rect 85669 6409 85681 6412
rect 85715 6409 85727 6443
rect 89438 6440 89444 6452
rect 85669 6403 85727 6409
rect 87248 6412 89444 6440
rect 70112 6375 70170 6381
rect 70112 6341 70124 6375
rect 70158 6372 70170 6375
rect 71777 6375 71835 6381
rect 71777 6372 71789 6375
rect 70158 6344 71789 6372
rect 70158 6341 70170 6344
rect 70112 6335 70170 6341
rect 71777 6341 71789 6344
rect 71823 6372 71835 6375
rect 87248 6372 87276 6412
rect 89438 6400 89444 6412
rect 89496 6400 89502 6452
rect 92198 6400 92204 6452
rect 92256 6440 92262 6452
rect 94498 6440 94504 6452
rect 92256 6412 94504 6440
rect 92256 6400 92262 6412
rect 94498 6400 94504 6412
rect 94556 6400 94562 6452
rect 102134 6400 102140 6452
rect 102192 6440 102198 6452
rect 106458 6440 106464 6452
rect 102192 6412 105400 6440
rect 106419 6412 106464 6440
rect 102192 6400 102198 6412
rect 105372 6381 105400 6412
rect 106458 6400 106464 6412
rect 106516 6400 106522 6452
rect 108758 6440 108764 6452
rect 108719 6412 108764 6440
rect 108758 6400 108764 6412
rect 108816 6400 108822 6452
rect 108850 6400 108856 6452
rect 108908 6440 108914 6452
rect 109589 6443 109647 6449
rect 109589 6440 109601 6443
rect 108908 6412 109601 6440
rect 108908 6400 108914 6412
rect 109589 6409 109601 6412
rect 109635 6440 109647 6443
rect 111334 6440 111340 6452
rect 109635 6412 111340 6440
rect 109635 6409 109647 6412
rect 109589 6403 109647 6409
rect 111334 6400 111340 6412
rect 111392 6400 111398 6452
rect 111610 6400 111616 6452
rect 111668 6440 111674 6452
rect 117130 6440 117136 6452
rect 111668 6412 116164 6440
rect 117091 6412 117136 6440
rect 111668 6400 111674 6412
rect 71823 6344 87276 6372
rect 87356 6375 87414 6381
rect 71823 6341 71835 6344
rect 71777 6335 71835 6341
rect 87356 6341 87368 6375
rect 87402 6372 87414 6375
rect 88153 6375 88211 6381
rect 88153 6372 88165 6375
rect 87402 6344 88165 6372
rect 87402 6341 87414 6344
rect 87356 6335 87414 6341
rect 88153 6341 88165 6344
rect 88199 6372 88211 6375
rect 105348 6375 105406 6381
rect 88199 6344 105308 6372
rect 88199 6341 88211 6344
rect 88153 6335 88211 6341
rect 69845 6307 69903 6313
rect 69845 6304 69857 6307
rect 69308 6276 69857 6304
rect 69845 6273 69857 6276
rect 69891 6273 69903 6307
rect 69845 6267 69903 6273
rect 73890 6264 73896 6316
rect 73948 6304 73954 6316
rect 75086 6304 75092 6316
rect 73948 6276 75092 6304
rect 73948 6264 73954 6276
rect 75086 6264 75092 6276
rect 75144 6264 75150 6316
rect 76121 6307 76179 6313
rect 76121 6273 76133 6307
rect 76167 6304 76179 6307
rect 76929 6307 76987 6313
rect 76929 6304 76941 6307
rect 76167 6276 76941 6304
rect 76167 6273 76179 6276
rect 76121 6267 76179 6273
rect 76929 6273 76941 6276
rect 76975 6304 76987 6307
rect 89622 6304 89628 6316
rect 76975 6276 89628 6304
rect 76975 6273 76987 6276
rect 76929 6267 76987 6273
rect 89622 6264 89628 6276
rect 89680 6264 89686 6316
rect 89800 6307 89858 6313
rect 89800 6273 89812 6307
rect 89846 6304 89858 6307
rect 91462 6304 91468 6316
rect 89846 6276 91468 6304
rect 89846 6273 89858 6276
rect 89800 6267 89858 6273
rect 91462 6264 91468 6276
rect 91520 6264 91526 6316
rect 92109 6307 92167 6313
rect 92109 6304 92121 6307
rect 91563 6276 92121 6304
rect 76377 6239 76435 6245
rect 76377 6205 76389 6239
rect 76423 6236 76435 6239
rect 76466 6236 76472 6248
rect 76423 6208 76472 6236
rect 76423 6205 76435 6208
rect 76377 6199 76435 6205
rect 76466 6196 76472 6208
rect 76524 6236 76530 6248
rect 77110 6236 77116 6248
rect 76524 6208 77116 6236
rect 76524 6196 76530 6208
rect 77110 6196 77116 6208
rect 77168 6236 77174 6248
rect 80422 6236 80428 6248
rect 77168 6208 80428 6236
rect 77168 6196 77174 6208
rect 80422 6196 80428 6208
rect 80480 6236 80486 6248
rect 81066 6236 81072 6248
rect 80480 6208 81072 6236
rect 80480 6196 80486 6208
rect 81066 6196 81072 6208
rect 81124 6196 81130 6248
rect 87601 6239 87659 6245
rect 87601 6205 87613 6239
rect 87647 6236 87659 6239
rect 88426 6236 88432 6248
rect 87647 6208 88432 6236
rect 87647 6205 87659 6208
rect 87601 6199 87659 6205
rect 71225 6171 71283 6177
rect 66732 6140 69428 6168
rect 63552 6072 65564 6100
rect 69400 6100 69428 6140
rect 71225 6137 71237 6171
rect 71271 6168 71283 6171
rect 79134 6168 79140 6180
rect 71271 6140 75500 6168
rect 71271 6137 71283 6140
rect 71225 6131 71283 6137
rect 73706 6100 73712 6112
rect 69400 6072 73712 6100
rect 63552 6060 63558 6072
rect 73706 6060 73712 6072
rect 73764 6060 73770 6112
rect 75472 6100 75500 6140
rect 76392 6140 79140 6168
rect 76392 6100 76420 6140
rect 79134 6128 79140 6140
rect 79192 6128 79198 6180
rect 80698 6128 80704 6180
rect 80756 6168 80762 6180
rect 86221 6171 86279 6177
rect 86221 6168 86233 6171
rect 80756 6140 86233 6168
rect 80756 6128 80762 6140
rect 86221 6137 86233 6140
rect 86267 6137 86279 6171
rect 86221 6131 86279 6137
rect 75472 6072 76420 6100
rect 85574 6060 85580 6112
rect 85632 6100 85638 6112
rect 87616 6100 87644 6199
rect 88426 6196 88432 6208
rect 88484 6236 88490 6248
rect 88981 6239 89039 6245
rect 88981 6236 88993 6239
rect 88484 6208 88993 6236
rect 88484 6196 88490 6208
rect 88981 6205 88993 6208
rect 89027 6236 89039 6239
rect 89530 6236 89536 6248
rect 89027 6208 89536 6236
rect 89027 6205 89039 6208
rect 88981 6199 89039 6205
rect 89530 6196 89536 6208
rect 89588 6196 89594 6248
rect 90542 6196 90548 6248
rect 90600 6236 90606 6248
rect 91563 6236 91591 6276
rect 92109 6273 92121 6276
rect 92155 6304 92167 6307
rect 93210 6304 93216 6316
rect 92155 6276 93216 6304
rect 92155 6273 92167 6276
rect 92109 6267 92167 6273
rect 93210 6264 93216 6276
rect 93268 6264 93274 6316
rect 97350 6313 97356 6316
rect 97344 6304 97356 6313
rect 97311 6276 97356 6304
rect 97344 6267 97356 6276
rect 97350 6264 97356 6267
rect 97408 6264 97414 6316
rect 101582 6304 101588 6316
rect 101543 6276 101588 6304
rect 101582 6264 101588 6276
rect 101640 6264 101646 6316
rect 101858 6304 101864 6316
rect 101819 6276 101864 6304
rect 101858 6264 101864 6276
rect 101916 6264 101922 6316
rect 105081 6307 105139 6313
rect 105081 6273 105093 6307
rect 105127 6304 105139 6307
rect 105170 6304 105176 6316
rect 105127 6276 105176 6304
rect 105127 6273 105139 6276
rect 105081 6267 105139 6273
rect 105170 6264 105176 6276
rect 105228 6264 105234 6316
rect 105280 6304 105308 6344
rect 105348 6341 105360 6375
rect 105394 6341 105406 6375
rect 105348 6335 105406 6341
rect 107194 6332 107200 6384
rect 107252 6372 107258 6384
rect 107626 6375 107684 6381
rect 107626 6372 107638 6375
rect 107252 6344 107638 6372
rect 107252 6332 107258 6344
rect 107626 6341 107638 6344
rect 107672 6341 107684 6375
rect 107626 6335 107684 6341
rect 107838 6332 107844 6384
rect 107896 6372 107902 6384
rect 108868 6372 108896 6400
rect 110690 6372 110696 6384
rect 107896 6344 108896 6372
rect 109006 6344 110696 6372
rect 107896 6332 107902 6344
rect 107010 6304 107016 6316
rect 105280 6276 107016 6304
rect 107010 6264 107016 6276
rect 107068 6264 107074 6316
rect 107378 6304 107384 6316
rect 107339 6276 107384 6304
rect 107378 6264 107384 6276
rect 107436 6264 107442 6316
rect 90600 6208 91591 6236
rect 90600 6196 90606 6208
rect 91830 6196 91836 6248
rect 91888 6236 91894 6248
rect 91925 6239 91983 6245
rect 91925 6236 91937 6239
rect 91888 6208 91937 6236
rect 91888 6196 91894 6208
rect 91925 6205 91937 6208
rect 91971 6236 91983 6239
rect 94038 6236 94044 6248
rect 91971 6208 94044 6236
rect 91971 6205 91983 6208
rect 91925 6199 91983 6205
rect 94038 6196 94044 6208
rect 94096 6196 94102 6248
rect 96614 6196 96620 6248
rect 96672 6236 96678 6248
rect 97077 6239 97135 6245
rect 97077 6236 97089 6239
rect 96672 6208 97089 6236
rect 96672 6196 96678 6208
rect 97077 6205 97089 6208
rect 97123 6205 97135 6239
rect 100754 6236 100760 6248
rect 97077 6199 97135 6205
rect 98472 6208 100760 6236
rect 98472 6177 98500 6208
rect 100754 6196 100760 6208
rect 100812 6196 100818 6248
rect 100846 6196 100852 6248
rect 100904 6236 100910 6248
rect 100941 6239 100999 6245
rect 100941 6236 100953 6239
rect 100904 6208 100953 6236
rect 100904 6196 100910 6208
rect 100941 6205 100953 6208
rect 100987 6236 100999 6239
rect 101876 6236 101904 6264
rect 100987 6208 101904 6236
rect 100987 6205 100999 6208
rect 100941 6199 100999 6205
rect 106090 6196 106096 6248
rect 106148 6236 106154 6248
rect 107102 6236 107108 6248
rect 106148 6208 107108 6236
rect 106148 6196 106154 6208
rect 107102 6196 107108 6208
rect 107160 6196 107166 6248
rect 109006 6236 109034 6344
rect 110690 6332 110696 6344
rect 110748 6332 110754 6384
rect 111245 6375 111303 6381
rect 111245 6341 111257 6375
rect 111291 6372 111303 6375
rect 111426 6372 111432 6384
rect 111291 6344 111432 6372
rect 111291 6341 111303 6344
rect 111245 6335 111303 6341
rect 111426 6332 111432 6344
rect 111484 6332 111490 6384
rect 111978 6332 111984 6384
rect 112036 6372 112042 6384
rect 116136 6372 116164 6412
rect 117130 6400 117136 6412
rect 117188 6400 117194 6452
rect 119893 6443 119951 6449
rect 119893 6440 119905 6443
rect 118666 6412 119905 6440
rect 118666 6372 118694 6412
rect 119893 6409 119905 6412
rect 119939 6409 119951 6443
rect 119893 6403 119951 6409
rect 120534 6400 120540 6452
rect 120592 6440 120598 6452
rect 121638 6440 121644 6452
rect 120592 6412 121644 6440
rect 120592 6400 120598 6412
rect 121638 6400 121644 6412
rect 121696 6400 121702 6452
rect 121733 6443 121791 6449
rect 121733 6409 121745 6443
rect 121779 6409 121791 6443
rect 121733 6403 121791 6409
rect 112036 6344 116072 6372
rect 116136 6344 118694 6372
rect 112036 6332 112042 6344
rect 114005 6307 114063 6313
rect 114005 6273 114017 6307
rect 114051 6273 114063 6307
rect 114005 6267 114063 6273
rect 114189 6307 114247 6313
rect 114189 6273 114201 6307
rect 114235 6304 114247 6307
rect 114554 6304 114560 6316
rect 114235 6276 114560 6304
rect 114235 6273 114247 6276
rect 114189 6267 114247 6273
rect 108408 6208 109034 6236
rect 90913 6171 90971 6177
rect 90913 6137 90925 6171
rect 90959 6168 90971 6171
rect 98457 6171 98515 6177
rect 90959 6140 97120 6168
rect 90959 6137 90971 6140
rect 90913 6131 90971 6137
rect 85632 6072 87644 6100
rect 92293 6103 92351 6109
rect 85632 6060 85638 6072
rect 92293 6069 92305 6103
rect 92339 6100 92351 6103
rect 93118 6100 93124 6112
rect 92339 6072 93124 6100
rect 92339 6069 92351 6072
rect 92293 6063 92351 6069
rect 93118 6060 93124 6072
rect 93176 6060 93182 6112
rect 93854 6060 93860 6112
rect 93912 6100 93918 6112
rect 94314 6100 94320 6112
rect 93912 6072 94320 6100
rect 93912 6060 93918 6072
rect 94314 6060 94320 6072
rect 94372 6060 94378 6112
rect 96614 6100 96620 6112
rect 96575 6072 96620 6100
rect 96614 6060 96620 6072
rect 96672 6060 96678 6112
rect 97092 6100 97120 6140
rect 98457 6137 98469 6171
rect 98503 6137 98515 6171
rect 105078 6168 105084 6180
rect 98457 6131 98515 6137
rect 99346 6140 105084 6168
rect 99346 6100 99374 6140
rect 105078 6128 105084 6140
rect 105136 6128 105142 6180
rect 97092 6072 99374 6100
rect 100938 6060 100944 6112
rect 100996 6100 101002 6112
rect 108408 6100 108436 6208
rect 114020 6168 114048 6267
rect 114554 6264 114560 6276
rect 114612 6304 114618 6316
rect 114922 6304 114928 6316
rect 114612 6276 114928 6304
rect 114612 6264 114618 6276
rect 114922 6264 114928 6276
rect 114980 6264 114986 6316
rect 115842 6264 115848 6316
rect 115900 6313 115906 6316
rect 115900 6304 115912 6313
rect 116044 6304 116072 6344
rect 119062 6332 119068 6384
rect 119120 6372 119126 6384
rect 119249 6375 119307 6381
rect 119249 6372 119261 6375
rect 119120 6344 119261 6372
rect 119120 6332 119126 6344
rect 119249 6341 119261 6344
rect 119295 6341 119307 6375
rect 121748 6372 121776 6403
rect 121914 6400 121920 6452
rect 121972 6440 121978 6452
rect 121972 6412 123239 6440
rect 121972 6400 121978 6412
rect 119249 6335 119307 6341
rect 120184 6344 121776 6372
rect 120184 6304 120212 6344
rect 121822 6332 121828 6384
rect 121880 6372 121886 6384
rect 122742 6372 122748 6384
rect 121880 6344 122748 6372
rect 121880 6332 121886 6344
rect 122742 6332 122748 6344
rect 122800 6372 122806 6384
rect 123211 6372 123239 6412
rect 123846 6400 123852 6452
rect 123904 6440 123910 6452
rect 126146 6440 126152 6452
rect 123904 6412 126152 6440
rect 123904 6400 123910 6412
rect 126146 6400 126152 6412
rect 126204 6400 126210 6452
rect 126698 6400 126704 6452
rect 126756 6440 126762 6452
rect 126885 6443 126943 6449
rect 126885 6440 126897 6443
rect 126756 6412 126897 6440
rect 126756 6400 126762 6412
rect 126885 6409 126897 6412
rect 126931 6409 126943 6443
rect 127986 6440 127992 6452
rect 126885 6403 126943 6409
rect 126992 6412 127992 6440
rect 126992 6372 127020 6412
rect 127986 6400 127992 6412
rect 128044 6400 128050 6452
rect 128538 6400 128544 6452
rect 128596 6440 128602 6452
rect 129550 6440 129556 6452
rect 128596 6412 128952 6440
rect 129511 6412 129556 6440
rect 128596 6400 128602 6412
rect 128262 6372 128268 6384
rect 122800 6344 123156 6372
rect 123211 6344 127020 6372
rect 127360 6344 128268 6372
rect 122800 6332 122806 6344
rect 115900 6276 115945 6304
rect 116044 6276 120212 6304
rect 121017 6307 121075 6313
rect 115900 6267 115912 6276
rect 121017 6273 121029 6307
rect 121063 6304 121075 6307
rect 122558 6304 122564 6316
rect 121063 6276 122564 6304
rect 121063 6273 121075 6276
rect 121017 6267 121075 6273
rect 115900 6264 115906 6267
rect 122558 6264 122564 6276
rect 122616 6264 122622 6316
rect 123128 6313 123156 6344
rect 122857 6307 122915 6313
rect 122857 6273 122869 6307
rect 122903 6304 122915 6307
rect 123113 6307 123171 6313
rect 122903 6276 123064 6304
rect 122903 6273 122915 6276
rect 122857 6267 122915 6273
rect 116118 6236 116124 6248
rect 116079 6208 116124 6236
rect 116118 6196 116124 6208
rect 116176 6196 116182 6248
rect 116673 6239 116731 6245
rect 116673 6205 116685 6239
rect 116719 6236 116731 6239
rect 119890 6236 119896 6248
rect 116719 6208 119896 6236
rect 116719 6205 116731 6208
rect 116673 6199 116731 6205
rect 113284 6140 114048 6168
rect 100996 6072 108436 6100
rect 100996 6060 101002 6072
rect 111886 6060 111892 6112
rect 111944 6100 111950 6112
rect 113284 6109 113312 6140
rect 114646 6128 114652 6180
rect 114704 6168 114710 6180
rect 114741 6171 114799 6177
rect 114741 6168 114753 6171
rect 114704 6140 114753 6168
rect 114704 6128 114710 6140
rect 114741 6137 114753 6140
rect 114787 6137 114799 6171
rect 114741 6131 114799 6137
rect 113269 6103 113327 6109
rect 113269 6100 113281 6103
rect 111944 6072 113281 6100
rect 111944 6060 111950 6072
rect 113269 6069 113281 6072
rect 113315 6069 113327 6103
rect 113818 6100 113824 6112
rect 113779 6072 113824 6100
rect 113269 6063 113327 6069
rect 113818 6060 113824 6072
rect 113876 6060 113882 6112
rect 115842 6060 115848 6112
rect 115900 6100 115906 6112
rect 116688 6100 116716 6199
rect 119890 6196 119896 6208
rect 119948 6196 119954 6248
rect 121273 6239 121331 6245
rect 121273 6205 121285 6239
rect 121319 6236 121331 6239
rect 121822 6236 121828 6248
rect 121319 6208 121828 6236
rect 121319 6205 121331 6208
rect 121273 6199 121331 6205
rect 121822 6196 121828 6208
rect 121880 6196 121886 6248
rect 123036 6236 123064 6276
rect 123113 6273 123125 6307
rect 123159 6304 123171 6307
rect 124858 6304 124864 6316
rect 123159 6276 124864 6304
rect 123159 6273 123171 6276
rect 123113 6267 123171 6273
rect 124858 6264 124864 6276
rect 124916 6304 124922 6316
rect 125226 6304 125232 6316
rect 124916 6276 125232 6304
rect 124916 6264 124922 6276
rect 125226 6264 125232 6276
rect 125284 6304 125290 6316
rect 127360 6313 127388 6344
rect 128262 6332 128268 6344
rect 128320 6332 128326 6384
rect 128924 6372 128952 6412
rect 129550 6400 129556 6412
rect 129608 6400 129614 6452
rect 130194 6440 130200 6452
rect 130155 6412 130200 6440
rect 130194 6400 130200 6412
rect 130252 6440 130258 6452
rect 135070 6440 135076 6452
rect 130252 6412 134104 6440
rect 130252 6400 130258 6412
rect 129001 6375 129059 6381
rect 129001 6372 129013 6375
rect 128924 6344 129013 6372
rect 129001 6341 129013 6344
rect 129047 6341 129059 6375
rect 129001 6335 129059 6341
rect 130562 6332 130568 6384
rect 130620 6372 130626 6384
rect 131574 6372 131580 6384
rect 130620 6344 131580 6372
rect 130620 6332 130626 6344
rect 131574 6332 131580 6344
rect 131632 6332 131638 6384
rect 125505 6307 125563 6313
rect 125505 6304 125517 6307
rect 125284 6276 125517 6304
rect 125284 6264 125290 6276
rect 125505 6273 125517 6276
rect 125551 6273 125563 6307
rect 125505 6267 125563 6273
rect 125772 6307 125830 6313
rect 125772 6273 125784 6307
rect 125818 6304 125830 6307
rect 127345 6307 127403 6313
rect 127345 6304 127357 6307
rect 125818 6276 127357 6304
rect 125818 6273 125830 6276
rect 125772 6267 125830 6273
rect 127345 6273 127357 6276
rect 127391 6273 127403 6307
rect 127345 6267 127403 6273
rect 123294 6236 123300 6248
rect 123036 6208 123300 6236
rect 123294 6196 123300 6208
rect 123352 6236 123358 6248
rect 123938 6236 123944 6248
rect 123352 6208 123944 6236
rect 123352 6196 123358 6208
rect 123938 6196 123944 6208
rect 123996 6196 124002 6248
rect 116762 6128 116768 6180
rect 116820 6168 116826 6180
rect 116820 6140 120396 6168
rect 116820 6128 116826 6140
rect 118234 6100 118240 6112
rect 115900 6072 116716 6100
rect 118195 6072 118240 6100
rect 115900 6060 115906 6072
rect 118234 6060 118240 6072
rect 118292 6060 118298 6112
rect 118789 6103 118847 6109
rect 118789 6069 118801 6103
rect 118835 6100 118847 6103
rect 119706 6100 119712 6112
rect 118835 6072 119712 6100
rect 118835 6069 118847 6072
rect 118789 6063 118847 6069
rect 119706 6060 119712 6072
rect 119764 6060 119770 6112
rect 120368 6100 120396 6140
rect 123110 6128 123116 6180
rect 123168 6168 123174 6180
rect 123665 6171 123723 6177
rect 123665 6168 123677 6171
rect 123168 6140 123677 6168
rect 123168 6128 123174 6140
rect 123665 6137 123677 6140
rect 123711 6168 123723 6171
rect 123846 6168 123852 6180
rect 123711 6140 123852 6168
rect 123711 6137 123723 6140
rect 123665 6131 123723 6137
rect 123846 6128 123852 6140
rect 123904 6128 123910 6180
rect 124398 6168 124404 6180
rect 124359 6140 124404 6168
rect 124398 6128 124404 6140
rect 124456 6128 124462 6180
rect 124214 6100 124220 6112
rect 120368 6072 124220 6100
rect 124214 6060 124220 6072
rect 124272 6060 124278 6112
rect 125520 6100 125548 6267
rect 127526 6264 127532 6316
rect 127584 6304 127590 6316
rect 129274 6304 129280 6316
rect 127584 6276 129280 6304
rect 127584 6264 127590 6276
rect 129274 6264 129280 6276
rect 129332 6264 129338 6316
rect 129366 6264 129372 6316
rect 129424 6304 129430 6316
rect 134076 6304 134104 6412
rect 134260 6412 135076 6440
rect 134260 6384 134288 6412
rect 135070 6400 135076 6412
rect 135128 6400 135134 6452
rect 136910 6400 136916 6452
rect 136968 6440 136974 6452
rect 137649 6443 137707 6449
rect 137649 6440 137661 6443
rect 136968 6412 137661 6440
rect 136968 6400 136974 6412
rect 137649 6409 137661 6412
rect 137695 6409 137707 6443
rect 139670 6440 139676 6452
rect 137649 6403 137707 6409
rect 138768 6412 139676 6440
rect 134242 6372 134248 6384
rect 134203 6344 134248 6372
rect 134242 6332 134248 6344
rect 134300 6332 134306 6384
rect 134797 6375 134855 6381
rect 134797 6341 134809 6375
rect 134843 6372 134855 6375
rect 135898 6372 135904 6384
rect 134843 6344 135904 6372
rect 134843 6341 134855 6344
rect 134797 6335 134855 6341
rect 135898 6332 135904 6344
rect 135956 6372 135962 6384
rect 138198 6372 138204 6384
rect 135956 6344 138204 6372
rect 135956 6332 135962 6344
rect 138198 6332 138204 6344
rect 138256 6332 138262 6384
rect 138658 6304 138664 6316
rect 129424 6276 133716 6304
rect 134076 6276 138664 6304
rect 129424 6264 129430 6276
rect 127989 6239 128047 6245
rect 127989 6205 128001 6239
rect 128035 6236 128047 6239
rect 128078 6236 128084 6248
rect 128035 6208 128084 6236
rect 128035 6205 128047 6208
rect 127989 6199 128047 6205
rect 128078 6196 128084 6208
rect 128136 6196 128142 6248
rect 128262 6196 128268 6248
rect 128320 6236 128326 6248
rect 130838 6236 130844 6248
rect 128320 6208 130844 6236
rect 128320 6196 128326 6208
rect 130838 6196 130844 6208
rect 130896 6196 130902 6248
rect 130933 6239 130991 6245
rect 130933 6205 130945 6239
rect 130979 6236 130991 6239
rect 132218 6236 132224 6248
rect 130979 6208 132224 6236
rect 130979 6205 130991 6208
rect 130933 6199 130991 6205
rect 126514 6128 126520 6180
rect 126572 6168 126578 6180
rect 130948 6168 130976 6199
rect 132218 6196 132224 6208
rect 132276 6196 132282 6248
rect 132589 6239 132647 6245
rect 132589 6205 132601 6239
rect 132635 6236 132647 6239
rect 132770 6236 132776 6248
rect 132635 6208 132776 6236
rect 132635 6205 132647 6208
rect 132589 6199 132647 6205
rect 132770 6196 132776 6208
rect 132828 6236 132834 6248
rect 132954 6236 132960 6248
rect 132828 6208 132960 6236
rect 132828 6196 132834 6208
rect 132954 6196 132960 6208
rect 133012 6196 133018 6248
rect 133046 6196 133052 6248
rect 133104 6236 133110 6248
rect 133601 6239 133659 6245
rect 133601 6236 133613 6239
rect 133104 6208 133613 6236
rect 133104 6196 133110 6208
rect 133601 6205 133613 6208
rect 133647 6205 133659 6239
rect 133688 6236 133716 6276
rect 138658 6264 138664 6276
rect 138716 6264 138722 6316
rect 138768 6236 138796 6412
rect 139670 6400 139676 6412
rect 139728 6400 139734 6452
rect 139854 6400 139860 6452
rect 139912 6440 139918 6452
rect 143350 6440 143356 6452
rect 139912 6412 143356 6440
rect 139912 6400 139918 6412
rect 143350 6400 143356 6412
rect 143408 6400 143414 6452
rect 143902 6400 143908 6452
rect 143960 6440 143966 6452
rect 145006 6440 145012 6452
rect 143960 6412 145012 6440
rect 143960 6400 143966 6412
rect 145006 6400 145012 6412
rect 145064 6400 145070 6452
rect 145650 6440 145656 6452
rect 145611 6412 145656 6440
rect 145650 6400 145656 6412
rect 145708 6400 145714 6452
rect 146294 6400 146300 6452
rect 146352 6440 146358 6452
rect 147582 6440 147588 6452
rect 146352 6412 147588 6440
rect 146352 6400 146358 6412
rect 147582 6400 147588 6412
rect 147640 6400 147646 6452
rect 148226 6400 148232 6452
rect 148284 6440 148290 6452
rect 148873 6443 148931 6449
rect 148873 6440 148885 6443
rect 148284 6412 148885 6440
rect 148284 6400 148290 6412
rect 148873 6409 148885 6412
rect 148919 6409 148931 6443
rect 148873 6403 148931 6409
rect 149146 6400 149152 6452
rect 149204 6440 149210 6452
rect 149790 6440 149796 6452
rect 149204 6412 149796 6440
rect 149204 6400 149210 6412
rect 149790 6400 149796 6412
rect 149848 6400 149854 6452
rect 149882 6400 149888 6452
rect 149940 6440 149946 6452
rect 150069 6443 150127 6449
rect 150069 6440 150081 6443
rect 149940 6412 150081 6440
rect 149940 6400 149946 6412
rect 150069 6409 150081 6412
rect 150115 6409 150127 6443
rect 150069 6403 150127 6409
rect 150434 6400 150440 6452
rect 150492 6440 150498 6452
rect 152645 6443 152703 6449
rect 152645 6440 152657 6443
rect 150492 6412 152657 6440
rect 150492 6400 150498 6412
rect 152645 6409 152657 6412
rect 152691 6409 152703 6443
rect 152645 6403 152703 6409
rect 152918 6400 152924 6452
rect 152976 6440 152982 6452
rect 157429 6443 157487 6449
rect 157429 6440 157441 6443
rect 152976 6412 157441 6440
rect 152976 6400 152982 6412
rect 157429 6409 157441 6412
rect 157475 6409 157487 6443
rect 157429 6403 157487 6409
rect 138845 6375 138903 6381
rect 138845 6341 138857 6375
rect 138891 6372 138903 6375
rect 141234 6372 141240 6384
rect 138891 6344 141240 6372
rect 138891 6341 138903 6344
rect 138845 6335 138903 6341
rect 133688 6208 138796 6236
rect 133601 6199 133659 6205
rect 126572 6140 130976 6168
rect 126572 6128 126578 6140
rect 131574 6128 131580 6180
rect 131632 6168 131638 6180
rect 138860 6168 138888 6335
rect 141234 6332 141240 6344
rect 141292 6332 141298 6384
rect 141326 6332 141332 6384
rect 141384 6372 141390 6384
rect 143718 6372 143724 6384
rect 141384 6344 143724 6372
rect 141384 6332 141390 6344
rect 143718 6332 143724 6344
rect 143776 6332 143782 6384
rect 143810 6332 143816 6384
rect 143868 6372 143874 6384
rect 147738 6375 147796 6381
rect 147738 6372 147750 6375
rect 143868 6344 147750 6372
rect 143868 6332 143874 6344
rect 147738 6341 147750 6344
rect 147784 6341 147796 6375
rect 147738 6335 147796 6341
rect 147858 6332 147864 6384
rect 147916 6372 147922 6384
rect 155129 6375 155187 6381
rect 147916 6344 155080 6372
rect 147916 6332 147922 6344
rect 142798 6304 142804 6316
rect 142759 6276 142804 6304
rect 142798 6264 142804 6276
rect 142856 6264 142862 6316
rect 142890 6264 142896 6316
rect 142948 6304 142954 6316
rect 144086 6304 144092 6316
rect 142948 6276 144092 6304
rect 142948 6264 142954 6276
rect 144086 6264 144092 6276
rect 144144 6264 144150 6316
rect 144569 6307 144627 6313
rect 144569 6273 144581 6307
rect 144615 6304 144627 6307
rect 144730 6304 144736 6316
rect 144615 6276 144736 6304
rect 144615 6273 144627 6276
rect 144569 6267 144627 6273
rect 144730 6264 144736 6276
rect 144788 6264 144794 6316
rect 144825 6307 144883 6313
rect 144825 6273 144837 6307
rect 144871 6304 144883 6307
rect 144914 6304 144920 6316
rect 144871 6276 144920 6304
rect 144871 6273 144883 6276
rect 144825 6267 144883 6273
rect 144914 6264 144920 6276
rect 144972 6304 144978 6316
rect 145650 6304 145656 6316
rect 144972 6276 145656 6304
rect 144972 6264 144978 6276
rect 145650 6264 145656 6276
rect 145708 6264 145714 6316
rect 145926 6264 145932 6316
rect 145984 6304 145990 6316
rect 146777 6307 146835 6313
rect 146777 6304 146789 6307
rect 145984 6276 146789 6304
rect 145984 6264 145990 6276
rect 146777 6273 146789 6276
rect 146823 6304 146835 6307
rect 146938 6304 146944 6316
rect 146823 6276 146944 6304
rect 146823 6273 146835 6276
rect 146777 6267 146835 6273
rect 146938 6264 146944 6276
rect 146996 6264 147002 6316
rect 147122 6264 147128 6316
rect 147180 6304 147186 6316
rect 149146 6304 149152 6316
rect 147180 6276 149152 6304
rect 147180 6264 147186 6276
rect 149146 6264 149152 6276
rect 149204 6264 149210 6316
rect 149330 6304 149336 6316
rect 149291 6276 149336 6304
rect 149330 6264 149336 6276
rect 149388 6264 149394 6316
rect 150250 6304 150256 6316
rect 150211 6276 150256 6304
rect 150250 6264 150256 6276
rect 150308 6264 150314 6316
rect 150989 6307 151047 6313
rect 150989 6273 151001 6307
rect 151035 6304 151047 6307
rect 151078 6304 151084 6316
rect 151035 6276 151084 6304
rect 151035 6273 151047 6276
rect 150989 6267 151047 6273
rect 151078 6264 151084 6276
rect 151136 6264 151142 6316
rect 151817 6307 151875 6313
rect 151817 6273 151829 6307
rect 151863 6304 151875 6307
rect 152366 6304 152372 6316
rect 151863 6276 152372 6304
rect 151863 6273 151875 6276
rect 151817 6267 151875 6273
rect 152366 6264 152372 6276
rect 152424 6264 152430 6316
rect 152829 6307 152887 6313
rect 152829 6273 152841 6307
rect 152875 6304 152887 6307
rect 153378 6304 153384 6316
rect 152875 6276 153384 6304
rect 152875 6273 152887 6276
rect 152829 6267 152887 6273
rect 153378 6264 153384 6276
rect 153436 6264 153442 6316
rect 153657 6307 153715 6313
rect 153657 6273 153669 6307
rect 153703 6304 153715 6307
rect 153746 6304 153752 6316
rect 153703 6276 153752 6304
rect 153703 6273 153715 6276
rect 153657 6267 153715 6273
rect 153746 6264 153752 6276
rect 153804 6264 153810 6316
rect 154022 6264 154028 6316
rect 154080 6304 154086 6316
rect 154482 6304 154488 6316
rect 154080 6276 154488 6304
rect 154080 6264 154086 6276
rect 154482 6264 154488 6276
rect 154540 6264 154546 6316
rect 154853 6307 154911 6313
rect 154853 6273 154865 6307
rect 154899 6273 154911 6307
rect 154853 6267 154911 6273
rect 154945 6307 155003 6313
rect 154945 6273 154957 6307
rect 154991 6273 155003 6307
rect 155052 6304 155080 6344
rect 155129 6341 155141 6375
rect 155175 6372 155187 6375
rect 157794 6372 157800 6384
rect 155175 6344 157800 6372
rect 155175 6341 155187 6344
rect 155129 6335 155187 6341
rect 157794 6332 157800 6344
rect 157852 6332 157858 6384
rect 158438 6372 158444 6384
rect 158088 6344 158444 6372
rect 156141 6307 156199 6313
rect 156141 6304 156153 6307
rect 155052 6276 156153 6304
rect 154945 6267 155003 6273
rect 156141 6273 156153 6276
rect 156187 6273 156199 6307
rect 156141 6267 156199 6273
rect 139670 6196 139676 6248
rect 139728 6236 139734 6248
rect 140501 6239 140559 6245
rect 140501 6236 140513 6239
rect 139728 6208 140513 6236
rect 139728 6196 139734 6208
rect 140501 6205 140513 6208
rect 140547 6236 140559 6239
rect 140682 6236 140688 6248
rect 140547 6208 140688 6236
rect 140547 6205 140559 6208
rect 140501 6199 140559 6205
rect 140682 6196 140688 6208
rect 140740 6196 140746 6248
rect 147030 6236 147036 6248
rect 143368 6208 143663 6236
rect 146991 6208 147036 6236
rect 131632 6140 138888 6168
rect 131632 6128 131638 6140
rect 138934 6128 138940 6180
rect 138992 6168 138998 6180
rect 143368 6168 143396 6208
rect 138992 6140 143396 6168
rect 138992 6128 138998 6140
rect 127618 6100 127624 6112
rect 125520 6072 127624 6100
rect 127618 6060 127624 6072
rect 127676 6060 127682 6112
rect 128538 6100 128544 6112
rect 128499 6072 128544 6100
rect 128538 6060 128544 6072
rect 128596 6060 128602 6112
rect 128722 6060 128728 6112
rect 128780 6100 128786 6112
rect 131206 6100 131212 6112
rect 128780 6072 131212 6100
rect 128780 6060 128786 6072
rect 131206 6060 131212 6072
rect 131264 6060 131270 6112
rect 131482 6100 131488 6112
rect 131443 6072 131488 6100
rect 131482 6060 131488 6072
rect 131540 6060 131546 6112
rect 132037 6103 132095 6109
rect 132037 6069 132049 6103
rect 132083 6100 132095 6103
rect 132310 6100 132316 6112
rect 132083 6072 132316 6100
rect 132083 6069 132095 6072
rect 132037 6063 132095 6069
rect 132310 6060 132316 6072
rect 132368 6060 132374 6112
rect 132954 6060 132960 6112
rect 133012 6100 133018 6112
rect 133049 6103 133107 6109
rect 133049 6100 133061 6103
rect 133012 6072 133061 6100
rect 133012 6060 133018 6072
rect 133049 6069 133061 6072
rect 133095 6100 133107 6103
rect 135254 6100 135260 6112
rect 133095 6072 135260 6100
rect 133095 6069 133107 6072
rect 133049 6063 133107 6069
rect 135254 6060 135260 6072
rect 135312 6060 135318 6112
rect 135809 6103 135867 6109
rect 135809 6069 135821 6103
rect 135855 6100 135867 6103
rect 136082 6100 136088 6112
rect 135855 6072 136088 6100
rect 135855 6069 135867 6072
rect 135809 6063 135867 6069
rect 136082 6060 136088 6072
rect 136140 6060 136146 6112
rect 136361 6103 136419 6109
rect 136361 6069 136373 6103
rect 136407 6100 136419 6103
rect 136634 6100 136640 6112
rect 136407 6072 136640 6100
rect 136407 6069 136419 6072
rect 136361 6063 136419 6069
rect 136634 6060 136640 6072
rect 136692 6100 136698 6112
rect 136821 6103 136879 6109
rect 136821 6100 136833 6103
rect 136692 6072 136833 6100
rect 136692 6060 136698 6072
rect 136821 6069 136833 6072
rect 136867 6100 136879 6103
rect 137922 6100 137928 6112
rect 136867 6072 137928 6100
rect 136867 6069 136879 6072
rect 136821 6063 136879 6069
rect 137922 6060 137928 6072
rect 137980 6100 137986 6112
rect 138201 6103 138259 6109
rect 138201 6100 138213 6103
rect 137980 6072 138213 6100
rect 137980 6060 137986 6072
rect 138201 6069 138213 6072
rect 138247 6069 138259 6103
rect 138201 6063 138259 6069
rect 139397 6103 139455 6109
rect 139397 6069 139409 6103
rect 139443 6100 139455 6103
rect 139854 6100 139860 6112
rect 139443 6072 139860 6100
rect 139443 6069 139455 6072
rect 139397 6063 139455 6069
rect 139854 6060 139860 6072
rect 139912 6060 139918 6112
rect 139949 6103 140007 6109
rect 139949 6069 139961 6103
rect 139995 6100 140007 6103
rect 140038 6100 140044 6112
rect 139995 6072 140044 6100
rect 139995 6069 140007 6072
rect 139949 6063 140007 6069
rect 140038 6060 140044 6072
rect 140096 6100 140102 6112
rect 140406 6100 140412 6112
rect 140096 6072 140412 6100
rect 140096 6060 140102 6072
rect 140406 6060 140412 6072
rect 140464 6060 140470 6112
rect 140590 6060 140596 6112
rect 140648 6100 140654 6112
rect 143445 6103 143503 6109
rect 143445 6100 143457 6103
rect 140648 6072 143457 6100
rect 140648 6060 140654 6072
rect 143445 6069 143457 6072
rect 143491 6069 143503 6103
rect 143635 6100 143663 6208
rect 147030 6196 147036 6208
rect 147088 6196 147094 6248
rect 147493 6239 147551 6245
rect 147493 6205 147505 6239
rect 147539 6205 147551 6239
rect 147493 6199 147551 6205
rect 145926 6168 145932 6180
rect 144886 6140 145932 6168
rect 144886 6100 144914 6140
rect 145926 6128 145932 6140
rect 145984 6128 145990 6180
rect 143635 6072 144914 6100
rect 143445 6063 143503 6069
rect 146386 6060 146392 6112
rect 146444 6100 146450 6112
rect 147398 6100 147404 6112
rect 146444 6072 147404 6100
rect 146444 6060 146450 6072
rect 147398 6060 147404 6072
rect 147456 6100 147462 6112
rect 147508 6100 147536 6199
rect 148502 6196 148508 6248
rect 148560 6236 148566 6248
rect 152918 6236 152924 6248
rect 148560 6208 152924 6236
rect 148560 6196 148566 6208
rect 152918 6196 152924 6208
rect 152976 6196 152982 6248
rect 153470 6196 153476 6248
rect 153528 6236 153534 6248
rect 153528 6208 154068 6236
rect 153528 6196 153534 6208
rect 148778 6128 148784 6180
rect 148836 6168 148842 6180
rect 150066 6168 150072 6180
rect 148836 6140 150072 6168
rect 148836 6128 148842 6140
rect 150066 6128 150072 6140
rect 150124 6128 150130 6180
rect 151630 6168 151636 6180
rect 150176 6140 151492 6168
rect 151591 6140 151636 6168
rect 147456 6072 147536 6100
rect 147456 6060 147462 6072
rect 147766 6060 147772 6112
rect 147824 6100 147830 6112
rect 149238 6100 149244 6112
rect 147824 6072 149244 6100
rect 147824 6060 147830 6072
rect 149238 6060 149244 6072
rect 149296 6060 149302 6112
rect 149514 6100 149520 6112
rect 149475 6072 149520 6100
rect 149514 6060 149520 6072
rect 149572 6100 149578 6112
rect 150176 6100 150204 6140
rect 149572 6072 150204 6100
rect 149572 6060 149578 6072
rect 150250 6060 150256 6112
rect 150308 6100 150314 6112
rect 150805 6103 150863 6109
rect 150805 6100 150817 6103
rect 150308 6072 150817 6100
rect 150308 6060 150314 6072
rect 150805 6069 150817 6072
rect 150851 6069 150863 6103
rect 151464 6100 151492 6140
rect 151630 6128 151636 6140
rect 151688 6128 151694 6180
rect 153930 6168 153936 6180
rect 151740 6140 153936 6168
rect 151740 6100 151768 6140
rect 153930 6128 153936 6140
rect 153988 6128 153994 6180
rect 154040 6168 154068 6208
rect 154868 6168 154896 6267
rect 154040 6140 154896 6168
rect 154960 6168 154988 6267
rect 156414 6264 156420 6316
rect 156472 6304 156478 6316
rect 156969 6307 157027 6313
rect 156969 6304 156981 6307
rect 156472 6276 156981 6304
rect 156472 6264 156478 6276
rect 156969 6273 156981 6276
rect 157015 6273 157027 6307
rect 156969 6267 157027 6273
rect 157613 6307 157671 6313
rect 157613 6273 157625 6307
rect 157659 6304 157671 6307
rect 158088 6304 158116 6344
rect 158438 6332 158444 6344
rect 158496 6332 158502 6384
rect 157659 6276 158116 6304
rect 157659 6273 157671 6276
rect 157613 6267 157671 6273
rect 158162 6264 158168 6316
rect 158220 6304 158226 6316
rect 158257 6307 158315 6313
rect 158257 6304 158269 6307
rect 158220 6276 158269 6304
rect 158220 6264 158226 6276
rect 158257 6273 158269 6276
rect 158303 6273 158315 6307
rect 158257 6267 158315 6273
rect 155218 6196 155224 6248
rect 155276 6236 155282 6248
rect 155957 6239 156015 6245
rect 155957 6236 155969 6239
rect 155276 6208 155969 6236
rect 155276 6196 155282 6208
rect 155957 6205 155969 6208
rect 156003 6236 156015 6239
rect 156782 6236 156788 6248
rect 156003 6208 156788 6236
rect 156003 6205 156015 6208
rect 155957 6199 156015 6205
rect 156782 6196 156788 6208
rect 156840 6196 156846 6248
rect 155310 6168 155316 6180
rect 154960 6140 155316 6168
rect 155310 6128 155316 6140
rect 155368 6128 155374 6180
rect 151464 6072 151768 6100
rect 150805 6063 150863 6069
rect 152642 6060 152648 6112
rect 152700 6100 152706 6112
rect 153654 6100 153660 6112
rect 152700 6072 153660 6100
rect 152700 6060 152706 6072
rect 153654 6060 153660 6072
rect 153712 6100 153718 6112
rect 153749 6103 153807 6109
rect 153749 6100 153761 6103
rect 153712 6072 153761 6100
rect 153712 6060 153718 6072
rect 153749 6069 153761 6072
rect 153795 6069 153807 6103
rect 153749 6063 153807 6069
rect 154298 6060 154304 6112
rect 154356 6100 154362 6112
rect 155862 6100 155868 6112
rect 154356 6072 155868 6100
rect 154356 6060 154362 6072
rect 155862 6060 155868 6072
rect 155920 6060 155926 6112
rect 156322 6100 156328 6112
rect 156283 6072 156328 6100
rect 156322 6060 156328 6072
rect 156380 6060 156386 6112
rect 156782 6100 156788 6112
rect 156743 6072 156788 6100
rect 156782 6060 156788 6072
rect 156840 6060 156846 6112
rect 157058 6060 157064 6112
rect 157116 6100 157122 6112
rect 158073 6103 158131 6109
rect 158073 6100 158085 6103
rect 157116 6072 158085 6100
rect 157116 6060 157122 6072
rect 158073 6069 158085 6072
rect 158119 6069 158131 6103
rect 158073 6063 158131 6069
rect 1104 6010 158884 6032
rect 1104 5958 20672 6010
rect 20724 5958 20736 6010
rect 20788 5958 20800 6010
rect 20852 5958 20864 6010
rect 20916 5958 20928 6010
rect 20980 5958 60117 6010
rect 60169 5958 60181 6010
rect 60233 5958 60245 6010
rect 60297 5958 60309 6010
rect 60361 5958 60373 6010
rect 60425 5958 99562 6010
rect 99614 5958 99626 6010
rect 99678 5958 99690 6010
rect 99742 5958 99754 6010
rect 99806 5958 99818 6010
rect 99870 5958 139007 6010
rect 139059 5958 139071 6010
rect 139123 5958 139135 6010
rect 139187 5958 139199 6010
rect 139251 5958 139263 6010
rect 139315 5958 158884 6010
rect 1104 5936 158884 5958
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 4948 5868 5365 5896
rect 4948 5856 4954 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5776 5868 5825 5896
rect 5776 5856 5782 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15252 5868 16129 5896
rect 15252 5856 15258 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 16574 5856 16580 5908
rect 16632 5896 16638 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 16632 5868 16957 5896
rect 16632 5856 16638 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 18138 5896 18144 5908
rect 16945 5859 17003 5865
rect 17328 5868 18144 5896
rect 17328 5840 17356 5868
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 18874 5896 18880 5908
rect 18371 5868 18880 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19576 5868 19625 5896
rect 19576 5856 19582 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 21821 5899 21879 5905
rect 21821 5896 21833 5899
rect 20404 5868 21833 5896
rect 20404 5856 20410 5868
rect 21821 5865 21833 5868
rect 21867 5896 21879 5899
rect 22002 5896 22008 5908
rect 21867 5868 22008 5896
rect 21867 5865 21879 5868
rect 21821 5859 21879 5865
rect 22002 5856 22008 5868
rect 22060 5856 22066 5908
rect 22462 5856 22468 5908
rect 22520 5896 22526 5908
rect 24026 5896 24032 5908
rect 22520 5868 24032 5896
rect 22520 5856 22526 5868
rect 24026 5856 24032 5868
rect 24084 5856 24090 5908
rect 24765 5899 24823 5905
rect 24765 5865 24777 5899
rect 24811 5896 24823 5899
rect 24854 5896 24860 5908
rect 24811 5868 24860 5896
rect 24811 5865 24823 5868
rect 24765 5859 24823 5865
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 28902 5856 28908 5908
rect 28960 5896 28966 5908
rect 30009 5899 30067 5905
rect 30009 5896 30021 5899
rect 28960 5868 30021 5896
rect 28960 5856 28966 5868
rect 30009 5865 30021 5868
rect 30055 5865 30067 5899
rect 30009 5859 30067 5865
rect 30374 5856 30380 5908
rect 30432 5896 30438 5908
rect 32306 5896 32312 5908
rect 30432 5868 32168 5896
rect 32219 5868 32312 5896
rect 30432 5856 30438 5868
rect 17310 5828 17316 5840
rect 16500 5800 17316 5828
rect 16500 5769 16528 5800
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 17494 5788 17500 5840
rect 17552 5828 17558 5840
rect 30466 5828 30472 5840
rect 17552 5800 30472 5828
rect 17552 5788 17558 5800
rect 30466 5788 30472 5800
rect 30524 5788 30530 5840
rect 30558 5788 30564 5840
rect 30616 5828 30622 5840
rect 32030 5828 32036 5840
rect 30616 5800 32036 5828
rect 30616 5788 30622 5800
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 32140 5828 32168 5868
rect 32306 5856 32312 5868
rect 32364 5896 32370 5908
rect 33778 5896 33784 5908
rect 32364 5868 33784 5896
rect 32364 5856 32370 5868
rect 33778 5856 33784 5868
rect 33836 5856 33842 5908
rect 38013 5899 38071 5905
rect 33888 5868 37412 5896
rect 33888 5828 33916 5868
rect 32140 5800 33916 5828
rect 33962 5788 33968 5840
rect 34020 5828 34026 5840
rect 35989 5831 36047 5837
rect 35989 5828 36001 5831
rect 34020 5800 36001 5828
rect 34020 5788 34026 5800
rect 35989 5797 36001 5800
rect 36035 5797 36047 5831
rect 35989 5791 36047 5797
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 20254 5760 20260 5772
rect 16485 5723 16543 5729
rect 17144 5732 20260 5760
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4240 5695 4298 5701
rect 4240 5661 4252 5695
rect 4286 5692 4298 5695
rect 4614 5692 4620 5704
rect 4286 5664 4620 5692
rect 4286 5661 4298 5664
rect 4240 5655 4298 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6086 5692 6092 5704
rect 6043 5664 6092 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 14274 5692 14280 5704
rect 13771 5664 14280 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 13188 5624 13216 5655
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 17144 5701 17172 5732
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 25222 5760 25228 5772
rect 22060 5732 25228 5760
rect 22060 5720 22066 5732
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 25774 5720 25780 5772
rect 25832 5760 25838 5772
rect 35437 5763 35495 5769
rect 35437 5760 35449 5763
rect 25832 5732 35449 5760
rect 25832 5720 25838 5732
rect 35437 5729 35449 5732
rect 35483 5760 35495 5763
rect 37384 5760 37412 5868
rect 38013 5865 38025 5899
rect 38059 5896 38071 5899
rect 38654 5896 38660 5908
rect 38059 5868 38660 5896
rect 38059 5865 38071 5868
rect 38013 5859 38071 5865
rect 38654 5856 38660 5868
rect 38712 5856 38718 5908
rect 43254 5896 43260 5908
rect 43215 5868 43260 5896
rect 43254 5856 43260 5868
rect 43312 5856 43318 5908
rect 44450 5856 44456 5908
rect 44508 5896 44514 5908
rect 45465 5899 45523 5905
rect 45465 5896 45477 5899
rect 44508 5868 45477 5896
rect 44508 5856 44514 5868
rect 45465 5865 45477 5868
rect 45511 5865 45523 5899
rect 48498 5896 48504 5908
rect 45465 5859 45523 5865
rect 45664 5868 48504 5896
rect 37458 5788 37464 5840
rect 37516 5828 37522 5840
rect 43622 5828 43628 5840
rect 37516 5800 43628 5828
rect 37516 5788 37522 5800
rect 43622 5788 43628 5800
rect 43680 5788 43686 5840
rect 44634 5760 44640 5772
rect 35483 5732 36216 5760
rect 37384 5732 41414 5760
rect 44595 5732 44640 5760
rect 35483 5729 35495 5732
rect 35437 5723 35495 5729
rect 14544 5695 14602 5701
rect 14544 5661 14556 5695
rect 14590 5661 14602 5695
rect 14544 5655 14602 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 14366 5624 14372 5636
rect 13188 5596 14372 5624
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14568 5624 14596 5655
rect 14516 5596 14596 5624
rect 14516 5584 14522 5596
rect 15010 5584 15016 5636
rect 15068 5624 15074 5636
rect 16316 5624 16344 5655
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17770 5692 17776 5704
rect 17368 5664 17776 5692
rect 17368 5652 17374 5664
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 19794 5692 19800 5704
rect 19755 5664 19800 5692
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20036 5664 22094 5692
rect 20036 5652 20042 5664
rect 21082 5624 21088 5636
rect 15068 5596 15792 5624
rect 16316 5596 21088 5624
rect 15068 5584 15074 5596
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 9732 5528 11621 5556
rect 9732 5516 9738 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 11609 5519 11667 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15657 5559 15715 5565
rect 15657 5556 15669 5559
rect 15620 5528 15669 5556
rect 15620 5516 15626 5528
rect 15657 5525 15669 5528
rect 15703 5525 15715 5559
rect 15764 5556 15792 5596
rect 21082 5584 21088 5596
rect 21140 5584 21146 5636
rect 22066 5624 22094 5664
rect 22370 5652 22376 5704
rect 22428 5692 22434 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 22428 5664 24593 5692
rect 22428 5652 22434 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 28994 5652 29000 5704
rect 29052 5692 29058 5704
rect 30193 5695 30251 5701
rect 30193 5692 30205 5695
rect 29052 5664 30205 5692
rect 29052 5652 29058 5664
rect 30193 5661 30205 5664
rect 30239 5661 30251 5695
rect 30374 5692 30380 5704
rect 30335 5664 30380 5692
rect 30193 5655 30251 5661
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 34422 5692 34428 5704
rect 30524 5664 34428 5692
rect 30524 5652 30530 5664
rect 34422 5652 34428 5664
rect 34480 5652 34486 5704
rect 36188 5692 36216 5732
rect 37102 5695 37160 5701
rect 37102 5692 37114 5695
rect 36188 5664 37114 5692
rect 37102 5661 37114 5664
rect 37148 5661 37160 5695
rect 37102 5655 37160 5661
rect 37369 5695 37427 5701
rect 37369 5661 37381 5695
rect 37415 5661 37427 5695
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37369 5655 37427 5661
rect 23934 5624 23940 5636
rect 22066 5596 23940 5624
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 24026 5584 24032 5636
rect 24084 5624 24090 5636
rect 33962 5624 33968 5636
rect 24084 5596 33968 5624
rect 24084 5584 24090 5596
rect 33962 5584 33968 5596
rect 34020 5584 34026 5636
rect 34330 5584 34336 5636
rect 34388 5624 34394 5636
rect 37182 5624 37188 5636
rect 34388 5596 37188 5624
rect 34388 5584 34394 5596
rect 37182 5584 37188 5596
rect 37240 5624 37246 5636
rect 37384 5624 37412 5655
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 41230 5692 41236 5704
rect 37936 5664 41236 5692
rect 37240 5596 37412 5624
rect 37240 5584 37246 5596
rect 16758 5556 16764 5568
rect 15764 5528 16764 5556
rect 15657 5519 15715 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 17034 5516 17040 5568
rect 17092 5556 17098 5568
rect 18598 5556 18604 5568
rect 17092 5528 18604 5556
rect 17092 5516 17098 5528
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 22094 5556 22100 5568
rect 18748 5528 22100 5556
rect 18748 5516 18754 5528
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 22186 5516 22192 5568
rect 22244 5556 22250 5568
rect 26050 5556 26056 5568
rect 22244 5528 26056 5556
rect 22244 5516 22250 5528
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 30837 5559 30895 5565
rect 30837 5556 30849 5559
rect 30432 5528 30849 5556
rect 30432 5516 30438 5528
rect 30837 5525 30849 5528
rect 30883 5525 30895 5559
rect 30837 5519 30895 5525
rect 33042 5516 33048 5568
rect 33100 5556 33106 5568
rect 37936 5556 37964 5664
rect 41230 5652 41236 5664
rect 41288 5652 41294 5704
rect 41386 5692 41414 5732
rect 44634 5720 44640 5732
rect 44692 5720 44698 5772
rect 45664 5701 45692 5868
rect 48498 5856 48504 5868
rect 48556 5856 48562 5908
rect 48590 5856 48596 5908
rect 48648 5896 48654 5908
rect 52181 5899 52239 5905
rect 52181 5896 52193 5899
rect 48648 5868 52193 5896
rect 48648 5856 48654 5868
rect 52181 5865 52193 5868
rect 52227 5896 52239 5899
rect 59906 5896 59912 5908
rect 52227 5868 59912 5896
rect 52227 5865 52239 5868
rect 52181 5859 52239 5865
rect 59906 5856 59912 5868
rect 59964 5856 59970 5908
rect 66622 5896 66628 5908
rect 63880 5868 66628 5896
rect 47118 5788 47124 5840
rect 47176 5828 47182 5840
rect 47302 5828 47308 5840
rect 47176 5800 47308 5828
rect 47176 5788 47182 5800
rect 47302 5788 47308 5800
rect 47360 5788 47366 5840
rect 49050 5788 49056 5840
rect 49108 5828 49114 5840
rect 49237 5831 49295 5837
rect 49237 5828 49249 5831
rect 49108 5800 49249 5828
rect 49108 5788 49114 5800
rect 49237 5797 49249 5800
rect 49283 5797 49295 5831
rect 49237 5791 49295 5797
rect 45830 5760 45836 5772
rect 45791 5732 45836 5760
rect 45830 5720 45836 5732
rect 45888 5720 45894 5772
rect 46014 5720 46020 5772
rect 46072 5760 46078 5772
rect 47857 5763 47915 5769
rect 47857 5760 47869 5763
rect 46072 5732 47869 5760
rect 46072 5720 46078 5732
rect 47857 5729 47869 5732
rect 47903 5729 47915 5763
rect 47857 5723 47915 5729
rect 53561 5763 53619 5769
rect 53561 5729 53573 5763
rect 53607 5760 53619 5763
rect 54662 5760 54668 5772
rect 53607 5732 54668 5760
rect 53607 5729 53619 5732
rect 53561 5723 53619 5729
rect 54662 5720 54668 5732
rect 54720 5720 54726 5772
rect 63310 5720 63316 5772
rect 63368 5760 63374 5772
rect 63880 5769 63908 5868
rect 66622 5856 66628 5868
rect 66680 5856 66686 5908
rect 68922 5896 68928 5908
rect 68883 5868 68928 5896
rect 68922 5856 68928 5868
rect 68980 5856 68986 5908
rect 69290 5856 69296 5908
rect 69348 5896 69354 5908
rect 75914 5896 75920 5908
rect 69348 5868 75920 5896
rect 69348 5856 69354 5868
rect 75914 5856 75920 5868
rect 75972 5896 75978 5908
rect 76193 5899 76251 5905
rect 76193 5896 76205 5899
rect 75972 5868 76205 5896
rect 75972 5856 75978 5868
rect 76193 5865 76205 5868
rect 76239 5896 76251 5899
rect 76742 5896 76748 5908
rect 76239 5868 76748 5896
rect 76239 5865 76251 5868
rect 76193 5859 76251 5865
rect 76742 5856 76748 5868
rect 76800 5856 76806 5908
rect 90634 5856 90640 5908
rect 90692 5896 90698 5908
rect 91830 5896 91836 5908
rect 90692 5868 91836 5896
rect 90692 5856 90698 5868
rect 91830 5856 91836 5868
rect 91888 5856 91894 5908
rect 93964 5868 95372 5896
rect 65245 5831 65303 5837
rect 65245 5797 65257 5831
rect 65291 5828 65303 5831
rect 67634 5828 67640 5840
rect 65291 5800 67640 5828
rect 65291 5797 65303 5800
rect 65245 5791 65303 5797
rect 67634 5788 67640 5800
rect 67692 5788 67698 5840
rect 68465 5831 68523 5837
rect 68465 5797 68477 5831
rect 68511 5828 68523 5831
rect 69106 5828 69112 5840
rect 68511 5800 69112 5828
rect 68511 5797 68523 5800
rect 68465 5791 68523 5797
rect 69106 5788 69112 5800
rect 69164 5788 69170 5840
rect 72694 5828 72700 5840
rect 72655 5800 72700 5828
rect 72694 5788 72700 5800
rect 72752 5788 72758 5840
rect 79045 5831 79103 5837
rect 79045 5828 79057 5831
rect 76116 5800 79057 5828
rect 63865 5763 63923 5769
rect 63865 5760 63877 5763
rect 63368 5732 63877 5760
rect 63368 5720 63374 5732
rect 63865 5729 63877 5732
rect 63911 5729 63923 5763
rect 63865 5723 63923 5729
rect 65886 5720 65892 5772
rect 65944 5760 65950 5772
rect 66165 5763 66223 5769
rect 66165 5760 66177 5763
rect 65944 5732 66177 5760
rect 65944 5720 65950 5732
rect 66165 5729 66177 5732
rect 66211 5729 66223 5763
rect 66165 5723 66223 5729
rect 75457 5763 75515 5769
rect 75457 5729 75469 5763
rect 75503 5760 75515 5763
rect 76006 5760 76012 5772
rect 75503 5732 76012 5760
rect 75503 5729 75515 5732
rect 75457 5723 75515 5729
rect 76006 5720 76012 5732
rect 76064 5720 76070 5772
rect 45649 5695 45707 5701
rect 41386 5664 44496 5692
rect 38010 5584 38016 5636
rect 38068 5624 38074 5636
rect 44370 5627 44428 5633
rect 44370 5624 44382 5627
rect 38068 5596 44382 5624
rect 38068 5584 38074 5596
rect 44370 5593 44382 5596
rect 44416 5593 44428 5627
rect 44468 5624 44496 5664
rect 45649 5661 45661 5695
rect 45695 5661 45707 5695
rect 45649 5655 45707 5661
rect 47964 5664 54156 5692
rect 47964 5624 47992 5664
rect 48113 5627 48171 5633
rect 48113 5624 48125 5627
rect 44468 5596 47992 5624
rect 48047 5596 48125 5624
rect 44370 5587 44428 5593
rect 38562 5556 38568 5568
rect 33100 5528 37964 5556
rect 38523 5528 38568 5556
rect 33100 5516 33106 5528
rect 38562 5516 38568 5528
rect 38620 5516 38626 5568
rect 43622 5516 43628 5568
rect 43680 5556 43686 5568
rect 47210 5556 47216 5568
rect 43680 5528 47216 5556
rect 43680 5516 43686 5528
rect 47210 5516 47216 5528
rect 47268 5516 47274 5568
rect 47302 5516 47308 5568
rect 47360 5556 47366 5568
rect 48047 5556 48075 5596
rect 48113 5593 48125 5596
rect 48159 5593 48171 5627
rect 48113 5587 48171 5593
rect 53316 5627 53374 5633
rect 53316 5593 53328 5627
rect 53362 5624 53374 5627
rect 54128 5624 54156 5664
rect 54202 5652 54208 5704
rect 54260 5692 54266 5704
rect 58618 5692 58624 5704
rect 54260 5664 54305 5692
rect 58579 5664 58624 5692
rect 54260 5652 54266 5664
rect 58618 5652 58624 5664
rect 58676 5652 58682 5704
rect 63770 5652 63776 5704
rect 63828 5692 63834 5704
rect 64121 5695 64179 5701
rect 64121 5692 64133 5695
rect 63828 5664 64133 5692
rect 63828 5652 63834 5664
rect 64121 5661 64133 5664
rect 64167 5661 64179 5695
rect 64121 5655 64179 5661
rect 65981 5695 66039 5701
rect 65981 5661 65993 5695
rect 66027 5692 66039 5695
rect 66070 5692 66076 5704
rect 66027 5664 66076 5692
rect 66027 5661 66039 5664
rect 65981 5655 66039 5661
rect 66070 5652 66076 5664
rect 66128 5652 66134 5704
rect 66254 5652 66260 5704
rect 66312 5692 66318 5704
rect 70038 5695 70096 5701
rect 70038 5692 70050 5695
rect 66312 5664 70050 5692
rect 66312 5652 66318 5664
rect 70038 5661 70050 5664
rect 70084 5661 70096 5695
rect 70038 5655 70096 5661
rect 70305 5695 70363 5701
rect 70305 5661 70317 5695
rect 70351 5661 70363 5695
rect 70305 5655 70363 5661
rect 72881 5695 72939 5701
rect 72881 5661 72893 5695
rect 72927 5661 72939 5695
rect 72881 5655 72939 5661
rect 73065 5695 73123 5701
rect 73065 5661 73077 5695
rect 73111 5692 73123 5695
rect 73154 5692 73160 5704
rect 73111 5664 73160 5692
rect 73111 5661 73123 5664
rect 73065 5655 73123 5661
rect 62022 5624 62028 5636
rect 53362 5596 54064 5624
rect 54128 5596 62028 5624
rect 53362 5593 53374 5596
rect 53316 5587 53374 5593
rect 54036 5565 54064 5596
rect 62022 5584 62028 5596
rect 62080 5584 62086 5636
rect 69106 5584 69112 5636
rect 69164 5624 69170 5636
rect 70320 5624 70348 5655
rect 69164 5596 70348 5624
rect 72896 5624 72924 5655
rect 73154 5652 73160 5664
rect 73212 5652 73218 5704
rect 74166 5652 74172 5704
rect 74224 5692 74230 5704
rect 76116 5692 76144 5800
rect 79045 5797 79057 5800
rect 79091 5797 79103 5831
rect 79045 5791 79103 5797
rect 86402 5788 86408 5840
rect 86460 5828 86466 5840
rect 93854 5828 93860 5840
rect 86460 5800 93860 5828
rect 86460 5788 86466 5800
rect 93854 5788 93860 5800
rect 93912 5788 93918 5840
rect 80422 5760 80428 5772
rect 80383 5732 80428 5760
rect 80422 5720 80428 5732
rect 80480 5720 80486 5772
rect 76742 5692 76748 5704
rect 74224 5664 76144 5692
rect 76703 5664 76748 5692
rect 74224 5652 74230 5664
rect 76742 5652 76748 5664
rect 76800 5652 76806 5704
rect 78858 5652 78864 5704
rect 78916 5692 78922 5704
rect 80158 5695 80216 5701
rect 80158 5692 80170 5695
rect 78916 5664 80170 5692
rect 78916 5652 78922 5664
rect 80158 5661 80170 5664
rect 80204 5661 80216 5695
rect 81250 5692 81256 5704
rect 81211 5664 81256 5692
rect 80158 5655 80216 5661
rect 81250 5652 81256 5664
rect 81308 5652 81314 5704
rect 83274 5652 83280 5704
rect 83332 5692 83338 5704
rect 93964 5692 93992 5868
rect 95344 5828 95372 5868
rect 96614 5856 96620 5908
rect 96672 5896 96678 5908
rect 99377 5899 99435 5905
rect 99377 5896 99389 5899
rect 96672 5868 99389 5896
rect 96672 5856 96678 5868
rect 99377 5865 99389 5868
rect 99423 5896 99435 5899
rect 101306 5896 101312 5908
rect 99423 5868 101312 5896
rect 99423 5865 99435 5868
rect 99377 5859 99435 5865
rect 101306 5856 101312 5868
rect 101364 5856 101370 5908
rect 103422 5856 103428 5908
rect 103480 5896 103486 5908
rect 108850 5896 108856 5908
rect 103480 5868 108528 5896
rect 108811 5868 108856 5896
rect 103480 5856 103486 5868
rect 99926 5828 99932 5840
rect 95344 5800 99932 5828
rect 99926 5788 99932 5800
rect 99984 5788 99990 5840
rect 105078 5788 105084 5840
rect 105136 5828 105142 5840
rect 106642 5828 106648 5840
rect 105136 5800 106648 5828
rect 105136 5788 105142 5800
rect 106642 5788 106648 5800
rect 106700 5788 106706 5840
rect 108393 5831 108451 5837
rect 108393 5797 108405 5831
rect 108439 5797 108451 5831
rect 108500 5828 108528 5868
rect 108850 5856 108856 5868
rect 108908 5856 108914 5908
rect 116762 5896 116768 5908
rect 113836 5868 116768 5896
rect 113836 5828 113864 5868
rect 116762 5856 116768 5868
rect 116820 5856 116826 5908
rect 117406 5896 117412 5908
rect 117367 5868 117412 5896
rect 117406 5856 117412 5868
rect 117464 5856 117470 5908
rect 120534 5896 120540 5908
rect 117700 5868 120540 5896
rect 108500 5800 113864 5828
rect 114373 5831 114431 5837
rect 108393 5791 108451 5797
rect 114373 5797 114385 5831
rect 114419 5828 114431 5831
rect 114554 5828 114560 5840
rect 114419 5800 114560 5828
rect 114419 5797 114431 5800
rect 114373 5791 114431 5797
rect 101490 5720 101496 5772
rect 101548 5760 101554 5772
rect 106090 5760 106096 5772
rect 101548 5732 106096 5760
rect 101548 5720 101554 5732
rect 106090 5720 106096 5732
rect 106148 5720 106154 5772
rect 108408 5760 108436 5791
rect 114554 5788 114560 5800
rect 114612 5788 114618 5840
rect 115382 5828 115388 5840
rect 115343 5800 115388 5828
rect 115382 5788 115388 5800
rect 115440 5788 115446 5840
rect 117038 5788 117044 5840
rect 117096 5828 117102 5840
rect 117700 5828 117728 5868
rect 120534 5856 120540 5868
rect 120592 5856 120598 5908
rect 120810 5896 120816 5908
rect 120771 5868 120816 5896
rect 120810 5856 120816 5868
rect 120868 5856 120874 5908
rect 121914 5896 121920 5908
rect 121656 5868 121920 5896
rect 117096 5800 117728 5828
rect 118329 5831 118387 5837
rect 117096 5788 117102 5800
rect 118329 5797 118341 5831
rect 118375 5797 118387 5831
rect 118329 5791 118387 5797
rect 120353 5831 120411 5837
rect 120353 5797 120365 5831
rect 120399 5828 120411 5831
rect 121656 5828 121684 5868
rect 121914 5856 121920 5868
rect 121972 5856 121978 5908
rect 122466 5896 122472 5908
rect 122427 5868 122472 5896
rect 122466 5856 122472 5868
rect 122524 5856 122530 5908
rect 122558 5856 122564 5908
rect 122616 5896 122622 5908
rect 123113 5899 123171 5905
rect 123113 5896 123125 5899
rect 122616 5868 123125 5896
rect 122616 5856 122622 5868
rect 123113 5865 123125 5868
rect 123159 5896 123171 5899
rect 127526 5896 127532 5908
rect 123159 5868 127532 5896
rect 123159 5865 123171 5868
rect 123113 5859 123171 5865
rect 127526 5856 127532 5868
rect 127584 5856 127590 5908
rect 128354 5896 128360 5908
rect 127636 5868 128360 5896
rect 120399 5800 121684 5828
rect 120399 5797 120411 5800
rect 120353 5791 120411 5797
rect 108482 5760 108488 5772
rect 108408 5732 108488 5760
rect 108482 5720 108488 5732
rect 108540 5720 108546 5772
rect 116765 5763 116823 5769
rect 116765 5729 116777 5763
rect 116811 5760 116823 5763
rect 117130 5760 117136 5772
rect 116811 5732 117136 5760
rect 116811 5729 116823 5732
rect 116765 5723 116823 5729
rect 117130 5720 117136 5732
rect 117188 5720 117194 5772
rect 95326 5692 95332 5704
rect 83332 5664 93992 5692
rect 94056 5664 95188 5692
rect 95287 5664 95332 5692
rect 83332 5652 83338 5664
rect 73525 5627 73583 5633
rect 73525 5624 73537 5627
rect 72896 5596 73537 5624
rect 69164 5584 69170 5596
rect 73525 5593 73537 5596
rect 73571 5624 73583 5627
rect 74442 5624 74448 5636
rect 73571 5596 74448 5624
rect 73571 5593 73583 5596
rect 73525 5587 73583 5593
rect 74442 5584 74448 5596
rect 74500 5584 74506 5636
rect 75212 5627 75270 5633
rect 75212 5593 75224 5627
rect 75258 5624 75270 5627
rect 77202 5624 77208 5636
rect 75258 5596 77208 5624
rect 75258 5593 75270 5596
rect 75212 5587 75270 5593
rect 77202 5584 77208 5596
rect 77260 5584 77266 5636
rect 83001 5627 83059 5633
rect 83001 5593 83013 5627
rect 83047 5624 83059 5627
rect 94056 5624 94084 5664
rect 83047 5596 94084 5624
rect 83047 5593 83059 5596
rect 83001 5587 83059 5593
rect 94130 5584 94136 5636
rect 94188 5624 94194 5636
rect 95062 5627 95120 5633
rect 95062 5624 95074 5627
rect 94188 5596 95074 5624
rect 94188 5584 94194 5596
rect 95062 5593 95074 5596
rect 95108 5593 95120 5627
rect 95160 5624 95188 5664
rect 95326 5652 95332 5664
rect 95384 5652 95390 5704
rect 101306 5692 101312 5704
rect 99346 5664 101168 5692
rect 101267 5664 101312 5692
rect 99346 5624 99374 5664
rect 100938 5624 100944 5636
rect 95160 5596 99374 5624
rect 99760 5596 100944 5624
rect 95062 5587 95120 5593
rect 47360 5528 48075 5556
rect 54021 5559 54079 5565
rect 47360 5516 47366 5528
rect 54021 5525 54033 5559
rect 54067 5525 54079 5559
rect 58434 5556 58440 5568
rect 58395 5528 58440 5556
rect 54021 5519 54079 5525
rect 58434 5516 58440 5528
rect 58492 5516 58498 5568
rect 65794 5556 65800 5568
rect 65755 5528 65800 5556
rect 65794 5516 65800 5528
rect 65852 5516 65858 5568
rect 74077 5559 74135 5565
rect 74077 5525 74089 5559
rect 74123 5556 74135 5559
rect 75362 5556 75368 5568
rect 74123 5528 75368 5556
rect 74123 5525 74135 5528
rect 74077 5519 74135 5525
rect 75362 5516 75368 5528
rect 75420 5516 75426 5568
rect 76006 5516 76012 5568
rect 76064 5556 76070 5568
rect 78033 5559 78091 5565
rect 78033 5556 78045 5559
rect 76064 5528 78045 5556
rect 76064 5516 76070 5528
rect 78033 5525 78045 5528
rect 78079 5525 78091 5559
rect 93394 5556 93400 5568
rect 93355 5528 93400 5556
rect 78033 5519 78091 5525
rect 93394 5516 93400 5528
rect 93452 5516 93458 5568
rect 93854 5516 93860 5568
rect 93912 5556 93918 5568
rect 93949 5559 94007 5565
rect 93949 5556 93961 5559
rect 93912 5528 93961 5556
rect 93912 5516 93918 5528
rect 93949 5525 93961 5528
rect 93995 5525 94007 5559
rect 93949 5519 94007 5525
rect 94038 5516 94044 5568
rect 94096 5556 94102 5568
rect 99760 5556 99788 5596
rect 100938 5584 100944 5596
rect 100996 5584 101002 5636
rect 101042 5627 101100 5633
rect 101042 5593 101054 5627
rect 101088 5593 101100 5627
rect 101140 5624 101168 5664
rect 101306 5652 101312 5664
rect 101364 5652 101370 5704
rect 107013 5695 107071 5701
rect 107013 5661 107025 5695
rect 107059 5692 107071 5695
rect 107654 5692 107660 5704
rect 107059 5664 107660 5692
rect 107059 5661 107071 5664
rect 107013 5655 107071 5661
rect 107654 5652 107660 5664
rect 107712 5652 107718 5704
rect 113726 5652 113732 5704
rect 113784 5692 113790 5704
rect 118344 5692 118372 5791
rect 121730 5788 121736 5840
rect 121788 5828 121794 5840
rect 126514 5828 126520 5840
rect 121788 5800 126520 5828
rect 121788 5788 121794 5800
rect 126514 5788 126520 5800
rect 126572 5788 126578 5840
rect 127066 5828 127072 5840
rect 127027 5800 127072 5828
rect 127066 5788 127072 5800
rect 127124 5788 127130 5840
rect 123018 5760 123024 5772
rect 121196 5732 123024 5760
rect 121196 5704 121224 5732
rect 123018 5720 123024 5732
rect 123076 5720 123082 5772
rect 123665 5763 123723 5769
rect 123665 5729 123677 5763
rect 123711 5760 123723 5763
rect 123938 5760 123944 5772
rect 123711 5732 123944 5760
rect 123711 5729 123723 5732
rect 123665 5723 123723 5729
rect 123938 5720 123944 5732
rect 123996 5720 124002 5772
rect 124585 5763 124643 5769
rect 124585 5729 124597 5763
rect 124631 5760 124643 5763
rect 124950 5760 124956 5772
rect 124631 5732 124956 5760
rect 124631 5729 124643 5732
rect 124585 5723 124643 5729
rect 124950 5720 124956 5732
rect 125008 5720 125014 5772
rect 127636 5760 127664 5868
rect 128354 5856 128360 5868
rect 128412 5856 128418 5908
rect 129642 5856 129648 5908
rect 129700 5896 129706 5908
rect 131853 5899 131911 5905
rect 131853 5896 131865 5899
rect 129700 5868 131865 5896
rect 129700 5856 129706 5868
rect 131853 5865 131865 5868
rect 131899 5865 131911 5899
rect 132862 5896 132868 5908
rect 132823 5868 132868 5896
rect 131853 5859 131911 5865
rect 132862 5856 132868 5868
rect 132920 5856 132926 5908
rect 133966 5856 133972 5908
rect 134024 5896 134030 5908
rect 135254 5896 135260 5908
rect 134024 5868 135260 5896
rect 134024 5856 134030 5868
rect 135254 5856 135260 5868
rect 135312 5856 135318 5908
rect 135714 5896 135720 5908
rect 135675 5868 135720 5896
rect 135714 5856 135720 5868
rect 135772 5856 135778 5908
rect 136266 5896 136272 5908
rect 136179 5868 136272 5896
rect 136266 5856 136272 5868
rect 136324 5896 136330 5908
rect 137002 5896 137008 5908
rect 136324 5868 137008 5896
rect 136324 5856 136330 5868
rect 137002 5856 137008 5868
rect 137060 5856 137066 5908
rect 141326 5896 141332 5908
rect 137143 5868 141332 5896
rect 129001 5831 129059 5837
rect 129001 5828 129013 5831
rect 125060 5732 127664 5760
rect 128740 5800 129013 5828
rect 113784 5664 118372 5692
rect 118513 5695 118571 5701
rect 113784 5652 113790 5664
rect 118513 5661 118525 5695
rect 118559 5692 118571 5695
rect 118602 5692 118608 5704
rect 118559 5664 118608 5692
rect 118559 5661 118571 5664
rect 118513 5655 118571 5661
rect 118602 5652 118608 5664
rect 118660 5652 118666 5704
rect 118970 5692 118976 5704
rect 118931 5664 118976 5692
rect 118970 5652 118976 5664
rect 119028 5652 119034 5704
rect 120997 5695 121055 5701
rect 120997 5692 121009 5695
rect 119172 5664 121009 5692
rect 107280 5627 107338 5633
rect 101140 5596 104204 5624
rect 101042 5587 101100 5593
rect 99926 5556 99932 5568
rect 94096 5528 99788 5556
rect 99887 5528 99932 5556
rect 94096 5516 94102 5528
rect 99926 5516 99932 5528
rect 99984 5516 99990 5568
rect 101048 5556 101076 5587
rect 101950 5556 101956 5568
rect 101048 5528 101956 5556
rect 101950 5516 101956 5528
rect 102008 5516 102014 5568
rect 104176 5556 104204 5596
rect 107280 5593 107292 5627
rect 107326 5624 107338 5627
rect 107378 5624 107384 5636
rect 107326 5596 107384 5624
rect 107326 5593 107338 5596
rect 107280 5587 107338 5593
rect 107378 5584 107384 5596
rect 107436 5584 107442 5636
rect 112162 5624 112168 5636
rect 107488 5596 112168 5624
rect 107488 5556 107516 5596
rect 112162 5584 112168 5596
rect 112220 5584 112226 5636
rect 116520 5627 116578 5633
rect 116520 5593 116532 5627
rect 116566 5624 116578 5627
rect 117406 5624 117412 5636
rect 116566 5596 117412 5624
rect 116566 5593 116578 5596
rect 116520 5587 116578 5593
rect 117406 5584 117412 5596
rect 117464 5584 117470 5636
rect 104176 5528 107516 5556
rect 108022 5516 108028 5568
rect 108080 5556 108086 5568
rect 113542 5556 113548 5568
rect 108080 5528 113548 5556
rect 108080 5516 108086 5528
rect 113542 5516 113548 5528
rect 113600 5516 113606 5568
rect 113726 5516 113732 5568
rect 113784 5556 113790 5568
rect 119172 5556 119200 5664
rect 120997 5661 121009 5664
rect 121043 5661 121055 5695
rect 121178 5692 121184 5704
rect 121139 5664 121184 5692
rect 120997 5655 121055 5661
rect 121178 5652 121184 5664
rect 121236 5652 121242 5704
rect 121730 5652 121736 5704
rect 121788 5652 121794 5704
rect 125060 5692 125088 5732
rect 125778 5692 125784 5704
rect 121840 5664 125088 5692
rect 125739 5664 125784 5692
rect 119240 5627 119298 5633
rect 119240 5593 119252 5627
rect 119286 5624 119298 5627
rect 121748 5624 121776 5652
rect 119286 5596 121776 5624
rect 119286 5593 119298 5596
rect 119240 5587 119298 5593
rect 113784 5528 119200 5556
rect 113784 5516 113790 5528
rect 121362 5516 121368 5568
rect 121420 5556 121426 5568
rect 121840 5556 121868 5664
rect 125778 5652 125784 5664
rect 125836 5652 125842 5704
rect 126054 5652 126060 5704
rect 126112 5692 126118 5704
rect 127618 5692 127624 5704
rect 126112 5664 127480 5692
rect 127579 5664 127624 5692
rect 126112 5652 126118 5664
rect 123018 5584 123024 5636
rect 123076 5624 123082 5636
rect 123076 5596 125180 5624
rect 123076 5584 123082 5596
rect 121420 5528 121868 5556
rect 121420 5516 121426 5528
rect 122558 5516 122564 5568
rect 122616 5556 122622 5568
rect 124582 5556 124588 5568
rect 122616 5528 124588 5556
rect 122616 5516 122622 5528
rect 124582 5516 124588 5528
rect 124640 5516 124646 5568
rect 125042 5556 125048 5568
rect 125003 5528 125048 5556
rect 125042 5516 125048 5528
rect 125100 5516 125106 5568
rect 125152 5556 125180 5596
rect 125410 5584 125416 5636
rect 125468 5624 125474 5636
rect 127452 5624 127480 5664
rect 127618 5652 127624 5664
rect 127676 5652 127682 5704
rect 127894 5701 127900 5704
rect 127888 5692 127900 5701
rect 127855 5664 127900 5692
rect 127888 5655 127900 5664
rect 127894 5652 127900 5655
rect 127952 5652 127958 5704
rect 128740 5624 128768 5800
rect 129001 5797 129013 5800
rect 129047 5797 129059 5831
rect 129001 5791 129059 5797
rect 129090 5788 129096 5840
rect 129148 5828 129154 5840
rect 129737 5831 129795 5837
rect 129737 5828 129749 5831
rect 129148 5800 129749 5828
rect 129148 5788 129154 5800
rect 129737 5797 129749 5800
rect 129783 5828 129795 5831
rect 137143 5828 137171 5868
rect 141326 5856 141332 5868
rect 141384 5856 141390 5908
rect 142341 5899 142399 5905
rect 142341 5865 142353 5899
rect 142387 5896 142399 5899
rect 144914 5896 144920 5908
rect 142387 5868 144920 5896
rect 142387 5865 142399 5868
rect 142341 5859 142399 5865
rect 144914 5856 144920 5868
rect 144972 5856 144978 5908
rect 145282 5856 145288 5908
rect 145340 5896 145346 5908
rect 146297 5899 146355 5905
rect 145340 5868 145972 5896
rect 145340 5856 145346 5868
rect 137278 5828 137284 5840
rect 129783 5800 135254 5828
rect 129783 5797 129795 5800
rect 129737 5791 129795 5797
rect 131206 5720 131212 5772
rect 131264 5760 131270 5772
rect 132310 5760 132316 5772
rect 131264 5732 132316 5760
rect 131264 5720 131270 5732
rect 132310 5720 132316 5732
rect 132368 5760 132374 5772
rect 132954 5760 132960 5772
rect 132368 5732 132960 5760
rect 132368 5720 132374 5732
rect 132954 5720 132960 5732
rect 133012 5720 133018 5772
rect 135226 5760 135254 5800
rect 135548 5800 137171 5828
rect 137239 5800 137284 5828
rect 135548 5760 135576 5800
rect 137278 5788 137284 5800
rect 137336 5788 137342 5840
rect 138290 5788 138296 5840
rect 138348 5828 138354 5840
rect 138477 5831 138535 5837
rect 138477 5828 138489 5831
rect 138348 5800 138489 5828
rect 138348 5788 138354 5800
rect 138477 5797 138489 5800
rect 138523 5797 138535 5831
rect 138477 5791 138535 5797
rect 140038 5788 140044 5840
rect 140096 5828 140102 5840
rect 140317 5831 140375 5837
rect 140317 5828 140329 5831
rect 140096 5800 140329 5828
rect 140096 5788 140102 5800
rect 140317 5797 140329 5800
rect 140363 5797 140375 5831
rect 140317 5791 140375 5797
rect 144178 5788 144184 5840
rect 144236 5828 144242 5840
rect 144457 5831 144515 5837
rect 144457 5828 144469 5831
rect 144236 5800 144469 5828
rect 144236 5788 144242 5800
rect 144457 5797 144469 5800
rect 144503 5797 144515 5831
rect 144457 5791 144515 5797
rect 135226 5732 135576 5760
rect 137002 5720 137008 5772
rect 137060 5760 137066 5772
rect 138842 5760 138848 5772
rect 137060 5732 138848 5760
rect 137060 5720 137066 5732
rect 138842 5720 138848 5732
rect 138900 5720 138906 5772
rect 140961 5763 141019 5769
rect 140961 5760 140973 5763
rect 139872 5732 140973 5760
rect 130102 5652 130108 5704
rect 130160 5692 130166 5704
rect 130381 5695 130439 5701
rect 130381 5692 130393 5695
rect 130160 5664 130393 5692
rect 130160 5652 130166 5664
rect 130381 5661 130393 5664
rect 130427 5661 130439 5695
rect 130381 5655 130439 5661
rect 130838 5652 130844 5704
rect 130896 5692 130902 5704
rect 133966 5692 133972 5704
rect 130896 5664 133972 5692
rect 130896 5652 130902 5664
rect 133966 5652 133972 5664
rect 134024 5652 134030 5704
rect 134518 5692 134524 5704
rect 134479 5664 134524 5692
rect 134518 5652 134524 5664
rect 134576 5652 134582 5704
rect 136634 5692 136640 5704
rect 135088 5664 136640 5692
rect 130194 5624 130200 5636
rect 125468 5596 126836 5624
rect 127452 5596 128768 5624
rect 130155 5596 130200 5624
rect 125468 5584 125474 5596
rect 125597 5559 125655 5565
rect 125597 5556 125609 5559
rect 125152 5528 125609 5556
rect 125597 5525 125609 5528
rect 125643 5525 125655 5559
rect 125597 5519 125655 5525
rect 125686 5516 125692 5568
rect 125744 5556 125750 5568
rect 126238 5556 126244 5568
rect 125744 5528 126244 5556
rect 125744 5516 125750 5528
rect 126238 5516 126244 5528
rect 126296 5556 126302 5568
rect 126425 5559 126483 5565
rect 126425 5556 126437 5559
rect 126296 5528 126437 5556
rect 126296 5516 126302 5528
rect 126425 5525 126437 5528
rect 126471 5556 126483 5559
rect 126698 5556 126704 5568
rect 126471 5528 126704 5556
rect 126471 5525 126483 5528
rect 126425 5519 126483 5525
rect 126698 5516 126704 5528
rect 126756 5516 126762 5568
rect 126808 5556 126836 5596
rect 130194 5584 130200 5596
rect 130252 5584 130258 5636
rect 131298 5624 131304 5636
rect 131259 5596 131304 5624
rect 131298 5584 131304 5596
rect 131356 5584 131362 5636
rect 131942 5624 131948 5636
rect 131903 5596 131948 5624
rect 131942 5584 131948 5596
rect 132000 5584 132006 5636
rect 135088 5633 135116 5664
rect 136634 5652 136640 5664
rect 136692 5692 136698 5704
rect 136729 5695 136787 5701
rect 136729 5692 136741 5695
rect 136692 5664 136741 5692
rect 136692 5652 136698 5664
rect 136729 5661 136741 5664
rect 136775 5661 136787 5695
rect 136729 5655 136787 5661
rect 137922 5652 137928 5704
rect 137980 5692 137986 5704
rect 138017 5695 138075 5701
rect 138017 5692 138029 5695
rect 137980 5664 138029 5692
rect 137980 5652 137986 5664
rect 138017 5661 138029 5664
rect 138063 5692 138075 5695
rect 139302 5692 139308 5704
rect 138063 5664 139308 5692
rect 138063 5661 138075 5664
rect 138017 5655 138075 5661
rect 139302 5652 139308 5664
rect 139360 5692 139366 5704
rect 139872 5701 139900 5732
rect 140961 5729 140973 5732
rect 141007 5729 141019 5763
rect 140961 5723 141019 5729
rect 139857 5695 139915 5701
rect 139857 5692 139869 5695
rect 139360 5664 139869 5692
rect 139360 5652 139366 5664
rect 139857 5661 139869 5664
rect 139903 5661 139915 5695
rect 140498 5692 140504 5704
rect 140459 5664 140504 5692
rect 139857 5655 139915 5661
rect 140498 5652 140504 5664
rect 140556 5652 140562 5704
rect 140976 5692 141004 5723
rect 144086 5720 144092 5772
rect 144144 5760 144150 5772
rect 145944 5760 145972 5868
rect 146297 5865 146309 5899
rect 146343 5896 146355 5899
rect 147674 5896 147680 5908
rect 146343 5868 147680 5896
rect 146343 5865 146355 5868
rect 146297 5859 146355 5865
rect 147674 5856 147680 5868
rect 147732 5856 147738 5908
rect 156782 5896 156788 5908
rect 147876 5868 156788 5896
rect 147876 5760 147904 5868
rect 156782 5856 156788 5868
rect 156840 5856 156846 5908
rect 149422 5788 149428 5840
rect 149480 5828 149486 5840
rect 149609 5831 149667 5837
rect 149609 5828 149621 5831
rect 149480 5800 149621 5828
rect 149480 5788 149486 5800
rect 149609 5797 149621 5800
rect 149655 5828 149667 5831
rect 149882 5828 149888 5840
rect 149655 5800 149888 5828
rect 149655 5797 149667 5800
rect 149609 5791 149667 5797
rect 149882 5788 149888 5800
rect 149940 5788 149946 5840
rect 150618 5788 150624 5840
rect 150676 5828 150682 5840
rect 151633 5831 151691 5837
rect 151633 5828 151645 5831
rect 150676 5800 151645 5828
rect 150676 5788 150682 5800
rect 151633 5797 151645 5800
rect 151679 5797 151691 5831
rect 151633 5791 151691 5797
rect 152366 5788 152372 5840
rect 152424 5828 152430 5840
rect 153930 5828 153936 5840
rect 152424 5800 153936 5828
rect 152424 5788 152430 5800
rect 153930 5788 153936 5800
rect 153988 5788 153994 5840
rect 154025 5831 154083 5837
rect 154025 5797 154037 5831
rect 154071 5828 154083 5831
rect 154114 5828 154120 5840
rect 154071 5800 154120 5828
rect 154071 5797 154083 5800
rect 154025 5791 154083 5797
rect 154114 5788 154120 5800
rect 154172 5788 154178 5840
rect 154482 5828 154488 5840
rect 154224 5800 154488 5828
rect 144144 5732 145052 5760
rect 145944 5732 147904 5760
rect 144144 5720 144150 5732
rect 142430 5692 142436 5704
rect 140976 5664 142436 5692
rect 142430 5652 142436 5664
rect 142488 5692 142494 5704
rect 142798 5692 142804 5704
rect 142488 5664 142804 5692
rect 142488 5652 142494 5664
rect 142798 5652 142804 5664
rect 142856 5692 142862 5704
rect 143077 5695 143135 5701
rect 143077 5692 143089 5695
rect 142856 5664 143089 5692
rect 142856 5652 142862 5664
rect 143077 5661 143089 5664
rect 143123 5692 143135 5695
rect 144917 5695 144975 5701
rect 144917 5692 144929 5695
rect 143123 5664 144929 5692
rect 143123 5661 143135 5664
rect 143077 5655 143135 5661
rect 144917 5661 144929 5664
rect 144963 5661 144975 5695
rect 145024 5692 145052 5732
rect 149238 5720 149244 5772
rect 149296 5760 149302 5772
rect 150437 5763 150495 5769
rect 149296 5732 150296 5760
rect 149296 5720 149302 5732
rect 145024 5664 146340 5692
rect 144917 5655 144975 5661
rect 135073 5627 135131 5633
rect 135073 5624 135085 5627
rect 133432 5596 135085 5624
rect 128538 5556 128544 5568
rect 126808 5528 128544 5556
rect 128538 5516 128544 5528
rect 128596 5556 128602 5568
rect 131022 5556 131028 5568
rect 128596 5528 131028 5556
rect 128596 5516 128602 5528
rect 131022 5516 131028 5528
rect 131080 5516 131086 5568
rect 133046 5516 133052 5568
rect 133104 5556 133110 5568
rect 133432 5565 133460 5596
rect 135073 5593 135085 5596
rect 135119 5593 135131 5627
rect 135073 5587 135131 5593
rect 135530 5584 135536 5636
rect 135588 5624 135594 5636
rect 136910 5624 136916 5636
rect 135588 5596 136916 5624
rect 135588 5584 135594 5596
rect 136910 5584 136916 5596
rect 136968 5584 136974 5636
rect 139612 5627 139670 5633
rect 139612 5593 139624 5627
rect 139658 5624 139670 5627
rect 140038 5624 140044 5636
rect 139658 5596 140044 5624
rect 139658 5593 139670 5596
rect 139612 5587 139670 5593
rect 140038 5584 140044 5596
rect 140096 5584 140102 5636
rect 140774 5584 140780 5636
rect 140832 5624 140838 5636
rect 143350 5633 143356 5636
rect 141206 5627 141264 5633
rect 141206 5624 141218 5627
rect 140832 5596 141218 5624
rect 140832 5584 140838 5596
rect 141206 5593 141218 5596
rect 141252 5593 141264 5627
rect 143344 5624 143356 5633
rect 143311 5596 143356 5624
rect 141206 5587 141264 5593
rect 143344 5587 143356 5596
rect 143350 5584 143356 5587
rect 143408 5584 143414 5636
rect 145184 5627 145242 5633
rect 145184 5593 145196 5627
rect 145230 5624 145242 5627
rect 146202 5624 146208 5636
rect 145230 5596 146208 5624
rect 145230 5593 145242 5596
rect 145184 5587 145242 5593
rect 146202 5584 146208 5596
rect 146260 5584 146266 5636
rect 146312 5624 146340 5664
rect 146386 5652 146392 5704
rect 146444 5692 146450 5704
rect 146754 5692 146760 5704
rect 146444 5664 146760 5692
rect 146444 5652 146450 5664
rect 146754 5652 146760 5664
rect 146812 5652 146818 5704
rect 146938 5692 146944 5704
rect 146899 5664 146944 5692
rect 146938 5652 146944 5664
rect 146996 5652 147002 5704
rect 147030 5652 147036 5704
rect 147088 5692 147094 5704
rect 147398 5692 147404 5704
rect 147088 5664 147404 5692
rect 147088 5652 147094 5664
rect 147398 5652 147404 5664
rect 147456 5692 147462 5704
rect 148229 5695 148287 5701
rect 148229 5692 148241 5695
rect 147456 5664 148241 5692
rect 147456 5652 147462 5664
rect 148229 5661 148241 5664
rect 148275 5692 148287 5695
rect 148870 5692 148876 5704
rect 148275 5664 148876 5692
rect 148275 5661 148287 5664
rect 148229 5655 148287 5661
rect 148870 5652 148876 5664
rect 148928 5652 148934 5704
rect 149514 5652 149520 5704
rect 149572 5692 149578 5704
rect 150268 5701 150296 5732
rect 150437 5729 150449 5763
rect 150483 5760 150495 5763
rect 153102 5760 153108 5772
rect 150483 5732 153108 5760
rect 150483 5729 150495 5732
rect 150437 5723 150495 5729
rect 153102 5720 153108 5732
rect 153160 5720 153166 5772
rect 153194 5720 153200 5772
rect 153252 5760 153258 5772
rect 153252 5732 153884 5760
rect 153252 5720 153258 5732
rect 150069 5695 150127 5701
rect 150069 5692 150081 5695
rect 149572 5664 150081 5692
rect 149572 5652 149578 5664
rect 150069 5661 150081 5664
rect 150115 5661 150127 5695
rect 150069 5655 150127 5661
rect 150253 5695 150311 5701
rect 150253 5661 150265 5695
rect 150299 5661 150311 5695
rect 150253 5655 150311 5661
rect 151081 5695 151139 5701
rect 151081 5661 151093 5695
rect 151127 5692 151139 5695
rect 151538 5692 151544 5704
rect 151127 5664 151544 5692
rect 151127 5661 151139 5664
rect 151081 5655 151139 5661
rect 151538 5652 151544 5664
rect 151596 5652 151602 5704
rect 151817 5695 151875 5701
rect 151817 5661 151829 5695
rect 151863 5692 151875 5695
rect 151906 5692 151912 5704
rect 151863 5664 151912 5692
rect 151863 5661 151875 5664
rect 151817 5655 151875 5661
rect 151906 5652 151912 5664
rect 151964 5652 151970 5704
rect 152461 5695 152519 5701
rect 152461 5661 152473 5695
rect 152507 5692 152519 5695
rect 153562 5692 153568 5704
rect 152507 5664 153568 5692
rect 152507 5661 152519 5664
rect 152461 5655 152519 5661
rect 153562 5652 153568 5664
rect 153620 5652 153626 5704
rect 153654 5652 153660 5704
rect 153712 5692 153718 5704
rect 153856 5701 153884 5732
rect 153841 5695 153899 5701
rect 153712 5664 153757 5692
rect 153712 5652 153718 5664
rect 153841 5661 153853 5695
rect 153887 5661 153899 5695
rect 153841 5655 153899 5661
rect 154114 5652 154120 5704
rect 154172 5692 154178 5704
rect 154224 5692 154252 5800
rect 154482 5788 154488 5800
rect 154540 5788 154546 5840
rect 154942 5788 154948 5840
rect 155000 5828 155006 5840
rect 155313 5831 155371 5837
rect 155313 5828 155325 5831
rect 155000 5800 155325 5828
rect 155000 5788 155006 5800
rect 155313 5797 155325 5800
rect 155359 5797 155371 5831
rect 155313 5791 155371 5797
rect 156690 5788 156696 5840
rect 156748 5828 156754 5840
rect 156969 5831 157027 5837
rect 156969 5828 156981 5831
rect 156748 5800 156981 5828
rect 156748 5788 156754 5800
rect 156969 5797 156981 5800
rect 157015 5797 157027 5831
rect 156969 5791 157027 5797
rect 157242 5788 157248 5840
rect 157300 5828 157306 5840
rect 157613 5831 157671 5837
rect 157613 5828 157625 5831
rect 157300 5800 157625 5828
rect 157300 5788 157306 5800
rect 157613 5797 157625 5800
rect 157659 5797 157671 5831
rect 157613 5791 157671 5797
rect 154853 5763 154911 5769
rect 154853 5729 154865 5763
rect 154899 5760 154911 5763
rect 158254 5760 158260 5772
rect 154899 5732 158260 5760
rect 154899 5729 154911 5732
rect 154853 5723 154911 5729
rect 158254 5720 158260 5732
rect 158312 5720 158318 5772
rect 154172 5664 154252 5692
rect 154577 5695 154635 5701
rect 154172 5652 154178 5664
rect 154577 5661 154589 5695
rect 154623 5661 154635 5695
rect 154577 5655 154635 5661
rect 148474 5627 148532 5633
rect 148474 5624 148486 5627
rect 146312 5596 148486 5624
rect 148474 5593 148486 5596
rect 148520 5593 148532 5627
rect 151446 5624 151452 5636
rect 148474 5587 148532 5593
rect 149348 5596 151452 5624
rect 133417 5559 133475 5565
rect 133417 5556 133429 5559
rect 133104 5528 133429 5556
rect 133104 5516 133110 5528
rect 133417 5525 133429 5528
rect 133463 5525 133475 5559
rect 133417 5519 133475 5525
rect 133782 5516 133788 5568
rect 133840 5556 133846 5568
rect 136266 5556 136272 5568
rect 133840 5528 136272 5556
rect 133840 5516 133846 5528
rect 136266 5516 136272 5528
rect 136324 5516 136330 5568
rect 138658 5516 138664 5568
rect 138716 5556 138722 5568
rect 142614 5556 142620 5568
rect 138716 5528 142620 5556
rect 138716 5516 138722 5528
rect 142614 5516 142620 5528
rect 142672 5516 142678 5568
rect 143074 5516 143080 5568
rect 143132 5556 143138 5568
rect 146662 5556 146668 5568
rect 143132 5528 146668 5556
rect 143132 5516 143138 5528
rect 146662 5516 146668 5528
rect 146720 5516 146726 5568
rect 147125 5559 147183 5565
rect 147125 5525 147137 5559
rect 147171 5556 147183 5559
rect 147398 5556 147404 5568
rect 147171 5528 147404 5556
rect 147171 5525 147183 5528
rect 147125 5519 147183 5525
rect 147398 5516 147404 5528
rect 147456 5516 147462 5568
rect 147677 5559 147735 5565
rect 147677 5525 147689 5559
rect 147723 5556 147735 5559
rect 148318 5556 148324 5568
rect 147723 5528 148324 5556
rect 147723 5525 147735 5528
rect 147677 5519 147735 5525
rect 148318 5516 148324 5528
rect 148376 5556 148382 5568
rect 149348 5556 149376 5596
rect 151446 5584 151452 5596
rect 151504 5584 151510 5636
rect 154592 5624 154620 5655
rect 154666 5652 154672 5704
rect 154724 5692 154730 5704
rect 155494 5692 155500 5704
rect 154724 5664 154769 5692
rect 155455 5664 155500 5692
rect 154724 5652 154730 5664
rect 155494 5652 155500 5664
rect 155552 5652 155558 5704
rect 155589 5695 155647 5701
rect 155589 5661 155601 5695
rect 155635 5661 155647 5695
rect 155589 5655 155647 5661
rect 154592 5596 154804 5624
rect 148376 5528 149376 5556
rect 148376 5516 148382 5528
rect 149422 5516 149428 5568
rect 149480 5556 149486 5568
rect 149698 5556 149704 5568
rect 149480 5528 149704 5556
rect 149480 5516 149486 5528
rect 149698 5516 149704 5528
rect 149756 5516 149762 5568
rect 150158 5516 150164 5568
rect 150216 5556 150222 5568
rect 150897 5559 150955 5565
rect 150897 5556 150909 5559
rect 150216 5528 150909 5556
rect 150216 5516 150222 5528
rect 150897 5525 150909 5528
rect 150943 5525 150955 5559
rect 150897 5519 150955 5525
rect 151078 5516 151084 5568
rect 151136 5556 151142 5568
rect 152277 5559 152335 5565
rect 152277 5556 152289 5559
rect 151136 5528 152289 5556
rect 151136 5516 151142 5528
rect 152277 5525 152289 5528
rect 152323 5525 152335 5559
rect 154776 5556 154804 5596
rect 155402 5584 155408 5636
rect 155460 5624 155466 5636
rect 155604 5624 155632 5655
rect 155770 5652 155776 5704
rect 155828 5692 155834 5704
rect 156141 5695 156199 5701
rect 156141 5692 156153 5695
rect 155828 5664 156153 5692
rect 155828 5652 155834 5664
rect 156141 5661 156153 5664
rect 156187 5661 156199 5695
rect 156141 5655 156199 5661
rect 156325 5695 156383 5701
rect 156325 5661 156337 5695
rect 156371 5661 156383 5695
rect 157150 5692 157156 5704
rect 157111 5664 157156 5692
rect 156325 5655 156383 5661
rect 155460 5596 155632 5624
rect 155460 5584 155466 5596
rect 155862 5584 155868 5636
rect 155920 5624 155926 5636
rect 156340 5624 156368 5655
rect 157150 5652 157156 5664
rect 157208 5652 157214 5704
rect 157518 5652 157524 5704
rect 157576 5692 157582 5704
rect 157797 5695 157855 5701
rect 157797 5692 157809 5695
rect 157576 5664 157809 5692
rect 157576 5652 157582 5664
rect 157797 5661 157809 5664
rect 157843 5661 157855 5695
rect 157797 5655 157855 5661
rect 155920 5596 156368 5624
rect 156509 5627 156567 5633
rect 155920 5584 155926 5596
rect 156509 5593 156521 5627
rect 156555 5624 156567 5627
rect 156555 5596 157104 5624
rect 156555 5593 156567 5596
rect 156509 5587 156567 5593
rect 155420 5556 155448 5584
rect 154776 5528 155448 5556
rect 157076 5556 157104 5596
rect 158622 5556 158628 5568
rect 157076 5528 158628 5556
rect 152277 5519 152335 5525
rect 158622 5516 158628 5528
rect 158680 5516 158686 5568
rect 1104 5466 159043 5488
rect 1104 5414 40394 5466
rect 40446 5414 40458 5466
rect 40510 5414 40522 5466
rect 40574 5414 40586 5466
rect 40638 5414 40650 5466
rect 40702 5414 79839 5466
rect 79891 5414 79903 5466
rect 79955 5414 79967 5466
rect 80019 5414 80031 5466
rect 80083 5414 80095 5466
rect 80147 5414 119284 5466
rect 119336 5414 119348 5466
rect 119400 5414 119412 5466
rect 119464 5414 119476 5466
rect 119528 5414 119540 5466
rect 119592 5414 158729 5466
rect 158781 5414 158793 5466
rect 158845 5414 158857 5466
rect 158909 5414 158921 5466
rect 158973 5414 158985 5466
rect 159037 5414 159043 5466
rect 1104 5392 159043 5414
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 6638 5352 6644 5364
rect 5960 5324 6644 5352
rect 5960 5312 5966 5324
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 13633 5355 13691 5361
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 13722 5352 13728 5364
rect 13679 5324 13728 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 16298 5352 16304 5364
rect 13872 5324 16304 5352
rect 13872 5312 13878 5324
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16816 5324 16865 5352
rect 16816 5312 16822 5324
rect 16853 5321 16865 5324
rect 16899 5352 16911 5355
rect 17589 5355 17647 5361
rect 17589 5352 17601 5355
rect 16899 5324 17601 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 17589 5321 17601 5324
rect 17635 5321 17647 5355
rect 18138 5352 18144 5364
rect 18099 5324 18144 5352
rect 17589 5315 17647 5321
rect 18138 5312 18144 5324
rect 18196 5352 18202 5364
rect 18690 5352 18696 5364
rect 18196 5324 18696 5352
rect 18196 5312 18202 5324
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 19886 5352 19892 5364
rect 19847 5324 19892 5352
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 24121 5355 24179 5361
rect 22940 5324 23244 5352
rect 3878 5284 3884 5296
rect 3791 5256 3884 5284
rect 3804 5225 3832 5256
rect 3878 5244 3884 5256
rect 3936 5284 3942 5296
rect 14274 5284 14280 5296
rect 3936 5256 6040 5284
rect 3936 5244 3942 5256
rect 6012 5228 6040 5256
rect 12268 5256 14280 5284
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 4056 5219 4114 5225
rect 4056 5185 4068 5219
rect 4102 5216 4114 5219
rect 5902 5216 5908 5228
rect 4102 5188 5764 5216
rect 5863 5188 5908 5216
rect 4102 5185 4114 5188
rect 4056 5179 4114 5185
rect 5736 5148 5764 5188
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 12268 5225 12296 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17000 5256 21312 5284
rect 17000 5244 17006 5256
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 6052 5188 12265 5216
rect 6052 5176 6058 5188
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12520 5219 12578 5225
rect 12520 5185 12532 5219
rect 12566 5216 12578 5219
rect 12986 5216 12992 5228
rect 12566 5188 12992 5216
rect 12566 5185 12578 5188
rect 12520 5179 12578 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 15010 5216 15016 5228
rect 14971 5188 15016 5216
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 9674 5148 9680 5160
rect 5736 5120 9680 5148
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 15212 5148 15240 5179
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 17276 5188 19717 5216
rect 17276 5176 17282 5188
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 21284 5216 21312 5256
rect 21358 5244 21364 5296
rect 21416 5284 21422 5296
rect 22940 5284 22968 5324
rect 23014 5293 23020 5296
rect 21416 5256 22968 5284
rect 21416 5244 21422 5256
rect 23008 5247 23020 5293
rect 23072 5284 23078 5296
rect 23216 5284 23244 5324
rect 24121 5321 24133 5355
rect 24167 5352 24179 5355
rect 25498 5352 25504 5364
rect 24167 5324 25504 5352
rect 24167 5321 24179 5324
rect 24121 5315 24179 5321
rect 25498 5312 25504 5324
rect 25556 5352 25562 5364
rect 25958 5352 25964 5364
rect 25556 5324 25964 5352
rect 25556 5312 25562 5324
rect 25958 5312 25964 5324
rect 26016 5312 26022 5364
rect 27249 5355 27307 5361
rect 27249 5321 27261 5355
rect 27295 5352 27307 5355
rect 34514 5352 34520 5364
rect 27295 5324 34520 5352
rect 27295 5321 27307 5324
rect 27249 5315 27307 5321
rect 24581 5287 24639 5293
rect 24581 5284 24593 5287
rect 23072 5256 23108 5284
rect 23216 5256 24593 5284
rect 23014 5244 23020 5247
rect 23072 5244 23078 5256
rect 24581 5253 24593 5256
rect 24627 5284 24639 5287
rect 27264 5284 27292 5315
rect 34514 5312 34520 5324
rect 34572 5312 34578 5364
rect 35342 5352 35348 5364
rect 35303 5324 35348 5352
rect 35342 5312 35348 5324
rect 35400 5312 35406 5364
rect 43346 5312 43352 5364
rect 43404 5352 43410 5364
rect 48501 5355 48559 5361
rect 48501 5352 48513 5355
rect 43404 5324 48513 5352
rect 43404 5312 43410 5324
rect 48501 5321 48513 5324
rect 48547 5321 48559 5355
rect 48501 5315 48559 5321
rect 54297 5355 54355 5361
rect 54297 5321 54309 5355
rect 54343 5352 54355 5355
rect 55030 5352 55036 5364
rect 54343 5324 55036 5352
rect 54343 5321 54355 5324
rect 54297 5315 54355 5321
rect 55030 5312 55036 5324
rect 55088 5312 55094 5364
rect 62390 5352 62396 5364
rect 62351 5324 62396 5352
rect 62390 5312 62396 5324
rect 62448 5312 62454 5364
rect 63310 5352 63316 5364
rect 63271 5324 63316 5352
rect 63310 5312 63316 5324
rect 63368 5312 63374 5364
rect 65705 5355 65763 5361
rect 65705 5321 65717 5355
rect 65751 5352 65763 5355
rect 65886 5352 65892 5364
rect 65751 5324 65892 5352
rect 65751 5321 65763 5324
rect 65705 5315 65763 5321
rect 65886 5312 65892 5324
rect 65944 5312 65950 5364
rect 73154 5312 73160 5364
rect 73212 5352 73218 5364
rect 73525 5355 73583 5361
rect 73525 5352 73537 5355
rect 73212 5324 73537 5352
rect 73212 5312 73218 5324
rect 73525 5321 73537 5324
rect 73571 5352 73583 5355
rect 74350 5352 74356 5364
rect 73571 5324 74356 5352
rect 73571 5321 73583 5324
rect 73525 5315 73583 5321
rect 74350 5312 74356 5324
rect 74408 5312 74414 5364
rect 75914 5352 75920 5364
rect 75875 5324 75920 5352
rect 75914 5312 75920 5324
rect 75972 5312 75978 5364
rect 114094 5352 114100 5364
rect 76116 5324 114100 5352
rect 32306 5284 32312 5296
rect 24627 5256 27292 5284
rect 27356 5256 32312 5284
rect 24627 5253 24639 5256
rect 24581 5247 24639 5253
rect 21284 5188 24164 5216
rect 19705 5179 19763 5185
rect 15562 5148 15568 5160
rect 13688 5120 15148 5148
rect 15212 5120 15568 5148
rect 13688 5108 13694 5120
rect 5721 5083 5779 5089
rect 5721 5049 5733 5083
rect 5767 5080 5779 5083
rect 5767 5052 9076 5080
rect 5767 5049 5779 5052
rect 5721 5043 5779 5049
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 9048 5012 9076 5052
rect 12618 5012 12624 5024
rect 9048 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 14332 4984 14565 5012
rect 14332 4972 14338 4984
rect 14553 4981 14565 4984
rect 14599 5012 14611 5015
rect 14918 5012 14924 5024
rect 14599 4984 14924 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15120 5012 15148 5120
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 22462 5148 22468 5160
rect 15896 5120 22468 5148
rect 15896 5108 15902 5120
rect 22462 5108 22468 5120
rect 22520 5108 22526 5160
rect 22741 5151 22799 5157
rect 22741 5117 22753 5151
rect 22787 5117 22799 5151
rect 24136 5148 24164 5188
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 26145 5219 26203 5225
rect 26145 5216 26157 5219
rect 24728 5188 26157 5216
rect 24728 5176 24734 5188
rect 26145 5185 26157 5188
rect 26191 5216 26203 5219
rect 27356 5216 27384 5256
rect 32306 5244 32312 5256
rect 32364 5244 32370 5296
rect 33778 5244 33784 5296
rect 33836 5284 33842 5296
rect 34885 5287 34943 5293
rect 34885 5284 34897 5287
rect 33836 5256 34897 5284
rect 33836 5244 33842 5256
rect 34885 5253 34897 5256
rect 34931 5284 34943 5287
rect 45370 5284 45376 5296
rect 34931 5256 36768 5284
rect 45283 5256 45376 5284
rect 34931 5253 34943 5256
rect 34885 5247 34943 5253
rect 29650 5219 29708 5225
rect 29650 5216 29662 5219
rect 26191 5188 27384 5216
rect 27417 5188 29662 5216
rect 26191 5185 26203 5188
rect 26145 5179 26203 5185
rect 27417 5148 27445 5188
rect 29650 5185 29662 5188
rect 29696 5185 29708 5219
rect 29650 5179 29708 5185
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 31490 5219 31548 5225
rect 31490 5216 31502 5219
rect 30524 5188 31502 5216
rect 30524 5176 30530 5188
rect 31490 5185 31502 5188
rect 31536 5185 31548 5219
rect 31490 5179 31548 5185
rect 34241 5219 34299 5225
rect 34241 5185 34253 5219
rect 34287 5216 34299 5219
rect 35986 5216 35992 5228
rect 34287 5188 35992 5216
rect 34287 5185 34299 5188
rect 34241 5179 34299 5185
rect 35986 5176 35992 5188
rect 36044 5176 36050 5228
rect 36469 5219 36527 5225
rect 36469 5185 36481 5219
rect 36515 5216 36527 5219
rect 36630 5216 36636 5228
rect 36515 5188 36636 5216
rect 36515 5185 36527 5188
rect 36469 5179 36527 5185
rect 36630 5176 36636 5188
rect 36688 5176 36694 5228
rect 36740 5225 36768 5256
rect 45370 5244 45376 5256
rect 45428 5284 45434 5296
rect 45830 5284 45836 5296
rect 45428 5256 45836 5284
rect 45428 5244 45434 5256
rect 45830 5244 45836 5256
rect 45888 5244 45894 5296
rect 48314 5244 48320 5296
rect 48372 5284 48378 5296
rect 55646 5287 55704 5293
rect 55646 5284 55658 5287
rect 48372 5256 55658 5284
rect 48372 5244 48378 5256
rect 55646 5253 55658 5256
rect 55692 5253 55704 5287
rect 63328 5284 63356 5312
rect 55646 5247 55704 5253
rect 61028 5256 63356 5284
rect 36725 5219 36783 5225
rect 36725 5185 36737 5219
rect 36771 5216 36783 5219
rect 38562 5216 38568 5228
rect 36771 5188 38568 5216
rect 36771 5185 36783 5188
rect 36725 5179 36783 5185
rect 38562 5176 38568 5188
rect 38620 5176 38626 5228
rect 48682 5216 48688 5228
rect 48643 5188 48688 5216
rect 48682 5176 48688 5188
rect 48740 5176 48746 5228
rect 53184 5219 53242 5225
rect 53184 5185 53196 5219
rect 53230 5216 53242 5219
rect 58802 5216 58808 5228
rect 53230 5188 58808 5216
rect 53230 5185 53242 5188
rect 53184 5179 53242 5185
rect 58802 5176 58808 5188
rect 58860 5176 58866 5228
rect 61028 5225 61056 5256
rect 63586 5244 63592 5296
rect 63644 5284 63650 5296
rect 74997 5287 75055 5293
rect 63644 5256 74948 5284
rect 63644 5244 63650 5256
rect 61013 5219 61071 5225
rect 61013 5185 61025 5219
rect 61059 5185 61071 5219
rect 61013 5179 61071 5185
rect 61102 5176 61108 5228
rect 61160 5216 61166 5228
rect 61269 5219 61327 5225
rect 61269 5216 61281 5219
rect 61160 5188 61281 5216
rect 61160 5176 61166 5188
rect 61269 5185 61281 5188
rect 61315 5185 61327 5219
rect 61269 5179 61327 5185
rect 61746 5176 61752 5228
rect 61804 5216 61810 5228
rect 74810 5216 74816 5228
rect 61804 5188 74816 5216
rect 61804 5176 61810 5188
rect 74810 5176 74816 5188
rect 74868 5176 74874 5228
rect 74920 5216 74948 5256
rect 74997 5253 75009 5287
rect 75043 5284 75055 5287
rect 76006 5284 76012 5296
rect 75043 5256 76012 5284
rect 75043 5253 75055 5256
rect 74997 5247 75055 5253
rect 76006 5244 76012 5256
rect 76064 5244 76070 5296
rect 76116 5216 76144 5324
rect 114094 5312 114100 5324
rect 114152 5312 114158 5364
rect 115661 5355 115719 5361
rect 115661 5321 115673 5355
rect 115707 5352 115719 5355
rect 116026 5352 116032 5364
rect 115707 5324 116032 5352
rect 115707 5321 115719 5324
rect 115661 5315 115719 5321
rect 116026 5312 116032 5324
rect 116084 5312 116090 5364
rect 116305 5355 116363 5361
rect 116305 5321 116317 5355
rect 116351 5352 116363 5355
rect 118418 5352 118424 5364
rect 116351 5324 118424 5352
rect 116351 5321 116363 5324
rect 116305 5315 116363 5321
rect 118418 5312 118424 5324
rect 118476 5312 118482 5364
rect 118513 5355 118571 5361
rect 118513 5321 118525 5355
rect 118559 5352 118571 5355
rect 118694 5352 118700 5364
rect 118559 5324 118700 5352
rect 118559 5321 118571 5324
rect 118513 5315 118571 5321
rect 118694 5312 118700 5324
rect 118752 5312 118758 5364
rect 118878 5312 118884 5364
rect 118936 5352 118942 5364
rect 121273 5355 121331 5361
rect 121273 5352 121285 5355
rect 118936 5324 121285 5352
rect 118936 5312 118942 5324
rect 121273 5321 121285 5324
rect 121319 5352 121331 5355
rect 122650 5352 122656 5364
rect 121319 5324 122656 5352
rect 121319 5321 121331 5324
rect 121273 5315 121331 5321
rect 122650 5312 122656 5324
rect 122708 5312 122714 5364
rect 123110 5352 123116 5364
rect 123071 5324 123116 5352
rect 123110 5312 123116 5324
rect 123168 5312 123174 5364
rect 124493 5355 124551 5361
rect 124493 5321 124505 5355
rect 124539 5352 124551 5355
rect 125502 5352 125508 5364
rect 124539 5324 125508 5352
rect 124539 5321 124551 5324
rect 124493 5315 124551 5321
rect 125502 5312 125508 5324
rect 125560 5312 125566 5364
rect 126790 5312 126796 5364
rect 126848 5352 126854 5364
rect 127713 5355 127771 5361
rect 127713 5352 127725 5355
rect 126848 5324 127725 5352
rect 126848 5312 126854 5324
rect 127713 5321 127725 5324
rect 127759 5321 127771 5355
rect 127713 5315 127771 5321
rect 127802 5312 127808 5364
rect 127860 5352 127866 5364
rect 128078 5352 128084 5364
rect 127860 5324 128084 5352
rect 127860 5312 127866 5324
rect 128078 5312 128084 5324
rect 128136 5312 128142 5364
rect 128354 5312 128360 5364
rect 128412 5352 128418 5364
rect 129093 5355 129151 5361
rect 129093 5352 129105 5355
rect 128412 5324 129105 5352
rect 128412 5312 128418 5324
rect 129093 5321 129105 5324
rect 129139 5352 129151 5355
rect 129182 5352 129188 5364
rect 129139 5324 129188 5352
rect 129139 5321 129151 5324
rect 129093 5315 129151 5321
rect 129182 5312 129188 5324
rect 129240 5312 129246 5364
rect 129645 5355 129703 5361
rect 129645 5321 129657 5355
rect 129691 5352 129703 5355
rect 129734 5352 129740 5364
rect 129691 5324 129740 5352
rect 129691 5321 129703 5324
rect 129645 5315 129703 5321
rect 129734 5312 129740 5324
rect 129792 5312 129798 5364
rect 129826 5312 129832 5364
rect 129884 5352 129890 5364
rect 137370 5352 137376 5364
rect 129884 5324 137376 5352
rect 129884 5312 129890 5324
rect 137370 5312 137376 5324
rect 137428 5312 137434 5364
rect 137830 5352 137836 5364
rect 137791 5324 137836 5352
rect 137830 5312 137836 5324
rect 137888 5312 137894 5364
rect 138382 5352 138388 5364
rect 138343 5324 138388 5352
rect 138382 5312 138388 5324
rect 138440 5312 138446 5364
rect 139302 5352 139308 5364
rect 139263 5324 139308 5352
rect 139302 5312 139308 5324
rect 139360 5312 139366 5364
rect 139949 5355 140007 5361
rect 139949 5321 139961 5355
rect 139995 5352 140007 5355
rect 141510 5352 141516 5364
rect 139995 5324 141516 5352
rect 139995 5321 140007 5324
rect 139949 5315 140007 5321
rect 141510 5312 141516 5324
rect 141568 5312 141574 5364
rect 142706 5312 142712 5364
rect 142764 5352 142770 5364
rect 144638 5352 144644 5364
rect 142764 5324 143948 5352
rect 144599 5324 144644 5352
rect 142764 5312 142770 5324
rect 77205 5287 77263 5293
rect 77205 5253 77217 5287
rect 77251 5284 77263 5287
rect 81250 5284 81256 5296
rect 77251 5256 81256 5284
rect 77251 5253 77263 5256
rect 77205 5247 77263 5253
rect 81250 5244 81256 5256
rect 81308 5244 81314 5296
rect 93394 5284 93400 5296
rect 90744 5256 93400 5284
rect 74920 5188 76144 5216
rect 79045 5219 79103 5225
rect 79045 5185 79057 5219
rect 79091 5216 79103 5219
rect 81066 5216 81072 5228
rect 79091 5188 81072 5216
rect 79091 5185 79103 5188
rect 79045 5179 79103 5185
rect 81066 5176 81072 5188
rect 81124 5176 81130 5228
rect 82541 5219 82599 5225
rect 82541 5216 82553 5219
rect 81268 5188 82553 5216
rect 24136 5120 27445 5148
rect 29917 5151 29975 5157
rect 22741 5111 22799 5117
rect 29917 5117 29929 5151
rect 29963 5148 29975 5151
rect 30282 5148 30288 5160
rect 29963 5120 30288 5148
rect 29963 5117 29975 5120
rect 29917 5111 29975 5117
rect 15381 5083 15439 5089
rect 15381 5049 15393 5083
rect 15427 5080 15439 5083
rect 17218 5080 17224 5092
rect 15427 5052 17224 5080
rect 15427 5049 15439 5052
rect 15381 5043 15439 5049
rect 17218 5040 17224 5052
rect 17276 5040 17282 5092
rect 21910 5080 21916 5092
rect 17328 5052 21916 5080
rect 17328 5012 17356 5052
rect 21910 5040 21916 5052
rect 21968 5040 21974 5092
rect 22554 5040 22560 5092
rect 22612 5080 22618 5092
rect 22756 5080 22784 5111
rect 30282 5108 30288 5120
rect 30340 5108 30346 5160
rect 31754 5108 31760 5160
rect 31812 5148 31818 5160
rect 34330 5148 34336 5160
rect 31812 5120 34336 5148
rect 31812 5108 31818 5120
rect 34330 5108 34336 5120
rect 34388 5108 34394 5160
rect 51074 5108 51080 5160
rect 51132 5148 51138 5160
rect 52270 5148 52276 5160
rect 51132 5120 52276 5148
rect 51132 5108 51138 5120
rect 52270 5108 52276 5120
rect 52328 5148 52334 5160
rect 52917 5151 52975 5157
rect 52917 5148 52929 5151
rect 52328 5120 52929 5148
rect 52328 5108 52334 5120
rect 52917 5117 52929 5120
rect 52963 5117 52975 5151
rect 55398 5148 55404 5160
rect 55311 5120 55404 5148
rect 52917 5111 52975 5117
rect 34054 5080 34060 5092
rect 22612 5052 22784 5080
rect 34015 5052 34060 5080
rect 22612 5040 22618 5052
rect 15120 4984 17356 5012
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 22646 5012 22652 5024
rect 18288 4984 22652 5012
rect 18288 4972 18294 4984
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 22756 5012 22784 5052
rect 34054 5040 34060 5052
rect 34112 5040 34118 5092
rect 24670 5012 24676 5024
rect 22756 4984 24676 5012
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 25314 4972 25320 5024
rect 25372 5012 25378 5024
rect 28537 5015 28595 5021
rect 28537 5012 28549 5015
rect 25372 4984 28549 5012
rect 25372 4972 25378 4984
rect 28537 4981 28549 4984
rect 28583 4981 28595 5015
rect 30374 5012 30380 5024
rect 30335 4984 30380 5012
rect 28537 4975 28595 4981
rect 30374 4972 30380 4984
rect 30432 4972 30438 5024
rect 52932 5012 52960 5111
rect 55398 5108 55404 5120
rect 55456 5108 55462 5160
rect 75546 5108 75552 5160
rect 75604 5148 75610 5160
rect 81268 5148 81296 5188
rect 82541 5185 82553 5188
rect 82587 5185 82599 5219
rect 82541 5179 82599 5185
rect 88334 5176 88340 5228
rect 88392 5216 88398 5228
rect 90744 5225 90772 5256
rect 90729 5219 90787 5225
rect 90729 5216 90741 5219
rect 88392 5188 90741 5216
rect 88392 5176 88398 5188
rect 90729 5185 90741 5188
rect 90775 5185 90787 5219
rect 90729 5179 90787 5185
rect 92405 5219 92463 5225
rect 92405 5185 92417 5219
rect 92451 5216 92463 5219
rect 92566 5216 92572 5228
rect 92451 5188 92572 5216
rect 92451 5185 92463 5188
rect 92405 5179 92463 5185
rect 92566 5176 92572 5188
rect 92624 5176 92630 5228
rect 92676 5225 92704 5256
rect 93394 5244 93400 5256
rect 93452 5284 93458 5296
rect 95326 5284 95332 5296
rect 93452 5256 95332 5284
rect 93452 5244 93458 5256
rect 95326 5244 95332 5256
rect 95384 5244 95390 5296
rect 104888 5287 104946 5293
rect 104888 5253 104900 5287
rect 104934 5284 104946 5287
rect 106553 5287 106611 5293
rect 106553 5284 106565 5287
rect 104934 5256 106565 5284
rect 104934 5253 104946 5256
rect 104888 5247 104946 5253
rect 106553 5253 106565 5256
rect 106599 5284 106611 5287
rect 116946 5284 116952 5296
rect 106599 5256 116952 5284
rect 106599 5253 106611 5256
rect 106553 5247 106611 5253
rect 116946 5244 116952 5256
rect 117004 5244 117010 5296
rect 117130 5244 117136 5296
rect 117188 5284 117194 5296
rect 120166 5293 120172 5296
rect 120160 5284 120172 5293
rect 117188 5256 119936 5284
rect 120127 5256 120172 5284
rect 117188 5244 117194 5256
rect 92661 5219 92719 5225
rect 92661 5185 92673 5219
rect 92707 5185 92719 5219
rect 93118 5216 93124 5228
rect 93079 5188 93124 5216
rect 92661 5179 92719 5185
rect 93118 5176 93124 5188
rect 93176 5176 93182 5228
rect 93210 5176 93216 5228
rect 93268 5216 93274 5228
rect 96706 5216 96712 5228
rect 93268 5188 96712 5216
rect 93268 5176 93274 5188
rect 96706 5176 96712 5188
rect 96764 5176 96770 5228
rect 105170 5176 105176 5228
rect 105228 5216 105234 5228
rect 109126 5216 109132 5228
rect 105228 5188 109132 5216
rect 105228 5176 105234 5188
rect 109126 5176 109132 5188
rect 109184 5216 109190 5228
rect 109770 5216 109776 5228
rect 109184 5188 109776 5216
rect 109184 5176 109190 5188
rect 109770 5176 109776 5188
rect 109828 5176 109834 5228
rect 112349 5219 112407 5225
rect 112349 5185 112361 5219
rect 112395 5216 112407 5219
rect 113818 5216 113824 5228
rect 112395 5188 113824 5216
rect 112395 5185 112407 5188
rect 112349 5179 112407 5185
rect 113818 5176 113824 5188
rect 113876 5176 113882 5228
rect 114925 5219 114983 5225
rect 114925 5216 114937 5219
rect 114112 5188 114937 5216
rect 82357 5151 82415 5157
rect 82357 5148 82369 5151
rect 75604 5120 81296 5148
rect 81912 5120 82369 5148
rect 75604 5108 75610 5120
rect 55416 5012 55444 5108
rect 77202 5040 77208 5092
rect 77260 5080 77266 5092
rect 78861 5083 78919 5089
rect 78861 5080 78873 5083
rect 77260 5052 78873 5080
rect 77260 5040 77266 5052
rect 78861 5049 78873 5052
rect 78907 5049 78919 5083
rect 78861 5043 78919 5049
rect 81912 5024 81940 5120
rect 82357 5117 82369 5120
rect 82403 5148 82415 5151
rect 82998 5148 83004 5160
rect 82403 5120 83004 5148
rect 82403 5117 82415 5120
rect 82357 5111 82415 5117
rect 82998 5108 83004 5120
rect 83056 5108 83062 5160
rect 101306 5108 101312 5160
rect 101364 5148 101370 5160
rect 104618 5148 104624 5160
rect 101364 5120 104624 5148
rect 101364 5108 101370 5120
rect 104618 5108 104624 5120
rect 104676 5108 104682 5160
rect 110874 5108 110880 5160
rect 110932 5148 110938 5160
rect 110932 5120 112392 5148
rect 110932 5108 110938 5120
rect 88058 5040 88064 5092
rect 88116 5080 88122 5092
rect 93305 5083 93363 5089
rect 88116 5052 91416 5080
rect 88116 5040 88122 5052
rect 56778 5012 56784 5024
rect 52932 4984 55444 5012
rect 56739 4984 56784 5012
rect 56778 4972 56784 4984
rect 56836 4972 56842 5024
rect 81894 5012 81900 5024
rect 81855 4984 81900 5012
rect 81894 4972 81900 4984
rect 81952 4972 81958 5024
rect 82725 5015 82783 5021
rect 82725 4981 82737 5015
rect 82771 5012 82783 5015
rect 84286 5012 84292 5024
rect 82771 4984 84292 5012
rect 82771 4981 82783 4984
rect 82725 4975 82783 4981
rect 84286 4972 84292 4984
rect 84344 4972 84350 5024
rect 91094 4972 91100 5024
rect 91152 5012 91158 5024
rect 91281 5015 91339 5021
rect 91281 5012 91293 5015
rect 91152 4984 91293 5012
rect 91152 4972 91158 4984
rect 91281 4981 91293 4984
rect 91327 4981 91339 5015
rect 91388 5012 91416 5052
rect 93305 5049 93317 5083
rect 93351 5080 93363 5083
rect 94130 5080 94136 5092
rect 93351 5052 94136 5080
rect 93351 5049 93363 5052
rect 93305 5043 93363 5049
rect 94130 5040 94136 5052
rect 94188 5040 94194 5092
rect 111886 5080 111892 5092
rect 106016 5052 111892 5080
rect 106016 5021 106044 5052
rect 111886 5040 111892 5052
rect 111944 5040 111950 5092
rect 112364 5080 112392 5120
rect 113542 5108 113548 5160
rect 113600 5148 113606 5160
rect 114112 5157 114140 5188
rect 114925 5185 114937 5188
rect 114971 5185 114983 5219
rect 114925 5179 114983 5185
rect 117429 5219 117487 5225
rect 117429 5185 117441 5219
rect 117475 5216 117487 5219
rect 118050 5216 118056 5228
rect 117475 5188 118056 5216
rect 117475 5185 117487 5188
rect 117429 5179 117487 5185
rect 118050 5176 118056 5188
rect 118108 5176 118114 5228
rect 118326 5176 118332 5228
rect 118384 5216 118390 5228
rect 119908 5225 119936 5256
rect 120160 5247 120172 5256
rect 120166 5244 120172 5247
rect 120224 5244 120230 5296
rect 121822 5244 121828 5296
rect 121880 5284 121886 5296
rect 123849 5287 123907 5293
rect 123849 5284 123861 5287
rect 121880 5256 123861 5284
rect 121880 5244 121886 5256
rect 123849 5253 123861 5256
rect 123895 5284 123907 5287
rect 125042 5284 125048 5296
rect 123895 5256 125048 5284
rect 123895 5253 123907 5256
rect 123849 5247 123907 5253
rect 125042 5244 125048 5256
rect 125100 5284 125106 5296
rect 127066 5284 127072 5296
rect 125100 5256 127072 5284
rect 125100 5244 125106 5256
rect 127066 5244 127072 5256
rect 127124 5284 127130 5296
rect 132034 5284 132040 5296
rect 127124 5256 131528 5284
rect 131995 5256 132040 5284
rect 127124 5244 127130 5256
rect 131500 5228 131528 5256
rect 132034 5244 132040 5256
rect 132092 5284 132098 5296
rect 137186 5284 137192 5296
rect 132092 5256 137192 5284
rect 132092 5244 132098 5256
rect 137186 5244 137192 5256
rect 137244 5244 137250 5296
rect 137278 5244 137284 5296
rect 137336 5284 137342 5296
rect 137557 5287 137615 5293
rect 137557 5284 137569 5287
rect 137336 5256 137569 5284
rect 137336 5244 137342 5256
rect 137557 5253 137569 5256
rect 137603 5253 137615 5287
rect 140222 5284 140228 5296
rect 137557 5247 137615 5253
rect 138400 5256 140228 5284
rect 118697 5219 118755 5225
rect 118697 5216 118709 5219
rect 118384 5188 118709 5216
rect 118384 5176 118390 5188
rect 118697 5185 118709 5188
rect 118743 5185 118755 5219
rect 118697 5179 118755 5185
rect 119893 5219 119951 5225
rect 119893 5185 119905 5219
rect 119939 5185 119951 5219
rect 121989 5219 122047 5225
rect 121989 5216 122001 5219
rect 119893 5179 119951 5185
rect 120000 5188 122001 5216
rect 114097 5151 114155 5157
rect 114097 5148 114109 5151
rect 113600 5120 114109 5148
rect 113600 5108 113606 5120
rect 114097 5117 114109 5120
rect 114143 5117 114155 5151
rect 114097 5111 114155 5117
rect 114741 5151 114799 5157
rect 114741 5117 114753 5151
rect 114787 5148 114799 5151
rect 116026 5148 116032 5160
rect 114787 5120 116032 5148
rect 114787 5117 114799 5120
rect 114741 5111 114799 5117
rect 116026 5108 116032 5120
rect 116084 5108 116090 5160
rect 117685 5151 117743 5157
rect 117685 5117 117697 5151
rect 117731 5148 117743 5151
rect 117774 5148 117780 5160
rect 117731 5120 117780 5148
rect 117731 5117 117743 5120
rect 117685 5111 117743 5117
rect 117774 5108 117780 5120
rect 117832 5108 117838 5160
rect 117866 5108 117872 5160
rect 117924 5148 117930 5160
rect 120000 5148 120028 5188
rect 121989 5185 122001 5188
rect 122035 5185 122047 5219
rect 121989 5179 122047 5185
rect 124214 5176 124220 5228
rect 124272 5216 124278 5228
rect 125321 5219 125379 5225
rect 125321 5216 125333 5219
rect 124272 5188 125333 5216
rect 124272 5176 124278 5188
rect 125321 5185 125333 5188
rect 125367 5185 125379 5219
rect 125321 5179 125379 5185
rect 126698 5176 126704 5228
rect 126756 5216 126762 5228
rect 127158 5216 127164 5228
rect 126756 5188 127020 5216
rect 127119 5188 127164 5216
rect 126756 5176 126762 5188
rect 121730 5148 121736 5160
rect 117924 5120 120028 5148
rect 121691 5120 121736 5148
rect 117924 5108 117930 5120
rect 121730 5108 121736 5120
rect 121788 5108 121794 5160
rect 125042 5148 125048 5160
rect 125003 5120 125048 5148
rect 125042 5108 125048 5120
rect 125100 5108 125106 5160
rect 125134 5108 125140 5160
rect 125192 5148 125198 5160
rect 126992 5148 127020 5188
rect 127158 5176 127164 5188
rect 127216 5216 127222 5228
rect 127897 5219 127955 5225
rect 127897 5216 127909 5219
rect 127216 5188 127909 5216
rect 127216 5176 127222 5188
rect 127897 5185 127909 5188
rect 127943 5185 127955 5219
rect 128078 5216 128084 5228
rect 128039 5188 128084 5216
rect 127897 5179 127955 5185
rect 128078 5176 128084 5188
rect 128136 5176 128142 5228
rect 131390 5216 131396 5228
rect 131351 5188 131396 5216
rect 131390 5176 131396 5188
rect 131448 5176 131454 5228
rect 131482 5176 131488 5228
rect 131540 5216 131546 5228
rect 134794 5216 134800 5228
rect 131540 5188 134800 5216
rect 131540 5176 131546 5188
rect 134794 5176 134800 5188
rect 134852 5176 134858 5228
rect 136818 5216 136824 5228
rect 136779 5188 136824 5216
rect 136818 5176 136824 5188
rect 136876 5176 136882 5228
rect 136910 5176 136916 5228
rect 136968 5216 136974 5228
rect 138400 5216 138428 5256
rect 140222 5244 140228 5256
rect 140280 5284 140286 5296
rect 140280 5256 141924 5284
rect 140280 5244 140286 5256
rect 138566 5216 138572 5228
rect 136968 5188 138428 5216
rect 138527 5188 138572 5216
rect 136968 5176 136974 5188
rect 138566 5176 138572 5188
rect 138624 5176 138630 5228
rect 139762 5216 139768 5228
rect 139723 5188 139768 5216
rect 139762 5176 139768 5188
rect 139820 5176 139826 5228
rect 139854 5176 139860 5228
rect 139912 5216 139918 5228
rect 140038 5216 140044 5228
rect 139912 5188 140044 5216
rect 139912 5176 139918 5188
rect 140038 5176 140044 5188
rect 140096 5176 140102 5228
rect 141142 5176 141148 5228
rect 141200 5216 141206 5228
rect 141706 5219 141764 5225
rect 141706 5216 141718 5219
rect 141200 5188 141718 5216
rect 141200 5176 141206 5188
rect 141706 5185 141718 5188
rect 141752 5185 141764 5219
rect 141706 5179 141764 5185
rect 127986 5148 127992 5160
rect 125192 5120 126744 5148
rect 126992 5120 127992 5148
rect 125192 5108 125198 5120
rect 115842 5080 115848 5092
rect 112364 5052 115848 5080
rect 115842 5040 115848 5052
rect 115900 5040 115906 5092
rect 118142 5040 118148 5092
rect 118200 5080 118206 5092
rect 119062 5080 119068 5092
rect 118200 5052 119068 5080
rect 118200 5040 118206 5052
rect 119062 5040 119068 5052
rect 119120 5040 119126 5092
rect 122834 5040 122840 5092
rect 122892 5080 122898 5092
rect 125870 5080 125876 5092
rect 122892 5052 125876 5080
rect 122892 5040 122898 5052
rect 125870 5040 125876 5052
rect 125928 5040 125934 5092
rect 106001 5015 106059 5021
rect 106001 5012 106013 5015
rect 91388 4984 106013 5012
rect 91281 4975 91339 4981
rect 106001 4981 106013 4984
rect 106047 4981 106059 5015
rect 112162 5012 112168 5024
rect 112123 4984 112168 5012
rect 106001 4975 106059 4981
rect 112162 4972 112168 4984
rect 112220 4972 112226 5024
rect 115109 5015 115167 5021
rect 115109 4981 115121 5015
rect 115155 5012 115167 5015
rect 115474 5012 115480 5024
rect 115155 4984 115480 5012
rect 115155 4981 115167 4984
rect 115109 4975 115167 4981
rect 115474 4972 115480 4984
rect 115532 4972 115538 5024
rect 119246 5012 119252 5024
rect 119207 4984 119252 5012
rect 119246 4972 119252 4984
rect 119304 4972 119310 5024
rect 124030 4972 124036 5024
rect 124088 5012 124094 5024
rect 125410 5012 125416 5024
rect 124088 4984 125416 5012
rect 124088 4972 124094 4984
rect 125410 4972 125416 4984
rect 125468 4972 125474 5024
rect 126514 4972 126520 5024
rect 126572 5012 126578 5024
rect 126609 5015 126667 5021
rect 126609 5012 126621 5015
rect 126572 4984 126621 5012
rect 126572 4972 126578 4984
rect 126609 4981 126621 4984
rect 126655 4981 126667 5015
rect 126716 5012 126744 5120
rect 127986 5108 127992 5120
rect 128044 5108 128050 5160
rect 129734 5148 129740 5160
rect 128326 5120 129740 5148
rect 126790 5040 126796 5092
rect 126848 5080 126854 5092
rect 128326 5080 128354 5120
rect 129734 5108 129740 5120
rect 129792 5108 129798 5160
rect 131408 5148 131436 5176
rect 131666 5148 131672 5160
rect 131408 5120 131672 5148
rect 131666 5108 131672 5120
rect 131724 5108 131730 5160
rect 132494 5108 132500 5160
rect 132552 5148 132558 5160
rect 133601 5151 133659 5157
rect 133601 5148 133613 5151
rect 132552 5120 133613 5148
rect 132552 5108 132558 5120
rect 133601 5117 133613 5120
rect 133647 5117 133659 5151
rect 140958 5148 140964 5160
rect 133601 5111 133659 5117
rect 133708 5120 140964 5148
rect 130381 5083 130439 5089
rect 130381 5080 130393 5083
rect 126848 5052 128354 5080
rect 128924 5052 130393 5080
rect 126848 5040 126854 5052
rect 128924 5012 128952 5052
rect 130381 5049 130393 5052
rect 130427 5080 130439 5083
rect 133708 5080 133736 5120
rect 140958 5108 140964 5120
rect 141016 5108 141022 5160
rect 141896 5148 141924 5256
rect 142798 5244 142804 5296
rect 142856 5284 142862 5296
rect 142856 5256 143856 5284
rect 142856 5244 142862 5256
rect 141973 5219 142031 5225
rect 141973 5185 141985 5219
rect 142019 5216 142031 5219
rect 142338 5216 142344 5228
rect 142019 5188 142344 5216
rect 142019 5185 142031 5188
rect 141973 5179 142031 5185
rect 142338 5176 142344 5188
rect 142396 5176 142402 5228
rect 143828 5225 143856 5256
rect 143557 5219 143615 5225
rect 143557 5185 143569 5219
rect 143603 5216 143615 5219
rect 143813 5219 143871 5225
rect 143603 5188 143764 5216
rect 143603 5185 143615 5188
rect 143557 5179 143615 5185
rect 143736 5148 143764 5188
rect 143813 5185 143825 5219
rect 143859 5185 143871 5219
rect 143920 5216 143948 5324
rect 144638 5312 144644 5324
rect 144696 5312 144702 5364
rect 145558 5312 145564 5364
rect 145616 5352 145622 5364
rect 145653 5355 145711 5361
rect 145653 5352 145665 5355
rect 145616 5324 145665 5352
rect 145616 5312 145622 5324
rect 145653 5321 145665 5324
rect 145699 5321 145711 5355
rect 145653 5315 145711 5321
rect 146754 5312 146760 5364
rect 146812 5352 146818 5364
rect 147582 5352 147588 5364
rect 146812 5324 147588 5352
rect 146812 5312 146818 5324
rect 147582 5312 147588 5324
rect 147640 5352 147646 5364
rect 153013 5355 153071 5361
rect 147640 5324 151961 5352
rect 147640 5312 147646 5324
rect 144178 5244 144184 5296
rect 144236 5284 144242 5296
rect 147306 5284 147312 5296
rect 144236 5256 147312 5284
rect 144236 5244 144242 5256
rect 147306 5244 147312 5256
rect 147364 5244 147370 5296
rect 147674 5244 147680 5296
rect 147732 5284 147738 5296
rect 150250 5284 150256 5296
rect 147732 5256 150256 5284
rect 147732 5244 147738 5256
rect 150250 5244 150256 5256
rect 150308 5244 150314 5296
rect 150342 5244 150348 5296
rect 150400 5284 150406 5296
rect 151814 5284 151820 5296
rect 150400 5256 151820 5284
rect 150400 5244 150406 5256
rect 151814 5244 151820 5256
rect 151872 5244 151878 5296
rect 151933 5293 151961 5324
rect 153013 5321 153025 5355
rect 153059 5352 153071 5355
rect 155862 5352 155868 5364
rect 153059 5324 155868 5352
rect 153059 5321 153071 5324
rect 153013 5315 153071 5321
rect 155862 5312 155868 5324
rect 155920 5312 155926 5364
rect 156782 5352 156788 5364
rect 156743 5324 156788 5352
rect 156782 5312 156788 5324
rect 156840 5312 156846 5364
rect 157150 5312 157156 5364
rect 157208 5352 157214 5364
rect 158073 5355 158131 5361
rect 158073 5352 158085 5355
rect 157208 5324 158085 5352
rect 157208 5312 157214 5324
rect 158073 5321 158085 5324
rect 158119 5321 158131 5355
rect 158073 5315 158131 5321
rect 151918 5287 151976 5293
rect 151918 5253 151930 5287
rect 151964 5253 151976 5287
rect 154298 5284 154304 5296
rect 151918 5247 151976 5253
rect 152016 5256 154304 5284
rect 144805 5219 144863 5225
rect 144805 5216 144817 5219
rect 143920 5188 144817 5216
rect 143813 5179 143871 5185
rect 144805 5185 144817 5188
rect 144851 5185 144863 5219
rect 144805 5179 144863 5185
rect 145009 5219 145067 5225
rect 145009 5185 145021 5219
rect 145055 5216 145067 5219
rect 145282 5216 145288 5228
rect 145055 5188 145288 5216
rect 145055 5185 145067 5188
rect 145009 5179 145067 5185
rect 145282 5176 145288 5188
rect 145340 5176 145346 5228
rect 146777 5219 146835 5225
rect 146777 5185 146789 5219
rect 146823 5216 146835 5219
rect 146938 5216 146944 5228
rect 146823 5188 146944 5216
rect 146823 5185 146835 5188
rect 146777 5179 146835 5185
rect 146938 5176 146944 5188
rect 146996 5176 147002 5228
rect 147030 5176 147036 5228
rect 147088 5216 147094 5228
rect 148606 5220 148664 5225
rect 148606 5219 148824 5220
rect 147088 5188 147133 5216
rect 147088 5176 147094 5188
rect 148606 5185 148618 5219
rect 148652 5192 148824 5219
rect 148652 5185 148664 5192
rect 148606 5179 148664 5185
rect 145926 5148 145932 5160
rect 141896 5120 142844 5148
rect 143736 5120 145932 5148
rect 135714 5080 135720 5092
rect 130427 5052 133736 5080
rect 134168 5052 135720 5080
rect 130427 5049 130439 5052
rect 130381 5043 130439 5049
rect 130838 5012 130844 5024
rect 126716 4984 128952 5012
rect 130799 4984 130844 5012
rect 126609 4975 126667 4981
rect 130838 4972 130844 4984
rect 130896 4972 130902 5024
rect 132310 4972 132316 5024
rect 132368 5012 132374 5024
rect 132497 5015 132555 5021
rect 132497 5012 132509 5015
rect 132368 4984 132509 5012
rect 132368 4972 132374 4984
rect 132497 4981 132509 4984
rect 132543 4981 132555 5015
rect 133046 5012 133052 5024
rect 133007 4984 133052 5012
rect 132497 4975 132555 4981
rect 133046 4972 133052 4984
rect 133104 5012 133110 5024
rect 134168 5021 134196 5052
rect 135714 5040 135720 5052
rect 135772 5040 135778 5092
rect 140590 5080 140596 5092
rect 135916 5052 138014 5080
rect 140551 5052 140596 5080
rect 134153 5015 134211 5021
rect 134153 5012 134165 5015
rect 133104 4984 134165 5012
rect 133104 4972 133110 4984
rect 134153 4981 134165 4984
rect 134199 4981 134211 5015
rect 134794 5012 134800 5024
rect 134707 4984 134800 5012
rect 134153 4975 134211 4981
rect 134794 4972 134800 4984
rect 134852 5012 134858 5024
rect 135916 5012 135944 5052
rect 134852 4984 135944 5012
rect 136361 5015 136419 5021
rect 134852 4972 134858 4984
rect 136361 4981 136373 5015
rect 136407 5012 136419 5015
rect 136910 5012 136916 5024
rect 136407 4984 136916 5012
rect 136407 4981 136419 4984
rect 136361 4975 136419 4981
rect 136910 4972 136916 4984
rect 136968 4972 136974 5024
rect 137005 5015 137063 5021
rect 137005 4981 137017 5015
rect 137051 5012 137063 5015
rect 137554 5012 137560 5024
rect 137051 4984 137560 5012
rect 137051 4981 137063 4984
rect 137005 4975 137063 4981
rect 137554 4972 137560 4984
rect 137612 4972 137618 5024
rect 137986 5012 138014 5052
rect 140590 5040 140596 5052
rect 140648 5040 140654 5092
rect 139578 5012 139584 5024
rect 137986 4984 139584 5012
rect 139578 4972 139584 4984
rect 139636 4972 139642 5024
rect 139762 4972 139768 5024
rect 139820 5012 139826 5024
rect 142433 5015 142491 5021
rect 142433 5012 142445 5015
rect 139820 4984 142445 5012
rect 139820 4972 139826 4984
rect 142433 4981 142445 4984
rect 142479 5012 142491 5015
rect 142706 5012 142712 5024
rect 142479 4984 142712 5012
rect 142479 4981 142491 4984
rect 142433 4975 142491 4981
rect 142706 4972 142712 4984
rect 142764 4972 142770 5024
rect 142816 5012 142844 5120
rect 145926 5108 145932 5120
rect 145984 5108 145990 5160
rect 148796 5148 148824 5192
rect 148870 5176 148876 5228
rect 148928 5216 148934 5228
rect 148928 5188 148973 5216
rect 148928 5176 148934 5188
rect 149330 5176 149336 5228
rect 149388 5216 149394 5228
rect 149701 5219 149759 5225
rect 149701 5216 149713 5219
rect 149388 5188 149713 5216
rect 149388 5176 149394 5188
rect 149701 5185 149713 5188
rect 149747 5185 149759 5219
rect 149701 5179 149759 5185
rect 149790 5176 149796 5228
rect 149848 5216 149854 5228
rect 152016 5216 152044 5256
rect 154298 5244 154304 5256
rect 154356 5244 154362 5296
rect 154945 5287 155003 5293
rect 154546 5256 154896 5284
rect 149848 5188 152044 5216
rect 149848 5176 149854 5188
rect 152366 5176 152372 5228
rect 152424 5216 152430 5228
rect 152829 5219 152887 5225
rect 152829 5216 152841 5219
rect 152424 5188 152841 5216
rect 152424 5176 152430 5188
rect 152829 5185 152841 5188
rect 152875 5185 152887 5219
rect 152829 5179 152887 5185
rect 153657 5219 153715 5225
rect 153657 5185 153669 5219
rect 153703 5216 153715 5219
rect 154022 5216 154028 5228
rect 153703 5188 154028 5216
rect 153703 5185 153715 5188
rect 153657 5179 153715 5185
rect 154022 5176 154028 5188
rect 154080 5176 154086 5228
rect 148796 5120 151236 5148
rect 147122 5040 147128 5092
rect 147180 5080 147186 5092
rect 150342 5080 150348 5092
rect 147180 5052 147628 5080
rect 147180 5040 147186 5052
rect 145282 5012 145288 5024
rect 142816 4984 145288 5012
rect 145282 4972 145288 4984
rect 145340 4972 145346 5024
rect 145650 4972 145656 5024
rect 145708 5012 145714 5024
rect 147306 5012 147312 5024
rect 145708 4984 147312 5012
rect 145708 4972 145714 4984
rect 147306 4972 147312 4984
rect 147364 5012 147370 5024
rect 147493 5015 147551 5021
rect 147493 5012 147505 5015
rect 147364 4984 147505 5012
rect 147364 4972 147370 4984
rect 147493 4981 147505 4984
rect 147539 4981 147551 5015
rect 147600 5012 147628 5052
rect 148888 5052 150348 5080
rect 148888 5012 148916 5052
rect 150342 5040 150348 5052
rect 150400 5040 150406 5092
rect 147600 4984 148916 5012
rect 147493 4975 147551 4981
rect 149698 4972 149704 5024
rect 149756 5012 149762 5024
rect 149885 5015 149943 5021
rect 149885 5012 149897 5015
rect 149756 4984 149897 5012
rect 149756 4972 149762 4984
rect 149885 4981 149897 4984
rect 149931 4981 149943 5015
rect 150802 5012 150808 5024
rect 150763 4984 150808 5012
rect 149885 4975 149943 4981
rect 150802 4972 150808 4984
rect 150860 4972 150866 5024
rect 151208 5012 151236 5120
rect 152182 5108 152188 5160
rect 152240 5148 152246 5160
rect 152642 5148 152648 5160
rect 152240 5120 152333 5148
rect 152603 5120 152648 5148
rect 152240 5108 152246 5120
rect 152642 5108 152648 5120
rect 152700 5108 152706 5160
rect 153378 5108 153384 5160
rect 153436 5148 153442 5160
rect 154114 5148 154120 5160
rect 153436 5120 154120 5148
rect 153436 5108 153442 5120
rect 154114 5108 154120 5120
rect 154172 5148 154178 5160
rect 154546 5148 154574 5256
rect 154666 5216 154672 5228
rect 154627 5188 154672 5216
rect 154666 5176 154672 5188
rect 154724 5176 154730 5228
rect 154781 5219 154839 5225
rect 154781 5185 154793 5219
rect 154827 5216 154839 5219
rect 154868 5216 154896 5256
rect 154945 5253 154957 5287
rect 154991 5284 155003 5287
rect 159174 5284 159180 5296
rect 154991 5256 159180 5284
rect 154991 5253 155003 5256
rect 154945 5247 155003 5253
rect 159174 5244 159180 5256
rect 159232 5244 159238 5296
rect 154827 5188 154896 5216
rect 154827 5185 154839 5188
rect 154781 5179 154839 5185
rect 155770 5176 155776 5228
rect 155828 5216 155834 5228
rect 155957 5219 156015 5225
rect 155957 5216 155969 5219
rect 155828 5188 155969 5216
rect 155828 5176 155834 5188
rect 155957 5185 155969 5188
rect 156003 5185 156015 5219
rect 155957 5179 156015 5185
rect 156141 5219 156199 5225
rect 156141 5185 156153 5219
rect 156187 5185 156199 5219
rect 156141 5179 156199 5185
rect 154172 5120 154574 5148
rect 154172 5108 154178 5120
rect 152200 5080 152228 5108
rect 152550 5080 152556 5092
rect 152200 5052 152556 5080
rect 152550 5040 152556 5052
rect 152608 5040 152614 5092
rect 155310 5080 155316 5092
rect 152936 5052 155316 5080
rect 152936 5012 152964 5052
rect 155310 5040 155316 5052
rect 155368 5040 155374 5092
rect 155494 5040 155500 5092
rect 155552 5080 155558 5092
rect 156156 5080 156184 5179
rect 156598 5176 156604 5228
rect 156656 5216 156662 5228
rect 156969 5219 157027 5225
rect 156969 5216 156981 5219
rect 156656 5188 156981 5216
rect 156656 5176 156662 5188
rect 156969 5185 156981 5188
rect 157015 5185 157027 5219
rect 156969 5179 157027 5185
rect 157334 5176 157340 5228
rect 157392 5216 157398 5228
rect 157613 5219 157671 5225
rect 157613 5216 157625 5219
rect 157392 5188 157625 5216
rect 157392 5176 157398 5188
rect 157613 5185 157625 5188
rect 157659 5185 157671 5219
rect 157613 5179 157671 5185
rect 158257 5219 158315 5225
rect 158257 5185 158269 5219
rect 158303 5216 158315 5219
rect 158530 5216 158536 5228
rect 158303 5188 158536 5216
rect 158303 5185 158315 5188
rect 158257 5179 158315 5185
rect 158530 5176 158536 5188
rect 158588 5176 158594 5228
rect 155552 5052 156184 5080
rect 155552 5040 155558 5052
rect 151208 4984 152964 5012
rect 153010 4972 153016 5024
rect 153068 5012 153074 5024
rect 153473 5015 153531 5021
rect 153473 5012 153485 5015
rect 153068 4984 153485 5012
rect 153068 4972 153074 4984
rect 153473 4981 153485 4984
rect 153519 4981 153531 5015
rect 153473 4975 153531 4981
rect 154114 4972 154120 5024
rect 154172 5012 154178 5024
rect 154666 5012 154672 5024
rect 154172 4984 154672 5012
rect 154172 4972 154178 4984
rect 154666 4972 154672 4984
rect 154724 5012 154730 5024
rect 155402 5012 155408 5024
rect 154724 4984 155408 5012
rect 154724 4972 154730 4984
rect 155402 4972 155408 4984
rect 155460 4972 155466 5024
rect 156325 5015 156383 5021
rect 156325 4981 156337 5015
rect 156371 5012 156383 5015
rect 157058 5012 157064 5024
rect 156371 4984 157064 5012
rect 156371 4981 156383 4984
rect 156325 4975 156383 4981
rect 157058 4972 157064 4984
rect 157116 4972 157122 5024
rect 157242 4972 157248 5024
rect 157300 5012 157306 5024
rect 157429 5015 157487 5021
rect 157429 5012 157441 5015
rect 157300 4984 157441 5012
rect 157300 4972 157306 4984
rect 157429 4981 157441 4984
rect 157475 4981 157487 5015
rect 157429 4975 157487 4981
rect 1104 4922 158884 4944
rect 1104 4870 20672 4922
rect 20724 4870 20736 4922
rect 20788 4870 20800 4922
rect 20852 4870 20864 4922
rect 20916 4870 20928 4922
rect 20980 4870 60117 4922
rect 60169 4870 60181 4922
rect 60233 4870 60245 4922
rect 60297 4870 60309 4922
rect 60361 4870 60373 4922
rect 60425 4870 99562 4922
rect 99614 4870 99626 4922
rect 99678 4870 99690 4922
rect 99742 4870 99754 4922
rect 99806 4870 99818 4922
rect 99870 4870 139007 4922
rect 139059 4870 139071 4922
rect 139123 4870 139135 4922
rect 139187 4870 139199 4922
rect 139251 4870 139263 4922
rect 139315 4870 158884 4922
rect 1104 4848 158884 4870
rect 4982 4808 4988 4820
rect 4943 4780 4988 4808
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 5994 4808 6000 4820
rect 5767 4780 6000 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 12342 4808 12348 4820
rect 12303 4780 12348 4808
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12676 4780 12817 4808
rect 12676 4768 12682 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 13320 4780 13369 4808
rect 13320 4768 13326 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 13357 4771 13415 4777
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14424 4780 14841 4808
rect 14424 4768 14430 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 14829 4771 14887 4777
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15102 4808 15108 4820
rect 14976 4780 15108 4808
rect 14976 4768 14982 4780
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15933 4811 15991 4817
rect 15933 4777 15945 4811
rect 15979 4808 15991 4811
rect 18230 4808 18236 4820
rect 15979 4780 18236 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 14458 4740 14464 4752
rect 5224 4712 14464 4740
rect 5224 4700 5230 4712
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 15948 4740 15976 4771
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 22741 4811 22799 4817
rect 22741 4808 22753 4811
rect 19760 4780 22753 4808
rect 19760 4768 19766 4780
rect 22741 4777 22753 4780
rect 22787 4777 22799 4811
rect 24670 4808 24676 4820
rect 24631 4780 24676 4808
rect 22741 4771 22799 4777
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 25222 4808 25228 4820
rect 25183 4780 25228 4808
rect 25222 4768 25228 4780
rect 25280 4768 25286 4820
rect 26145 4811 26203 4817
rect 26145 4777 26157 4811
rect 26191 4808 26203 4811
rect 27062 4808 27068 4820
rect 26191 4780 27068 4808
rect 26191 4777 26203 4780
rect 26145 4771 26203 4777
rect 27062 4768 27068 4780
rect 27120 4768 27126 4820
rect 27798 4768 27804 4820
rect 27856 4808 27862 4820
rect 30742 4808 30748 4820
rect 27856 4780 30512 4808
rect 30703 4780 30748 4808
rect 27856 4768 27862 4780
rect 14568 4712 15976 4740
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 14568 4672 14596 4712
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 19484 4712 19840 4740
rect 19484 4700 19490 4712
rect 13688 4644 14596 4672
rect 13688 4632 13694 4644
rect 14826 4632 14832 4684
rect 14884 4672 14890 4684
rect 14884 4644 15240 4672
rect 14884 4632 14890 4644
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5350 4604 5356 4616
rect 5215 4576 5356 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 12158 4604 12164 4616
rect 12119 4576 12164 4604
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13814 4604 13820 4616
rect 13771 4576 13820 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 14936 4536 14964 4644
rect 15212 4613 15240 4644
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 12676 4508 14964 4536
rect 15028 4536 15056 4567
rect 17034 4564 17040 4616
rect 17092 4613 17098 4616
rect 17092 4604 17104 4613
rect 17313 4607 17371 4613
rect 17092 4576 17137 4604
rect 17092 4567 17104 4576
rect 17313 4573 17325 4607
rect 17359 4604 17371 4607
rect 17862 4604 17868 4616
rect 17359 4576 17868 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17092 4564 17098 4567
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 19812 4604 19840 4712
rect 22462 4700 22468 4752
rect 22520 4740 22526 4752
rect 30374 4740 30380 4752
rect 22520 4712 30380 4740
rect 22520 4700 22526 4712
rect 30374 4700 30380 4712
rect 30432 4700 30438 4752
rect 30484 4740 30512 4780
rect 30742 4768 30748 4780
rect 30800 4768 30806 4820
rect 45186 4808 45192 4820
rect 31726 4780 45192 4808
rect 31726 4740 31754 4780
rect 45186 4768 45192 4780
rect 45244 4768 45250 4820
rect 46106 4808 46112 4820
rect 46067 4780 46112 4808
rect 46106 4768 46112 4780
rect 46164 4768 46170 4820
rect 49234 4768 49240 4820
rect 49292 4808 49298 4820
rect 73154 4808 73160 4820
rect 49292 4780 73160 4808
rect 49292 4768 49298 4780
rect 73154 4768 73160 4780
rect 73212 4768 73218 4820
rect 73338 4808 73344 4820
rect 73299 4780 73344 4808
rect 73338 4768 73344 4780
rect 73396 4768 73402 4820
rect 81066 4768 81072 4820
rect 81124 4808 81130 4820
rect 81989 4811 82047 4817
rect 81989 4808 82001 4811
rect 81124 4780 82001 4808
rect 81124 4768 81130 4780
rect 81989 4777 82001 4780
rect 82035 4777 82047 4811
rect 81989 4771 82047 4777
rect 84473 4811 84531 4817
rect 84473 4777 84485 4811
rect 84519 4808 84531 4811
rect 87966 4808 87972 4820
rect 84519 4780 87972 4808
rect 84519 4777 84531 4780
rect 84473 4771 84531 4777
rect 87966 4768 87972 4780
rect 88024 4768 88030 4820
rect 88334 4808 88340 4820
rect 88295 4780 88340 4808
rect 88334 4768 88340 4780
rect 88392 4768 88398 4820
rect 90177 4811 90235 4817
rect 90177 4777 90189 4811
rect 90223 4808 90235 4811
rect 93670 4808 93676 4820
rect 90223 4780 93676 4808
rect 90223 4777 90235 4780
rect 90177 4771 90235 4777
rect 93670 4768 93676 4780
rect 93728 4768 93734 4820
rect 95326 4768 95332 4820
rect 95384 4808 95390 4820
rect 96065 4811 96123 4817
rect 96065 4808 96077 4811
rect 95384 4780 96077 4808
rect 95384 4768 95390 4780
rect 96065 4777 96077 4780
rect 96111 4777 96123 4811
rect 96065 4771 96123 4777
rect 98089 4811 98147 4817
rect 98089 4777 98101 4811
rect 98135 4808 98147 4811
rect 98178 4808 98184 4820
rect 98135 4780 98184 4808
rect 98135 4777 98147 4780
rect 98089 4771 98147 4777
rect 44174 4740 44180 4752
rect 30484 4712 31754 4740
rect 44135 4712 44180 4740
rect 44174 4700 44180 4712
rect 44232 4700 44238 4752
rect 50430 4740 50436 4752
rect 50391 4712 50436 4740
rect 50430 4700 50436 4712
rect 50488 4740 50494 4752
rect 50488 4712 51074 4740
rect 50488 4700 50494 4712
rect 22646 4632 22652 4684
rect 22704 4672 22710 4684
rect 23842 4672 23848 4684
rect 22704 4644 23848 4672
rect 22704 4632 22710 4644
rect 23842 4632 23848 4644
rect 23900 4632 23906 4684
rect 25222 4632 25228 4684
rect 25280 4672 25286 4684
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 25280 4644 25789 4672
rect 25280 4632 25286 4644
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 25777 4635 25835 4641
rect 29917 4675 29975 4681
rect 29917 4641 29929 4675
rect 29963 4672 29975 4675
rect 30558 4672 30564 4684
rect 29963 4644 30564 4672
rect 29963 4641 29975 4644
rect 29917 4635 29975 4641
rect 30558 4632 30564 4644
rect 30616 4672 30622 4684
rect 31018 4672 31024 4684
rect 30616 4644 31024 4672
rect 30616 4632 30622 4644
rect 31018 4632 31024 4644
rect 31076 4632 31082 4684
rect 20634 4607 20692 4613
rect 20634 4604 20646 4607
rect 18012 4576 19748 4604
rect 19812 4576 20646 4604
rect 18012 4564 18018 4576
rect 19720 4536 19748 4576
rect 20634 4573 20646 4576
rect 20680 4573 20692 4607
rect 20634 4567 20692 4573
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21174 4604 21180 4616
rect 20947 4576 21180 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21174 4564 21180 4576
rect 21232 4604 21238 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21232 4576 21373 4604
rect 21232 4564 21238 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 25314 4604 25320 4616
rect 21361 4567 21419 4573
rect 21468 4576 25320 4604
rect 21468 4536 21496 4576
rect 25314 4564 25320 4576
rect 25372 4564 25378 4616
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4604 26019 4607
rect 26605 4607 26663 4613
rect 26605 4604 26617 4607
rect 26007 4576 26617 4604
rect 26007 4573 26019 4576
rect 25961 4567 26019 4573
rect 26605 4573 26617 4576
rect 26651 4573 26663 4607
rect 30098 4604 30104 4616
rect 30059 4576 30104 4604
rect 26605 4567 26663 4573
rect 21634 4545 21640 4548
rect 21628 4536 21640 4545
rect 15028 4508 15240 4536
rect 12676 4496 12682 4508
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14369 4471 14427 4477
rect 14369 4468 14381 4471
rect 13872 4440 14381 4468
rect 13872 4428 13878 4440
rect 14369 4437 14381 4440
rect 14415 4468 14427 4471
rect 15010 4468 15016 4480
rect 14415 4440 15016 4468
rect 14415 4437 14427 4440
rect 14369 4431 14427 4437
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 15212 4468 15240 4508
rect 17236 4508 19656 4536
rect 19720 4508 21496 4536
rect 21595 4508 21640 4536
rect 17236 4468 17264 4508
rect 17862 4468 17868 4480
rect 15212 4440 17264 4468
rect 17823 4440 17868 4468
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 18874 4468 18880 4480
rect 18835 4440 18880 4468
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19518 4468 19524 4480
rect 19479 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19628 4468 19656 4508
rect 21628 4499 21640 4508
rect 21634 4496 21640 4499
rect 21692 4496 21698 4548
rect 25774 4496 25780 4548
rect 25832 4536 25838 4548
rect 25976 4536 26004 4567
rect 30098 4564 30104 4576
rect 30156 4564 30162 4616
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4604 30343 4607
rect 30929 4607 30987 4613
rect 30929 4604 30941 4607
rect 30331 4576 30941 4604
rect 30331 4573 30343 4576
rect 30285 4567 30343 4573
rect 30929 4573 30941 4576
rect 30975 4573 30987 4607
rect 30929 4567 30987 4573
rect 38562 4564 38568 4616
rect 38620 4604 38626 4616
rect 42337 4607 42395 4613
rect 42337 4604 42349 4607
rect 38620 4576 42349 4604
rect 38620 4564 38626 4576
rect 42337 4573 42349 4576
rect 42383 4604 42395 4607
rect 42797 4607 42855 4613
rect 42797 4604 42809 4607
rect 42383 4576 42809 4604
rect 42383 4573 42395 4576
rect 42337 4567 42395 4573
rect 42797 4573 42809 4576
rect 42843 4604 42855 4607
rect 42843 4576 45416 4604
rect 42843 4573 42855 4576
rect 42797 4567 42855 4573
rect 25832 4508 26004 4536
rect 43064 4539 43122 4545
rect 25832 4496 25838 4508
rect 43064 4505 43076 4539
rect 43110 4536 43122 4539
rect 43990 4536 43996 4548
rect 43110 4508 43996 4536
rect 43110 4505 43122 4508
rect 43064 4499 43122 4505
rect 43990 4496 43996 4508
rect 44048 4496 44054 4548
rect 45388 4536 45416 4576
rect 45462 4564 45468 4616
rect 45520 4604 45526 4616
rect 46293 4607 46351 4613
rect 46293 4604 46305 4607
rect 45520 4576 46305 4604
rect 45520 4564 45526 4576
rect 46293 4573 46305 4576
rect 46339 4573 46351 4607
rect 51046 4604 51074 4712
rect 81529 4675 81587 4681
rect 81529 4641 81541 4675
rect 81575 4672 81587 4675
rect 81894 4672 81900 4684
rect 81575 4644 81900 4672
rect 81575 4641 81587 4644
rect 81529 4635 81587 4641
rect 81894 4632 81900 4644
rect 81952 4672 81958 4684
rect 82357 4675 82415 4681
rect 82357 4672 82369 4675
rect 81952 4644 82369 4672
rect 81952 4632 81958 4644
rect 82357 4641 82369 4644
rect 82403 4641 82415 4675
rect 88352 4672 88380 4768
rect 88797 4675 88855 4681
rect 88797 4672 88809 4675
rect 88352 4644 88809 4672
rect 82357 4635 82415 4641
rect 88797 4641 88809 4644
rect 88843 4641 88855 4675
rect 96080 4672 96108 4771
rect 98178 4768 98184 4780
rect 98236 4768 98242 4820
rect 104529 4811 104587 4817
rect 104529 4777 104541 4811
rect 104575 4808 104587 4811
rect 104618 4808 104624 4820
rect 104575 4780 104624 4808
rect 104575 4777 104587 4780
rect 104529 4771 104587 4777
rect 104618 4768 104624 4780
rect 104676 4768 104682 4820
rect 108114 4768 108120 4820
rect 108172 4808 108178 4820
rect 108301 4811 108359 4817
rect 108301 4808 108313 4811
rect 108172 4780 108313 4808
rect 108172 4768 108178 4780
rect 108301 4777 108313 4780
rect 108347 4777 108359 4811
rect 108301 4771 108359 4777
rect 109494 4768 109500 4820
rect 109552 4808 109558 4820
rect 117222 4808 117228 4820
rect 109552 4780 117228 4808
rect 109552 4768 109558 4780
rect 117222 4768 117228 4780
rect 117280 4768 117286 4820
rect 117774 4808 117780 4820
rect 117735 4780 117780 4808
rect 117774 4768 117780 4780
rect 117832 4768 117838 4820
rect 118666 4780 118924 4808
rect 115106 4700 115112 4752
rect 115164 4740 115170 4752
rect 117866 4740 117872 4752
rect 115164 4712 117872 4740
rect 115164 4700 115170 4712
rect 117866 4700 117872 4712
rect 117924 4700 117930 4752
rect 118142 4700 118148 4752
rect 118200 4740 118206 4752
rect 118666 4740 118694 4780
rect 118200 4712 118694 4740
rect 118896 4740 118924 4780
rect 119062 4768 119068 4820
rect 119120 4808 119126 4820
rect 121822 4808 121828 4820
rect 119120 4780 121828 4808
rect 119120 4768 119126 4780
rect 121822 4768 121828 4780
rect 121880 4768 121886 4820
rect 121917 4811 121975 4817
rect 121917 4777 121929 4811
rect 121963 4808 121975 4811
rect 122466 4808 122472 4820
rect 121963 4780 122472 4808
rect 121963 4777 121975 4780
rect 121917 4771 121975 4777
rect 122466 4768 122472 4780
rect 122524 4768 122530 4820
rect 133141 4811 133199 4817
rect 133141 4808 133153 4811
rect 122944 4780 133153 4808
rect 122944 4740 122972 4780
rect 133141 4777 133153 4780
rect 133187 4777 133199 4811
rect 133141 4771 133199 4777
rect 118896 4712 122972 4740
rect 124309 4743 124367 4749
rect 118200 4700 118206 4712
rect 124309 4709 124321 4743
rect 124355 4740 124367 4743
rect 125318 4740 125324 4752
rect 124355 4712 125324 4740
rect 124355 4709 124367 4712
rect 124309 4703 124367 4709
rect 125318 4700 125324 4712
rect 125376 4700 125382 4752
rect 125410 4700 125416 4752
rect 125468 4740 125474 4752
rect 125873 4743 125931 4749
rect 125873 4740 125885 4743
rect 125468 4712 125885 4740
rect 125468 4700 125474 4712
rect 125873 4709 125885 4712
rect 125919 4709 125931 4743
rect 125873 4703 125931 4709
rect 125962 4700 125968 4752
rect 126020 4740 126026 4752
rect 127897 4743 127955 4749
rect 127897 4740 127909 4743
rect 126020 4712 127909 4740
rect 126020 4700 126026 4712
rect 127897 4709 127909 4712
rect 127943 4740 127955 4743
rect 127986 4740 127992 4752
rect 127943 4712 127992 4740
rect 127943 4709 127955 4712
rect 127897 4703 127955 4709
rect 127986 4700 127992 4712
rect 128044 4700 128050 4752
rect 130565 4743 130623 4749
rect 130565 4709 130577 4743
rect 130611 4740 130623 4743
rect 131482 4740 131488 4752
rect 130611 4712 131488 4740
rect 130611 4709 130623 4712
rect 130565 4703 130623 4709
rect 131482 4700 131488 4712
rect 131540 4700 131546 4752
rect 131758 4740 131764 4752
rect 131592 4712 131764 4740
rect 96614 4672 96620 4684
rect 96080 4644 96620 4672
rect 88797 4635 88855 4641
rect 96614 4632 96620 4644
rect 96672 4672 96678 4684
rect 96709 4675 96767 4681
rect 96709 4672 96721 4675
rect 96672 4644 96721 4672
rect 96672 4632 96678 4644
rect 96709 4641 96721 4644
rect 96755 4641 96767 4675
rect 113726 4672 113732 4684
rect 96709 4635 96767 4641
rect 109604 4644 113732 4672
rect 52098 4607 52156 4613
rect 52098 4604 52110 4607
rect 51046 4576 52110 4604
rect 46293 4567 46351 4573
rect 52098 4573 52110 4576
rect 52144 4573 52156 4607
rect 52098 4567 52156 4573
rect 52270 4564 52276 4616
rect 52328 4604 52334 4616
rect 52365 4607 52423 4613
rect 52365 4604 52377 4607
rect 52328 4576 52377 4604
rect 52328 4564 52334 4576
rect 52365 4573 52377 4576
rect 52411 4573 52423 4607
rect 52365 4567 52423 4573
rect 73157 4607 73215 4613
rect 73157 4573 73169 4607
rect 73203 4604 73215 4607
rect 73522 4604 73528 4616
rect 73203 4576 73528 4604
rect 73203 4573 73215 4576
rect 73157 4567 73215 4573
rect 73522 4564 73528 4576
rect 73580 4564 73586 4616
rect 82173 4607 82231 4613
rect 82173 4573 82185 4607
rect 82219 4573 82231 4607
rect 84286 4604 84292 4616
rect 84247 4576 84292 4604
rect 82173 4567 82231 4573
rect 47210 4536 47216 4548
rect 45388 4508 47216 4536
rect 47210 4496 47216 4508
rect 47268 4496 47274 4548
rect 76374 4536 76380 4548
rect 76335 4508 76380 4536
rect 76374 4496 76380 4508
rect 76432 4496 76438 4548
rect 82188 4536 82216 4567
rect 84286 4564 84292 4576
rect 84344 4564 84350 4616
rect 88886 4564 88892 4616
rect 88944 4604 88950 4616
rect 89053 4607 89111 4613
rect 89053 4604 89065 4607
rect 88944 4576 89065 4604
rect 88944 4564 88950 4576
rect 89053 4573 89065 4576
rect 89099 4573 89111 4607
rect 89053 4567 89111 4573
rect 92566 4564 92572 4616
rect 92624 4604 92630 4616
rect 92845 4607 92903 4613
rect 92845 4604 92857 4607
rect 92624 4576 92857 4604
rect 92624 4564 92630 4576
rect 92845 4573 92857 4576
rect 92891 4604 92903 4607
rect 92891 4576 99374 4604
rect 92891 4573 92903 4576
rect 92845 4567 92903 4573
rect 91922 4536 91928 4548
rect 82188 4508 89024 4536
rect 21818 4468 21824 4480
rect 19628 4440 21824 4468
rect 21818 4428 21824 4440
rect 21876 4428 21882 4480
rect 21910 4428 21916 4480
rect 21968 4468 21974 4480
rect 24762 4468 24768 4480
rect 21968 4440 24768 4468
rect 21968 4428 21974 4440
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 50985 4471 51043 4477
rect 50985 4468 50997 4471
rect 26292 4440 50997 4468
rect 26292 4428 26298 4440
rect 50985 4437 50997 4440
rect 51031 4437 51043 4471
rect 88996 4468 89024 4508
rect 89686 4508 91928 4536
rect 89686 4468 89714 4508
rect 91922 4496 91928 4508
rect 91980 4496 91986 4548
rect 96976 4539 97034 4545
rect 96976 4505 96988 4539
rect 97022 4536 97034 4539
rect 98546 4536 98552 4548
rect 97022 4508 98552 4536
rect 97022 4505 97034 4508
rect 96976 4499 97034 4505
rect 98546 4496 98552 4508
rect 98604 4496 98610 4548
rect 99346 4536 99374 4576
rect 101674 4564 101680 4616
rect 101732 4604 101738 4616
rect 105262 4604 105268 4616
rect 101732 4576 105268 4604
rect 101732 4564 101738 4576
rect 105262 4564 105268 4576
rect 105320 4564 105326 4616
rect 108482 4564 108488 4616
rect 108540 4604 108546 4616
rect 109425 4607 109483 4613
rect 109425 4604 109437 4607
rect 108540 4576 109437 4604
rect 108540 4564 108546 4576
rect 109425 4573 109437 4576
rect 109471 4604 109483 4607
rect 109604 4604 109632 4644
rect 113726 4632 113732 4644
rect 113784 4632 113790 4684
rect 114925 4675 114983 4681
rect 114925 4641 114937 4675
rect 114971 4672 114983 4675
rect 116118 4672 116124 4684
rect 114971 4644 116124 4672
rect 114971 4641 114983 4644
rect 114925 4635 114983 4641
rect 116118 4632 116124 4644
rect 116176 4672 116182 4684
rect 116762 4672 116768 4684
rect 116176 4644 116768 4672
rect 116176 4632 116182 4644
rect 116762 4632 116768 4644
rect 116820 4632 116826 4684
rect 118789 4675 118847 4681
rect 118789 4641 118801 4675
rect 118835 4672 118847 4675
rect 119246 4672 119252 4684
rect 118835 4644 119252 4672
rect 118835 4641 118847 4644
rect 118789 4635 118847 4641
rect 119246 4632 119252 4644
rect 119304 4632 119310 4684
rect 122742 4632 122748 4684
rect 122800 4672 122806 4684
rect 122929 4675 122987 4681
rect 122929 4672 122941 4675
rect 122800 4644 122941 4672
rect 122800 4632 122806 4644
rect 122929 4641 122941 4644
rect 122975 4641 122987 4675
rect 122929 4635 122987 4641
rect 109471 4576 109632 4604
rect 109681 4607 109739 4613
rect 109471 4573 109483 4576
rect 109425 4567 109483 4573
rect 109681 4573 109693 4607
rect 109727 4604 109739 4607
rect 109770 4604 109776 4616
rect 109727 4576 109776 4604
rect 109727 4573 109739 4576
rect 109681 4567 109739 4573
rect 109770 4564 109776 4576
rect 109828 4564 109834 4616
rect 114094 4564 114100 4616
rect 114152 4604 114158 4616
rect 118973 4607 119031 4613
rect 114152 4598 118740 4604
rect 114152 4576 118832 4598
rect 114152 4564 114158 4576
rect 118712 4570 118832 4576
rect 109218 4536 109224 4548
rect 99346 4508 109224 4536
rect 109218 4496 109224 4508
rect 109276 4496 109282 4548
rect 114646 4496 114652 4548
rect 114704 4545 114710 4548
rect 114704 4536 114716 4545
rect 114704 4508 114749 4536
rect 114704 4499 114716 4508
rect 114704 4496 114710 4499
rect 115382 4496 115388 4548
rect 115440 4536 115446 4548
rect 117682 4536 117688 4548
rect 115440 4508 117688 4536
rect 115440 4496 115446 4508
rect 117682 4496 117688 4508
rect 117740 4496 117746 4548
rect 118050 4496 118056 4548
rect 118108 4536 118114 4548
rect 118804 4536 118832 4570
rect 118973 4573 118985 4607
rect 119019 4604 119031 4607
rect 119617 4607 119675 4613
rect 119617 4604 119629 4607
rect 119019 4576 119629 4604
rect 119019 4573 119031 4576
rect 118973 4567 119031 4573
rect 119617 4573 119629 4576
rect 119663 4573 119675 4607
rect 122834 4604 122840 4616
rect 119617 4567 119675 4573
rect 120736 4576 122840 4604
rect 118988 4536 119016 4567
rect 120736 4536 120764 4576
rect 122834 4564 122840 4576
rect 122892 4564 122898 4616
rect 122944 4604 122972 4635
rect 124122 4632 124128 4684
rect 124180 4672 124186 4684
rect 126974 4672 126980 4684
rect 124180 4644 126980 4672
rect 124180 4632 124186 4644
rect 126974 4632 126980 4644
rect 127032 4632 127038 4684
rect 129366 4632 129372 4684
rect 129424 4672 129430 4684
rect 131592 4672 131620 4712
rect 131758 4700 131764 4712
rect 131816 4700 131822 4752
rect 133156 4740 133184 4771
rect 134610 4768 134616 4820
rect 134668 4808 134674 4820
rect 135070 4808 135076 4820
rect 134668 4780 135076 4808
rect 134668 4768 134674 4780
rect 135070 4768 135076 4780
rect 135128 4768 135134 4820
rect 135898 4768 135904 4820
rect 135956 4808 135962 4820
rect 135993 4811 136051 4817
rect 135993 4808 136005 4811
rect 135956 4780 136005 4808
rect 135956 4768 135962 4780
rect 135993 4777 136005 4780
rect 136039 4777 136051 4811
rect 135993 4771 136051 4777
rect 138566 4768 138572 4820
rect 138624 4808 138630 4820
rect 140225 4811 140283 4817
rect 140225 4808 140237 4811
rect 138624 4780 140237 4808
rect 138624 4768 138630 4780
rect 140225 4777 140237 4780
rect 140271 4777 140283 4811
rect 140225 4771 140283 4777
rect 143810 4768 143816 4820
rect 143868 4808 143874 4820
rect 146018 4808 146024 4820
rect 143868 4780 146024 4808
rect 143868 4768 143874 4780
rect 146018 4768 146024 4780
rect 146076 4808 146082 4820
rect 146113 4811 146171 4817
rect 146113 4808 146125 4811
rect 146076 4780 146125 4808
rect 146076 4768 146082 4780
rect 146113 4777 146125 4780
rect 146159 4777 146171 4811
rect 151262 4808 151268 4820
rect 146113 4771 146171 4777
rect 146220 4780 151268 4808
rect 133156 4712 133736 4740
rect 129424 4644 131620 4672
rect 131669 4675 131727 4681
rect 129424 4632 129430 4644
rect 131669 4641 131681 4675
rect 131715 4672 131727 4675
rect 132310 4672 132316 4684
rect 131715 4644 132316 4672
rect 131715 4641 131727 4644
rect 131669 4635 131727 4641
rect 132310 4632 132316 4644
rect 132368 4632 132374 4684
rect 133708 4672 133736 4712
rect 138290 4700 138296 4752
rect 138348 4740 138354 4752
rect 139026 4740 139032 4752
rect 138348 4712 139032 4740
rect 138348 4700 138354 4712
rect 139026 4700 139032 4712
rect 139084 4700 139090 4752
rect 139765 4743 139823 4749
rect 139765 4709 139777 4743
rect 139811 4740 139823 4743
rect 140774 4740 140780 4752
rect 139811 4712 140780 4740
rect 139811 4709 139823 4712
rect 139765 4703 139823 4709
rect 140774 4700 140780 4712
rect 140832 4700 140838 4752
rect 145282 4700 145288 4752
rect 145340 4740 145346 4752
rect 145558 4740 145564 4752
rect 145340 4712 145564 4740
rect 145340 4700 145346 4712
rect 145558 4700 145564 4712
rect 145616 4700 145622 4752
rect 145834 4700 145840 4752
rect 145892 4740 145898 4752
rect 146220 4740 146248 4780
rect 151262 4768 151268 4780
rect 151320 4768 151326 4820
rect 151446 4768 151452 4820
rect 151504 4808 151510 4820
rect 152826 4808 152832 4820
rect 151504 4780 152832 4808
rect 151504 4768 151510 4780
rect 152826 4768 152832 4780
rect 152884 4768 152890 4820
rect 152918 4768 152924 4820
rect 152976 4808 152982 4820
rect 156601 4811 156659 4817
rect 156601 4808 156613 4811
rect 152976 4780 156613 4808
rect 152976 4768 152982 4780
rect 156601 4777 156613 4780
rect 156647 4777 156659 4811
rect 156601 4771 156659 4777
rect 157981 4811 158039 4817
rect 157981 4777 157993 4811
rect 158027 4808 158039 4811
rect 159266 4808 159272 4820
rect 158027 4780 159272 4808
rect 158027 4777 158039 4780
rect 157981 4771 158039 4777
rect 159266 4768 159272 4780
rect 159324 4768 159330 4820
rect 150066 4740 150072 4752
rect 145892 4712 146248 4740
rect 150027 4712 150072 4740
rect 145892 4700 145898 4712
rect 150066 4700 150072 4712
rect 150124 4700 150130 4752
rect 152182 4700 152188 4752
rect 152240 4740 152246 4752
rect 152458 4740 152464 4752
rect 152240 4712 152464 4740
rect 152240 4700 152246 4712
rect 152458 4700 152464 4712
rect 152516 4700 152522 4752
rect 154298 4700 154304 4752
rect 154356 4740 154362 4752
rect 154393 4743 154451 4749
rect 154393 4740 154405 4743
rect 154356 4712 154405 4740
rect 154356 4700 154362 4712
rect 154393 4709 154405 4712
rect 154439 4709 154451 4743
rect 157242 4740 157248 4752
rect 154393 4703 154451 4709
rect 155420 4712 157248 4740
rect 137925 4675 137983 4681
rect 137925 4672 137937 4675
rect 133708 4644 133828 4672
rect 123938 4604 123944 4616
rect 122944 4576 123944 4604
rect 123938 4564 123944 4576
rect 123996 4604 124002 4616
rect 125321 4607 125379 4613
rect 125321 4604 125333 4607
rect 123996 4576 125333 4604
rect 123996 4564 124002 4576
rect 125321 4573 125333 4576
rect 125367 4604 125379 4607
rect 129277 4607 129335 4613
rect 129277 4604 129289 4607
rect 125367 4576 129289 4604
rect 125367 4573 125379 4576
rect 125321 4567 125379 4573
rect 129277 4573 129289 4576
rect 129323 4604 129335 4607
rect 129737 4607 129795 4613
rect 129737 4604 129749 4607
rect 129323 4576 129749 4604
rect 129323 4573 129335 4576
rect 129277 4567 129335 4573
rect 129737 4573 129749 4576
rect 129783 4604 129795 4607
rect 133046 4604 133052 4616
rect 129783 4576 133052 4604
rect 129783 4573 129795 4576
rect 129737 4567 129795 4573
rect 133046 4564 133052 4576
rect 133104 4564 133110 4616
rect 133598 4564 133604 4616
rect 133656 4604 133662 4616
rect 133693 4607 133751 4613
rect 133693 4604 133705 4607
rect 133656 4576 133705 4604
rect 133656 4564 133662 4576
rect 133693 4573 133705 4576
rect 133739 4573 133751 4607
rect 133800 4604 133828 4644
rect 137388 4644 137937 4672
rect 133949 4607 134007 4613
rect 133949 4604 133961 4607
rect 133800 4576 133961 4604
rect 133693 4567 133751 4573
rect 133949 4573 133961 4576
rect 133995 4573 134007 4607
rect 133949 4567 134007 4573
rect 135714 4564 135720 4616
rect 135772 4604 135778 4616
rect 137388 4613 137416 4644
rect 137925 4641 137937 4644
rect 137971 4641 137983 4675
rect 137925 4635 137983 4641
rect 138569 4675 138627 4681
rect 138569 4641 138581 4675
rect 138615 4672 138627 4675
rect 142430 4672 142436 4684
rect 138615 4644 140728 4672
rect 142391 4644 142436 4672
rect 138615 4641 138627 4644
rect 138569 4635 138627 4641
rect 137373 4607 137431 4613
rect 137373 4604 137385 4607
rect 135772 4576 137385 4604
rect 135772 4564 135778 4576
rect 137373 4573 137385 4576
rect 137419 4573 137431 4607
rect 138382 4604 138388 4616
rect 137373 4567 137431 4573
rect 137572 4576 138388 4604
rect 118108 4508 118694 4536
rect 118804 4508 119016 4536
rect 119080 4508 120764 4536
rect 120813 4539 120871 4545
rect 118108 4496 118114 4508
rect 88996 4440 89714 4468
rect 50985 4431 51043 4437
rect 101766 4428 101772 4480
rect 101824 4468 101830 4480
rect 112162 4468 112168 4480
rect 101824 4440 112168 4468
rect 101824 4428 101830 4440
rect 112162 4428 112168 4440
rect 112220 4428 112226 4480
rect 113542 4468 113548 4480
rect 113503 4440 113548 4468
rect 113542 4428 113548 4440
rect 113600 4428 113606 4480
rect 115477 4471 115535 4477
rect 115477 4437 115489 4471
rect 115523 4468 115535 4471
rect 115566 4468 115572 4480
rect 115523 4440 115572 4468
rect 115523 4437 115535 4440
rect 115477 4431 115535 4437
rect 115566 4428 115572 4440
rect 115624 4428 115630 4480
rect 115842 4428 115848 4480
rect 115900 4468 115906 4480
rect 118142 4468 118148 4480
rect 115900 4440 118148 4468
rect 115900 4428 115906 4440
rect 118142 4428 118148 4440
rect 118200 4428 118206 4480
rect 118666 4468 118694 4508
rect 119080 4468 119108 4508
rect 120813 4505 120825 4539
rect 120859 4536 120871 4539
rect 123196 4539 123254 4545
rect 120859 4508 123156 4536
rect 120859 4505 120871 4508
rect 120813 4499 120871 4505
rect 118666 4440 119108 4468
rect 119157 4471 119215 4477
rect 119157 4437 119169 4471
rect 119203 4468 119215 4471
rect 119246 4468 119252 4480
rect 119203 4440 119252 4468
rect 119203 4437 119215 4440
rect 119157 4431 119215 4437
rect 119246 4428 119252 4440
rect 119304 4428 119310 4480
rect 120261 4471 120319 4477
rect 120261 4437 120273 4471
rect 120307 4468 120319 4471
rect 120350 4468 120356 4480
rect 120307 4440 120356 4468
rect 120307 4437 120319 4440
rect 120261 4431 120319 4437
rect 120350 4428 120356 4440
rect 120408 4428 120414 4480
rect 121178 4428 121184 4480
rect 121236 4468 121242 4480
rect 121273 4471 121331 4477
rect 121273 4468 121285 4471
rect 121236 4440 121285 4468
rect 121236 4428 121242 4440
rect 121273 4437 121285 4440
rect 121319 4437 121331 4471
rect 123128 4468 123156 4508
rect 123196 4505 123208 4539
rect 123242 4536 123254 4539
rect 123242 4508 124904 4536
rect 123242 4505 123254 4508
rect 123196 4499 123254 4505
rect 124876 4480 124904 4508
rect 125410 4496 125416 4548
rect 125468 4536 125474 4548
rect 126425 4539 126483 4545
rect 126425 4536 126437 4539
rect 125468 4508 126437 4536
rect 125468 4496 125474 4508
rect 126425 4505 126437 4508
rect 126471 4536 126483 4539
rect 128906 4536 128912 4548
rect 126471 4508 128912 4536
rect 126471 4505 126483 4508
rect 126425 4499 126483 4505
rect 128906 4496 128912 4508
rect 128964 4496 128970 4548
rect 129032 4539 129090 4545
rect 129032 4505 129044 4539
rect 129078 4536 129090 4539
rect 129826 4536 129832 4548
rect 129078 4508 129832 4536
rect 129078 4505 129090 4508
rect 129032 4499 129090 4505
rect 129826 4496 129832 4508
rect 129884 4496 129890 4548
rect 137128 4539 137186 4545
rect 130396 4508 133276 4536
rect 124122 4468 124128 4480
rect 123128 4440 124128 4468
rect 121273 4431 121331 4437
rect 124122 4428 124128 4440
rect 124180 4428 124186 4480
rect 124858 4468 124864 4480
rect 124819 4440 124864 4468
rect 124858 4428 124864 4440
rect 124916 4428 124922 4480
rect 126514 4428 126520 4480
rect 126572 4468 126578 4480
rect 127802 4468 127808 4480
rect 126572 4440 127808 4468
rect 126572 4428 126578 4440
rect 127802 4428 127808 4440
rect 127860 4428 127866 4480
rect 127986 4428 127992 4480
rect 128044 4468 128050 4480
rect 130396 4468 130424 4508
rect 131114 4468 131120 4480
rect 128044 4440 130424 4468
rect 131075 4440 131120 4468
rect 128044 4428 128050 4440
rect 131114 4428 131120 4440
rect 131172 4428 131178 4480
rect 132221 4471 132279 4477
rect 132221 4437 132233 4471
rect 132267 4468 132279 4471
rect 132494 4468 132500 4480
rect 132267 4440 132500 4468
rect 132267 4437 132279 4440
rect 132221 4431 132279 4437
rect 132494 4428 132500 4440
rect 132552 4428 132558 4480
rect 133248 4468 133276 4508
rect 134076 4508 135254 4536
rect 134076 4468 134104 4508
rect 133248 4440 134104 4468
rect 135226 4468 135254 4508
rect 137128 4505 137140 4539
rect 137174 4536 137186 4539
rect 137572 4536 137600 4576
rect 138382 4564 138388 4576
rect 138440 4564 138446 4616
rect 137174 4508 137600 4536
rect 137174 4505 137186 4508
rect 137128 4499 137186 4505
rect 138584 4468 138612 4635
rect 139581 4607 139639 4613
rect 139581 4573 139593 4607
rect 139627 4604 139639 4607
rect 139946 4604 139952 4616
rect 139627 4576 139952 4604
rect 139627 4573 139639 4576
rect 139581 4567 139639 4573
rect 139946 4564 139952 4576
rect 140004 4564 140010 4616
rect 140409 4607 140467 4613
rect 140409 4573 140421 4607
rect 140455 4573 140467 4607
rect 140590 4604 140596 4616
rect 140551 4576 140596 4604
rect 140409 4567 140467 4573
rect 139026 4496 139032 4548
rect 139084 4536 139090 4548
rect 140424 4536 140452 4567
rect 140590 4564 140596 4576
rect 140648 4564 140654 4616
rect 140700 4604 140728 4644
rect 142430 4632 142436 4644
rect 142488 4632 142494 4684
rect 147490 4672 147496 4684
rect 142540 4644 143212 4672
rect 147451 4644 147496 4672
rect 142540 4604 142568 4644
rect 143074 4604 143080 4616
rect 140700 4576 142568 4604
rect 143035 4576 143080 4604
rect 143074 4564 143080 4576
rect 143132 4564 143138 4616
rect 143184 4604 143212 4644
rect 147490 4632 147496 4644
rect 147548 4672 147554 4684
rect 148229 4675 148287 4681
rect 148229 4672 148241 4675
rect 147548 4644 148241 4672
rect 147548 4632 147554 4644
rect 148229 4641 148241 4644
rect 148275 4641 148287 4675
rect 155420 4672 155448 4712
rect 157242 4700 157248 4712
rect 157300 4700 157306 4752
rect 148229 4635 148287 4641
rect 151372 4644 155448 4672
rect 155497 4675 155555 4681
rect 143261 4607 143319 4613
rect 143261 4604 143273 4607
rect 143184 4576 143273 4604
rect 143261 4573 143273 4576
rect 143307 4573 143319 4607
rect 143261 4567 143319 4573
rect 143350 4564 143356 4616
rect 143408 4604 143414 4616
rect 144178 4604 144184 4616
rect 143408 4576 144184 4604
rect 143408 4564 143414 4576
rect 144178 4564 144184 4576
rect 144236 4564 144242 4616
rect 144270 4564 144276 4616
rect 144328 4604 144334 4616
rect 144540 4607 144598 4613
rect 144328 4576 144373 4604
rect 144328 4564 144334 4576
rect 144540 4573 144552 4607
rect 144586 4604 144598 4607
rect 145834 4604 145840 4616
rect 144586 4576 145840 4604
rect 144586 4573 144598 4576
rect 144540 4567 144598 4573
rect 145834 4564 145840 4576
rect 145892 4564 145898 4616
rect 147674 4604 147680 4616
rect 147140 4576 147680 4604
rect 139084 4508 140452 4536
rect 142188 4539 142246 4545
rect 139084 4496 139090 4508
rect 142188 4505 142200 4539
rect 142234 4536 142246 4539
rect 147140 4536 147168 4576
rect 147674 4564 147680 4576
rect 147732 4564 147738 4616
rect 148496 4607 148554 4613
rect 148496 4573 148508 4607
rect 148542 4604 148554 4607
rect 151372 4604 151400 4644
rect 155497 4641 155509 4675
rect 155543 4672 155555 4675
rect 159358 4672 159364 4684
rect 155543 4644 159364 4672
rect 155543 4641 155555 4644
rect 155497 4635 155555 4641
rect 159358 4632 159364 4644
rect 159416 4632 159422 4684
rect 148542 4576 151400 4604
rect 151449 4607 151507 4613
rect 148542 4573 148554 4576
rect 148496 4567 148554 4573
rect 151449 4573 151461 4607
rect 151495 4604 151507 4607
rect 151814 4604 151820 4616
rect 151495 4576 151820 4604
rect 151495 4573 151507 4576
rect 151449 4567 151507 4573
rect 151814 4564 151820 4576
rect 151872 4564 151878 4616
rect 151909 4607 151967 4613
rect 151909 4573 151921 4607
rect 151955 4573 151967 4607
rect 152090 4604 152096 4616
rect 152051 4576 152096 4604
rect 151909 4567 151967 4573
rect 142234 4508 147168 4536
rect 147248 4539 147306 4545
rect 142234 4505 142246 4508
rect 142188 4499 142246 4505
rect 147248 4505 147260 4539
rect 147294 4536 147306 4539
rect 151078 4536 151084 4548
rect 147294 4508 151084 4536
rect 147294 4505 147306 4508
rect 147248 4499 147306 4505
rect 151078 4496 151084 4508
rect 151136 4496 151142 4548
rect 151182 4539 151240 4545
rect 151182 4505 151194 4539
rect 151228 4505 151240 4539
rect 151182 4499 151240 4505
rect 141050 4468 141056 4480
rect 135226 4440 138612 4468
rect 141011 4440 141056 4468
rect 141050 4428 141056 4440
rect 141108 4428 141114 4480
rect 141418 4428 141424 4480
rect 141476 4468 141482 4480
rect 145558 4468 145564 4480
rect 141476 4440 145564 4468
rect 141476 4428 141482 4440
rect 145558 4428 145564 4440
rect 145616 4428 145622 4480
rect 145653 4471 145711 4477
rect 145653 4437 145665 4471
rect 145699 4468 145711 4471
rect 146754 4468 146760 4480
rect 145699 4440 146760 4468
rect 145699 4437 145711 4440
rect 145653 4431 145711 4437
rect 146754 4428 146760 4440
rect 146812 4428 146818 4480
rect 146938 4428 146944 4480
rect 146996 4468 147002 4480
rect 149422 4468 149428 4480
rect 146996 4440 149428 4468
rect 146996 4428 147002 4440
rect 149422 4428 149428 4440
rect 149480 4468 149486 4480
rect 149609 4471 149667 4477
rect 149609 4468 149621 4471
rect 149480 4440 149621 4468
rect 149480 4428 149486 4440
rect 149609 4437 149621 4440
rect 149655 4437 149667 4471
rect 149609 4431 149667 4437
rect 149882 4428 149888 4480
rect 149940 4468 149946 4480
rect 151188 4468 151216 4499
rect 151630 4496 151636 4548
rect 151688 4536 151694 4548
rect 151924 4536 151952 4567
rect 152090 4564 152096 4576
rect 152148 4564 152154 4616
rect 153562 4604 153568 4616
rect 153523 4576 153568 4604
rect 153562 4564 153568 4576
rect 153620 4564 153626 4616
rect 153654 4564 153660 4616
rect 153712 4604 153718 4616
rect 153749 4607 153807 4613
rect 153749 4604 153761 4607
rect 153712 4576 153761 4604
rect 153712 4564 153718 4576
rect 153749 4573 153761 4576
rect 153795 4573 153807 4607
rect 154574 4604 154580 4616
rect 154535 4576 154580 4604
rect 153749 4567 153807 4573
rect 154574 4564 154580 4576
rect 154632 4564 154638 4616
rect 155126 4604 155132 4616
rect 155087 4576 155132 4604
rect 155126 4564 155132 4576
rect 155184 4564 155190 4616
rect 155218 4564 155224 4616
rect 155276 4604 155282 4616
rect 155313 4607 155371 4613
rect 155313 4604 155325 4607
rect 155276 4576 155325 4604
rect 155276 4564 155282 4576
rect 155313 4573 155325 4576
rect 155359 4573 155371 4607
rect 156138 4604 156144 4616
rect 156099 4576 156144 4604
rect 155313 4567 155371 4573
rect 156138 4564 156144 4576
rect 156196 4564 156202 4616
rect 156785 4607 156843 4613
rect 156785 4573 156797 4607
rect 156831 4604 156843 4607
rect 156874 4604 156880 4616
rect 156831 4576 156880 4604
rect 156831 4573 156843 4576
rect 156785 4567 156843 4573
rect 156874 4564 156880 4576
rect 156932 4564 156938 4616
rect 157429 4607 157487 4613
rect 157429 4573 157441 4607
rect 157475 4604 157487 4607
rect 157978 4604 157984 4616
rect 157475 4576 157984 4604
rect 157475 4573 157487 4576
rect 157429 4567 157487 4573
rect 157978 4564 157984 4576
rect 158036 4564 158042 4616
rect 151688 4508 151952 4536
rect 153933 4539 153991 4545
rect 151688 4496 151694 4508
rect 153933 4505 153945 4539
rect 153979 4536 153991 4539
rect 154942 4536 154948 4548
rect 153979 4508 154948 4536
rect 153979 4505 153991 4508
rect 153933 4499 153991 4505
rect 154942 4496 154948 4508
rect 155000 4496 155006 4548
rect 152274 4468 152280 4480
rect 149940 4440 151216 4468
rect 152235 4440 152280 4468
rect 149940 4428 149946 4440
rect 152274 4428 152280 4440
rect 152332 4428 152338 4480
rect 155310 4428 155316 4480
rect 155368 4468 155374 4480
rect 155957 4471 156015 4477
rect 155957 4468 155969 4471
rect 155368 4440 155969 4468
rect 155368 4428 155374 4440
rect 155957 4437 155969 4440
rect 156003 4437 156015 4471
rect 157242 4468 157248 4480
rect 157203 4440 157248 4468
rect 155957 4431 156015 4437
rect 157242 4428 157248 4440
rect 157300 4428 157306 4480
rect 1104 4378 159043 4400
rect 1104 4326 40394 4378
rect 40446 4326 40458 4378
rect 40510 4326 40522 4378
rect 40574 4326 40586 4378
rect 40638 4326 40650 4378
rect 40702 4326 79839 4378
rect 79891 4326 79903 4378
rect 79955 4326 79967 4378
rect 80019 4326 80031 4378
rect 80083 4326 80095 4378
rect 80147 4326 119284 4378
rect 119336 4326 119348 4378
rect 119400 4326 119412 4378
rect 119464 4326 119476 4378
rect 119528 4326 119540 4378
rect 119592 4326 158729 4378
rect 158781 4326 158793 4378
rect 158845 4326 158857 4378
rect 158909 4326 158921 4378
rect 158973 4326 158985 4378
rect 159037 4326 159043 4378
rect 1104 4304 159043 4326
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 19518 4264 19524 4276
rect 10468 4236 19524 4264
rect 10468 4224 10474 4236
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 42613 4267 42671 4273
rect 42613 4264 42625 4267
rect 20220 4236 42625 4264
rect 20220 4224 20226 4236
rect 42613 4233 42625 4236
rect 42659 4233 42671 4267
rect 42613 4227 42671 4233
rect 43070 4224 43076 4276
rect 43128 4264 43134 4276
rect 56778 4264 56784 4276
rect 43128 4236 56784 4264
rect 43128 4224 43134 4236
rect 56778 4224 56784 4236
rect 56836 4224 56842 4276
rect 62301 4267 62359 4273
rect 62301 4233 62313 4267
rect 62347 4264 62359 4267
rect 63310 4264 63316 4276
rect 62347 4236 63316 4264
rect 62347 4233 62359 4236
rect 62301 4227 62359 4233
rect 12618 4196 12624 4208
rect 12579 4168 12624 4196
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 14274 4196 14280 4208
rect 13832 4168 14280 4196
rect 13832 4140 13860 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 16816 4168 16865 4196
rect 16816 4156 16822 4168
rect 16853 4165 16865 4168
rect 16899 4165 16911 4199
rect 16853 4159 16911 4165
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 21174 4196 21180 4208
rect 18932 4168 21180 4196
rect 18932 4156 18938 4168
rect 21174 4156 21180 4168
rect 21232 4156 21238 4208
rect 23658 4156 23664 4208
rect 23716 4196 23722 4208
rect 30377 4199 30435 4205
rect 23716 4168 24880 4196
rect 23716 4156 23722 4168
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 9122 4128 9128 4140
rect 8343 4100 9128 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10962 4128 10968 4140
rect 9640 4100 10968 4128
rect 9640 4088 9646 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 13814 4128 13820 4140
rect 13727 4100 13820 4128
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14073 4131 14131 4137
rect 14073 4128 14085 4131
rect 13964 4100 14085 4128
rect 13964 4088 13970 4100
rect 14073 4097 14085 4100
rect 14119 4097 14131 4131
rect 15654 4128 15660 4140
rect 15615 4100 15660 4128
rect 14073 4091 14131 4097
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16776 4128 16804 4156
rect 17678 4128 17684 4140
rect 16071 4100 16804 4128
rect 17639 4100 17684 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4060 12403 4063
rect 13722 4060 13728 4072
rect 12391 4032 13728 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 8113 3995 8171 4001
rect 8113 3992 8125 3995
rect 6880 3964 8125 3992
rect 6880 3952 6886 3964
rect 8113 3961 8125 3964
rect 8159 3961 8171 3995
rect 15856 3992 15884 4091
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18506 4128 18512 4140
rect 17920 4100 18512 4128
rect 17920 4088 17926 4100
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18782 4137 18788 4140
rect 18776 4091 18788 4137
rect 18840 4128 18846 4140
rect 18840 4100 18876 4128
rect 18782 4088 18788 4091
rect 18840 4088 18846 4100
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20349 4131 20407 4137
rect 20349 4128 20361 4131
rect 20128 4100 20361 4128
rect 20128 4088 20134 4100
rect 20349 4097 20361 4100
rect 20395 4097 20407 4131
rect 20349 4091 20407 4097
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 24578 4128 24584 4140
rect 20496 4100 24584 4128
rect 20496 4088 20502 4100
rect 24578 4088 24584 4100
rect 24636 4088 24642 4140
rect 24852 4128 24880 4168
rect 30377 4165 30389 4199
rect 30423 4196 30435 4199
rect 30558 4196 30564 4208
rect 30423 4168 30564 4196
rect 30423 4165 30435 4168
rect 30377 4159 30435 4165
rect 30558 4156 30564 4168
rect 30616 4156 30622 4208
rect 50982 4196 50988 4208
rect 42996 4168 43576 4196
rect 42886 4128 42892 4140
rect 24852 4100 42892 4128
rect 42886 4088 42892 4100
rect 42944 4088 42950 4140
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 30558 4060 30564 4072
rect 19576 4032 30564 4060
rect 19576 4020 19582 4032
rect 30558 4020 30564 4032
rect 30616 4020 30622 4072
rect 31846 4020 31852 4072
rect 31904 4060 31910 4072
rect 37182 4060 37188 4072
rect 31904 4032 37188 4060
rect 31904 4020 31910 4032
rect 37182 4020 37188 4032
rect 37240 4020 37246 4072
rect 41966 4060 41972 4072
rect 41927 4032 41972 4060
rect 41966 4020 41972 4032
rect 42024 4060 42030 4072
rect 42996 4060 43024 4168
rect 43548 4128 43576 4168
rect 47780 4168 48075 4196
rect 43726 4131 43784 4137
rect 43726 4128 43738 4131
rect 43548 4100 43738 4128
rect 43726 4097 43738 4100
rect 43772 4097 43784 4131
rect 43726 4091 43784 4097
rect 43993 4131 44051 4137
rect 43993 4097 44005 4131
rect 44039 4128 44051 4131
rect 44174 4128 44180 4140
rect 44039 4100 44180 4128
rect 44039 4097 44051 4100
rect 43993 4091 44051 4097
rect 44174 4088 44180 4100
rect 44232 4128 44238 4140
rect 44634 4128 44640 4140
rect 44232 4100 44640 4128
rect 44232 4088 44238 4100
rect 44634 4088 44640 4100
rect 44692 4088 44698 4140
rect 45278 4088 45284 4140
rect 45336 4128 45342 4140
rect 47780 4128 47808 4168
rect 47946 4128 47952 4140
rect 45336 4100 47808 4128
rect 47907 4100 47952 4128
rect 45336 4088 45342 4100
rect 47946 4088 47952 4100
rect 48004 4088 48010 4140
rect 48047 4128 48075 4168
rect 50908 4168 50988 4196
rect 50908 4137 50936 4168
rect 50982 4156 50988 4168
rect 51040 4156 51046 4208
rect 50893 4131 50951 4137
rect 48047 4100 50844 4128
rect 49786 4060 49792 4072
rect 42024 4032 43024 4060
rect 45388 4032 49792 4060
rect 42024 4020 42030 4032
rect 30466 3992 30472 4004
rect 15856 3964 18552 3992
rect 8113 3955 8171 3961
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3924 11762 3936
rect 12618 3924 12624 3936
rect 11756 3896 12624 3924
rect 11756 3884 11762 3896
rect 12618 3884 12624 3896
rect 12676 3924 12682 3936
rect 13262 3924 13268 3936
rect 12676 3896 13268 3924
rect 12676 3884 12682 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13357 3927 13415 3933
rect 13357 3893 13369 3927
rect 13403 3924 13415 3927
rect 13538 3924 13544 3936
rect 13403 3896 13544 3924
rect 13403 3893 13415 3896
rect 13357 3887 13415 3893
rect 13538 3884 13544 3896
rect 13596 3924 13602 3936
rect 15194 3924 15200 3936
rect 13596 3896 15200 3924
rect 13596 3884 13602 3896
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 17865 3927 17923 3933
rect 17865 3893 17877 3927
rect 17911 3924 17923 3927
rect 18414 3924 18420 3936
rect 17911 3896 18420 3924
rect 17911 3893 17923 3896
rect 17865 3887 17923 3893
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18524 3924 18552 3964
rect 19904 3964 30472 3992
rect 19904 3933 19932 3964
rect 30466 3952 30472 3964
rect 30524 3952 30530 4004
rect 30834 3952 30840 4004
rect 30892 3992 30898 4004
rect 30892 3964 32904 3992
rect 30892 3952 30898 3964
rect 32876 3936 32904 3964
rect 34422 3952 34428 4004
rect 34480 3992 34486 4004
rect 34480 3964 43116 3992
rect 34480 3952 34486 3964
rect 19889 3927 19947 3933
rect 19889 3924 19901 3927
rect 18524 3896 19901 3924
rect 19889 3893 19901 3896
rect 19935 3893 19947 3927
rect 21174 3924 21180 3936
rect 21135 3896 21180 3924
rect 19889 3887 19947 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 31110 3884 31116 3936
rect 31168 3924 31174 3936
rect 31754 3924 31760 3936
rect 31168 3896 31760 3924
rect 31168 3884 31174 3896
rect 31754 3884 31760 3896
rect 31812 3884 31818 3936
rect 32858 3924 32864 3936
rect 32819 3896 32864 3924
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 43088 3924 43116 3964
rect 45388 3924 45416 4032
rect 49786 4020 49792 4032
rect 49844 4020 49850 4072
rect 50816 4060 50844 4100
rect 50893 4097 50905 4131
rect 50939 4097 50951 4131
rect 55410 4131 55468 4137
rect 55410 4128 55422 4131
rect 50893 4091 50951 4097
rect 51046 4100 55422 4128
rect 51046 4060 51074 4100
rect 55410 4097 55422 4100
rect 55456 4097 55468 4131
rect 55410 4091 55468 4097
rect 61493 4131 61551 4137
rect 61493 4097 61505 4131
rect 61539 4128 61551 4131
rect 61749 4131 61807 4137
rect 61539 4100 61700 4128
rect 61539 4097 61551 4100
rect 61493 4091 61551 4097
rect 50816 4032 51074 4060
rect 55677 4063 55735 4069
rect 55677 4029 55689 4063
rect 55723 4060 55735 4063
rect 56137 4063 56195 4069
rect 56137 4060 56149 4063
rect 55723 4032 56149 4060
rect 55723 4029 55735 4032
rect 55677 4023 55735 4029
rect 56137 4029 56149 4032
rect 56183 4060 56195 4063
rect 58526 4060 58532 4072
rect 56183 4032 58532 4060
rect 56183 4029 56195 4032
rect 56137 4023 56195 4029
rect 45462 3952 45468 4004
rect 45520 3992 45526 4004
rect 54297 3995 54355 4001
rect 54297 3992 54309 3995
rect 45520 3964 54309 3992
rect 45520 3952 45526 3964
rect 54297 3961 54309 3964
rect 54343 3961 54355 3995
rect 54297 3955 54355 3961
rect 43088 3896 45416 3924
rect 47578 3884 47584 3936
rect 47636 3924 47642 3936
rect 47765 3927 47823 3933
rect 47765 3924 47777 3927
rect 47636 3896 47777 3924
rect 47636 3884 47642 3896
rect 47765 3893 47777 3896
rect 47811 3893 47823 3927
rect 47765 3887 47823 3893
rect 48958 3884 48964 3936
rect 49016 3924 49022 3936
rect 50709 3927 50767 3933
rect 50709 3924 50721 3927
rect 49016 3896 50721 3924
rect 49016 3884 49022 3896
rect 50709 3893 50721 3896
rect 50755 3893 50767 3927
rect 50709 3887 50767 3893
rect 54662 3884 54668 3936
rect 54720 3924 54726 3936
rect 55692 3924 55720 4023
rect 58526 4020 58532 4032
rect 58584 4020 58590 4072
rect 61672 4060 61700 4100
rect 61749 4097 61761 4131
rect 61795 4128 61807 4131
rect 62114 4128 62120 4140
rect 61795 4100 62120 4128
rect 61795 4097 61807 4100
rect 61749 4091 61807 4097
rect 62114 4088 62120 4100
rect 62172 4128 62178 4140
rect 62316 4128 62344 4227
rect 63310 4224 63316 4236
rect 63368 4224 63374 4276
rect 98546 4224 98552 4276
rect 98604 4264 98610 4276
rect 110322 4264 110328 4276
rect 98604 4236 110328 4264
rect 98604 4224 98610 4236
rect 110322 4224 110328 4236
rect 110380 4224 110386 4276
rect 113726 4224 113732 4276
rect 113784 4264 113790 4276
rect 118786 4264 118792 4276
rect 113784 4236 118792 4264
rect 113784 4224 113790 4236
rect 118786 4224 118792 4236
rect 118844 4224 118850 4276
rect 125042 4264 125048 4276
rect 125003 4236 125048 4264
rect 125042 4224 125048 4236
rect 125100 4224 125106 4276
rect 127526 4224 127532 4276
rect 127584 4264 127590 4276
rect 127584 4236 133092 4264
rect 127584 4224 127590 4236
rect 105170 4196 105176 4208
rect 104820 4168 105176 4196
rect 62172 4100 62344 4128
rect 75917 4131 75975 4137
rect 62172 4088 62178 4100
rect 75917 4097 75929 4131
rect 75963 4128 75975 4131
rect 76374 4128 76380 4140
rect 75963 4100 76380 4128
rect 75963 4097 75975 4100
rect 75917 4091 75975 4097
rect 76374 4088 76380 4100
rect 76432 4088 76438 4140
rect 78950 4088 78956 4140
rect 79008 4128 79014 4140
rect 79413 4131 79471 4137
rect 79413 4128 79425 4131
rect 79008 4100 79425 4128
rect 79008 4088 79014 4100
rect 79413 4097 79425 4100
rect 79459 4097 79471 4131
rect 79413 4091 79471 4097
rect 104621 4131 104679 4137
rect 104621 4097 104633 4131
rect 104667 4128 104679 4131
rect 104820 4128 104848 4168
rect 105170 4156 105176 4168
rect 105228 4156 105234 4208
rect 105262 4156 105268 4208
rect 105320 4196 105326 4208
rect 105320 4168 111647 4196
rect 105320 4156 105326 4168
rect 104667 4100 104848 4128
rect 104888 4131 104946 4137
rect 104667 4097 104679 4100
rect 104621 4091 104679 4097
rect 104888 4097 104900 4131
rect 104934 4128 104946 4131
rect 106461 4131 106519 4137
rect 106461 4128 106473 4131
rect 104934 4100 106473 4128
rect 104934 4097 104946 4100
rect 104888 4091 104946 4097
rect 106461 4097 106473 4100
rect 106507 4128 106519 4131
rect 106550 4128 106556 4140
rect 106507 4100 106556 4128
rect 106507 4097 106519 4100
rect 106461 4091 106519 4097
rect 106550 4088 106556 4100
rect 106608 4088 106614 4140
rect 108781 4131 108839 4137
rect 108781 4097 108793 4131
rect 108827 4128 108839 4131
rect 109310 4128 109316 4140
rect 108827 4100 109316 4128
rect 108827 4097 108839 4100
rect 108781 4091 108839 4097
rect 109310 4088 109316 4100
rect 109368 4088 109374 4140
rect 110713 4131 110771 4137
rect 110713 4097 110725 4131
rect 110759 4128 110771 4131
rect 111150 4128 111156 4140
rect 110759 4100 111156 4128
rect 110759 4097 110771 4100
rect 110713 4091 110771 4097
rect 111150 4088 111156 4100
rect 111208 4088 111214 4140
rect 64874 4060 64880 4072
rect 61672 4032 64880 4060
rect 64874 4020 64880 4032
rect 64932 4020 64938 4072
rect 76006 4020 76012 4072
rect 76064 4060 76070 4072
rect 76193 4063 76251 4069
rect 76193 4060 76205 4063
rect 76064 4032 76205 4060
rect 76064 4020 76070 4032
rect 76193 4029 76205 4032
rect 76239 4060 76251 4063
rect 76653 4063 76711 4069
rect 76653 4060 76665 4063
rect 76239 4032 76665 4060
rect 76239 4029 76251 4032
rect 76193 4023 76251 4029
rect 76653 4029 76665 4032
rect 76699 4029 76711 4063
rect 109034 4060 109040 4072
rect 108995 4032 109040 4060
rect 76653 4023 76711 4029
rect 109034 4020 109040 4032
rect 109092 4020 109098 4072
rect 110966 4060 110972 4072
rect 110927 4032 110972 4060
rect 110966 4020 110972 4032
rect 111024 4060 111030 4072
rect 111429 4063 111487 4069
rect 111429 4060 111441 4063
rect 111024 4032 111441 4060
rect 111024 4020 111030 4032
rect 111429 4029 111441 4032
rect 111475 4029 111487 4063
rect 111619 4060 111647 4168
rect 114186 4156 114192 4208
rect 114244 4196 114250 4208
rect 114244 4168 118740 4196
rect 114244 4156 114250 4168
rect 114646 4088 114652 4140
rect 114704 4128 114710 4140
rect 115566 4128 115572 4140
rect 114704 4100 115572 4128
rect 114704 4088 114710 4100
rect 115566 4088 115572 4100
rect 115624 4088 115630 4140
rect 115750 4088 115756 4140
rect 115808 4128 115814 4140
rect 118234 4128 118240 4140
rect 115808 4100 118096 4128
rect 118195 4100 118240 4128
rect 115808 4088 115814 4100
rect 113726 4060 113732 4072
rect 111619 4032 113732 4060
rect 111429 4023 111487 4029
rect 55766 3952 55772 4004
rect 55824 3992 55830 4004
rect 93026 3992 93032 4004
rect 55824 3964 60734 3992
rect 55824 3952 55830 3964
rect 54720 3896 55720 3924
rect 60369 3927 60427 3933
rect 54720 3884 54726 3896
rect 60369 3893 60381 3927
rect 60415 3924 60427 3927
rect 60458 3924 60464 3936
rect 60415 3896 60464 3924
rect 60415 3893 60427 3896
rect 60369 3887 60427 3893
rect 60458 3884 60464 3896
rect 60516 3884 60522 3936
rect 60706 3924 60734 3964
rect 80026 3964 93032 3992
rect 66254 3924 66260 3936
rect 60706 3896 66260 3924
rect 66254 3884 66260 3896
rect 66312 3884 66318 3936
rect 74810 3924 74816 3936
rect 74771 3896 74816 3924
rect 74810 3884 74816 3896
rect 74868 3884 74874 3936
rect 79597 3927 79655 3933
rect 79597 3893 79609 3927
rect 79643 3924 79655 3927
rect 80026 3924 80054 3964
rect 93026 3952 93032 3964
rect 93084 3952 93090 4004
rect 107654 3992 107660 4004
rect 105832 3964 107660 3992
rect 79643 3896 80054 3924
rect 79643 3893 79655 3896
rect 79597 3887 79655 3893
rect 84838 3884 84844 3936
rect 84896 3924 84902 3936
rect 91554 3924 91560 3936
rect 84896 3896 91560 3924
rect 84896 3884 84902 3896
rect 91554 3884 91560 3896
rect 91612 3884 91618 3936
rect 102962 3884 102968 3936
rect 103020 3924 103026 3936
rect 105832 3924 105860 3964
rect 107654 3952 107660 3964
rect 107712 3952 107718 4004
rect 109589 3995 109647 4001
rect 109589 3961 109601 3995
rect 109635 3992 109647 3995
rect 109678 3992 109684 4004
rect 109635 3964 109684 3992
rect 109635 3961 109647 3964
rect 109589 3955 109647 3961
rect 109678 3952 109684 3964
rect 109736 3952 109742 4004
rect 105998 3924 106004 3936
rect 103020 3896 105860 3924
rect 105959 3896 106004 3924
rect 103020 3884 103026 3896
rect 105998 3884 106004 3896
rect 106056 3884 106062 3936
rect 111444 3924 111472 4023
rect 113726 4020 113732 4032
rect 113784 4020 113790 4072
rect 116762 4020 116768 4072
rect 116820 4060 116826 4072
rect 118068 4060 118096 4100
rect 118234 4088 118240 4100
rect 118292 4088 118298 4140
rect 118418 4128 118424 4140
rect 118379 4100 118424 4128
rect 118418 4088 118424 4100
rect 118476 4088 118482 4140
rect 118602 4128 118608 4140
rect 118563 4100 118608 4128
rect 118602 4088 118608 4100
rect 118660 4088 118666 4140
rect 118712 4128 118740 4168
rect 119154 4156 119160 4208
rect 119212 4196 119218 4208
rect 119249 4199 119307 4205
rect 119249 4196 119261 4199
rect 119212 4168 119261 4196
rect 119212 4156 119218 4168
rect 119249 4165 119261 4168
rect 119295 4165 119307 4199
rect 128170 4196 128176 4208
rect 119249 4159 119307 4165
rect 119632 4168 128176 4196
rect 119632 4128 119660 4168
rect 128170 4156 128176 4168
rect 128228 4156 128234 4208
rect 128262 4156 128268 4208
rect 128320 4196 128326 4208
rect 128817 4199 128875 4205
rect 128817 4196 128829 4199
rect 128320 4168 128829 4196
rect 128320 4156 128326 4168
rect 128817 4165 128829 4168
rect 128863 4196 128875 4199
rect 131666 4196 131672 4208
rect 128863 4168 130424 4196
rect 128863 4165 128875 4168
rect 128817 4159 128875 4165
rect 118712 4100 119660 4128
rect 120905 4131 120963 4137
rect 120905 4097 120917 4131
rect 120951 4128 120963 4131
rect 121457 4131 121515 4137
rect 121457 4128 121469 4131
rect 120951 4100 121469 4128
rect 120951 4097 120963 4100
rect 120905 4091 120963 4097
rect 121457 4097 121469 4100
rect 121503 4128 121515 4131
rect 122742 4128 122748 4140
rect 121503 4100 122748 4128
rect 121503 4097 121515 4100
rect 121457 4091 121515 4097
rect 122742 4088 122748 4100
rect 122800 4088 122806 4140
rect 122834 4088 122840 4140
rect 122892 4128 122898 4140
rect 123294 4128 123300 4140
rect 122892 4100 123300 4128
rect 122892 4088 122898 4100
rect 123294 4088 123300 4100
rect 123352 4088 123358 4140
rect 123593 4131 123651 4137
rect 123593 4097 123605 4131
rect 123639 4128 123651 4131
rect 123849 4131 123907 4137
rect 123639 4100 123800 4128
rect 123639 4097 123651 4100
rect 123593 4091 123651 4097
rect 123772 4060 123800 4100
rect 123849 4097 123861 4131
rect 123895 4128 123907 4131
rect 123938 4128 123944 4140
rect 123895 4100 123944 4128
rect 123895 4097 123907 4100
rect 123849 4091 123907 4097
rect 123938 4088 123944 4100
rect 123996 4128 124002 4140
rect 124309 4131 124367 4137
rect 124309 4128 124321 4131
rect 123996 4100 124321 4128
rect 123996 4088 124002 4100
rect 124309 4097 124321 4100
rect 124355 4097 124367 4131
rect 125226 4128 125232 4140
rect 125187 4100 125232 4128
rect 124309 4091 124367 4097
rect 125226 4088 125232 4100
rect 125284 4088 125290 4140
rect 125318 4088 125324 4140
rect 125376 4128 125382 4140
rect 126057 4131 126115 4137
rect 126057 4128 126069 4131
rect 125376 4100 126069 4128
rect 125376 4088 125382 4100
rect 126057 4097 126069 4100
rect 126103 4097 126115 4131
rect 126057 4091 126115 4097
rect 126146 4088 126152 4140
rect 126204 4128 126210 4140
rect 126324 4131 126382 4137
rect 126324 4128 126336 4131
rect 126204 4100 126336 4128
rect 126204 4088 126210 4100
rect 126324 4097 126336 4100
rect 126370 4128 126382 4131
rect 126370 4100 127940 4128
rect 126370 4097 126382 4100
rect 126324 4091 126382 4097
rect 125413 4063 125471 4069
rect 116820 4032 118004 4060
rect 118068 4032 122880 4060
rect 123772 4032 123984 4060
rect 116820 4020 116826 4032
rect 111610 3952 111616 4004
rect 111668 3992 111674 4004
rect 117976 3992 118004 4032
rect 118970 3992 118976 4004
rect 111668 3964 117912 3992
rect 117976 3964 118976 3992
rect 111668 3952 111674 3964
rect 117774 3924 117780 3936
rect 111444 3896 117780 3924
rect 117774 3884 117780 3896
rect 117832 3884 117838 3936
rect 117884 3924 117912 3964
rect 118970 3952 118976 3964
rect 119028 3992 119034 4004
rect 120994 3992 121000 4004
rect 119028 3964 121000 3992
rect 119028 3952 119034 3964
rect 120994 3952 121000 3964
rect 121052 3952 121058 4004
rect 122469 3995 122527 4001
rect 122469 3961 122481 3995
rect 122515 3992 122527 3995
rect 122742 3992 122748 4004
rect 122515 3964 122748 3992
rect 122515 3961 122527 3964
rect 122469 3955 122527 3961
rect 122742 3952 122748 3964
rect 122800 3952 122806 4004
rect 119157 3927 119215 3933
rect 119157 3924 119169 3927
rect 117884 3896 119169 3924
rect 119157 3893 119169 3896
rect 119203 3893 119215 3927
rect 119157 3887 119215 3893
rect 119246 3884 119252 3936
rect 119304 3924 119310 3936
rect 119893 3927 119951 3933
rect 119893 3924 119905 3927
rect 119304 3896 119905 3924
rect 119304 3884 119310 3896
rect 119893 3893 119905 3896
rect 119939 3924 119951 3927
rect 120074 3924 120080 3936
rect 119939 3896 120080 3924
rect 119939 3893 119951 3896
rect 119893 3887 119951 3893
rect 120074 3884 120080 3896
rect 120132 3924 120138 3936
rect 121178 3924 121184 3936
rect 120132 3896 121184 3924
rect 120132 3884 120138 3896
rect 121178 3884 121184 3896
rect 121236 3884 121242 3936
rect 122006 3924 122012 3936
rect 121967 3896 122012 3924
rect 122006 3884 122012 3896
rect 122064 3884 122070 3936
rect 122852 3924 122880 4032
rect 123956 3992 123984 4032
rect 125413 4029 125425 4063
rect 125459 4060 125471 4063
rect 125502 4060 125508 4072
rect 125459 4032 125508 4060
rect 125459 4029 125471 4032
rect 125413 4023 125471 4029
rect 125502 4020 125508 4032
rect 125560 4020 125566 4072
rect 127912 4069 127940 4100
rect 127986 4088 127992 4140
rect 128044 4128 128050 4140
rect 130396 4128 130424 4168
rect 131224 4168 131672 4196
rect 131224 4128 131252 4168
rect 131666 4156 131672 4168
rect 131724 4156 131730 4208
rect 133064 4196 133092 4236
rect 133230 4224 133236 4276
rect 133288 4264 133294 4276
rect 140130 4264 140136 4276
rect 133288 4236 140136 4264
rect 133288 4224 133294 4236
rect 140130 4224 140136 4236
rect 140188 4224 140194 4276
rect 141142 4264 141148 4276
rect 141103 4236 141148 4264
rect 141142 4224 141148 4236
rect 141200 4224 141206 4276
rect 157242 4264 157248 4276
rect 144779 4236 157248 4264
rect 137922 4196 137928 4208
rect 133064 4168 137928 4196
rect 137922 4156 137928 4168
rect 137980 4156 137986 4208
rect 143350 4196 143356 4208
rect 142816 4168 143356 4196
rect 128044 4100 130332 4128
rect 130396 4100 131252 4128
rect 131321 4131 131379 4137
rect 128044 4088 128050 4100
rect 127897 4063 127955 4069
rect 127897 4029 127909 4063
rect 127943 4060 127955 4063
rect 129918 4060 129924 4072
rect 127943 4032 129924 4060
rect 127943 4029 127955 4032
rect 127897 4023 127955 4029
rect 129918 4020 129924 4032
rect 129976 4020 129982 4072
rect 126054 3992 126060 4004
rect 123956 3964 126060 3992
rect 126054 3952 126060 3964
rect 126112 3952 126118 4004
rect 127434 3992 127440 4004
rect 127395 3964 127440 3992
rect 127434 3952 127440 3964
rect 127492 3952 127498 4004
rect 130197 3995 130255 4001
rect 130197 3992 130209 3995
rect 127544 3964 130209 3992
rect 127544 3924 127572 3964
rect 130197 3961 130209 3964
rect 130243 3961 130255 3995
rect 130197 3955 130255 3961
rect 122852 3896 127572 3924
rect 127618 3884 127624 3936
rect 127676 3924 127682 3936
rect 127986 3924 127992 3936
rect 127676 3896 127992 3924
rect 127676 3884 127682 3896
rect 127986 3884 127992 3896
rect 128044 3884 128050 3936
rect 128998 3884 129004 3936
rect 129056 3924 129062 3936
rect 129277 3927 129335 3933
rect 129277 3924 129289 3927
rect 129056 3896 129289 3924
rect 129056 3884 129062 3896
rect 129277 3893 129289 3896
rect 129323 3893 129335 3927
rect 130304 3924 130332 4100
rect 131321 4097 131333 4131
rect 131367 4128 131379 4131
rect 131758 4128 131764 4140
rect 131367 4100 131764 4128
rect 131367 4097 131379 4100
rect 131321 4091 131379 4097
rect 131758 4088 131764 4100
rect 131816 4088 131822 4140
rect 138290 4137 138296 4140
rect 133161 4131 133219 4137
rect 133161 4097 133173 4131
rect 133207 4128 133219 4131
rect 133207 4100 135576 4128
rect 133207 4097 133219 4100
rect 133161 4091 133219 4097
rect 131577 4063 131635 4069
rect 131577 4029 131589 4063
rect 131623 4060 131635 4063
rect 132034 4060 132040 4072
rect 131623 4032 132040 4060
rect 131623 4029 131635 4032
rect 131577 4023 131635 4029
rect 132034 4020 132040 4032
rect 132092 4020 132098 4072
rect 133417 4063 133475 4069
rect 133417 4029 133429 4063
rect 133463 4060 133475 4063
rect 133598 4060 133604 4072
rect 133463 4032 133604 4060
rect 133463 4029 133475 4032
rect 133417 4023 133475 4029
rect 133598 4020 133604 4032
rect 133656 4020 133662 4072
rect 133966 4020 133972 4072
rect 134024 4060 134030 4072
rect 134153 4063 134211 4069
rect 134153 4060 134165 4063
rect 134024 4032 134165 4060
rect 134024 4020 134030 4032
rect 134153 4029 134165 4032
rect 134199 4060 134211 4063
rect 134242 4060 134248 4072
rect 134199 4032 134248 4060
rect 134199 4029 134211 4032
rect 134153 4023 134211 4029
rect 134242 4020 134248 4032
rect 134300 4020 134306 4072
rect 134797 4063 134855 4069
rect 134797 4029 134809 4063
rect 134843 4060 134855 4063
rect 134978 4060 134984 4072
rect 134843 4032 134984 4060
rect 134843 4029 134855 4032
rect 134797 4023 134855 4029
rect 134978 4020 134984 4032
rect 135036 4020 135042 4072
rect 131758 3952 131764 4004
rect 131816 3992 131822 4004
rect 131816 3964 132540 3992
rect 131816 3952 131822 3964
rect 132037 3927 132095 3933
rect 132037 3924 132049 3927
rect 130304 3896 132049 3924
rect 129277 3887 129335 3893
rect 132037 3893 132049 3896
rect 132083 3893 132095 3927
rect 132512 3924 132540 3964
rect 135254 3924 135260 3936
rect 132512 3896 135260 3924
rect 132037 3887 132095 3893
rect 135254 3884 135260 3896
rect 135312 3884 135318 3936
rect 135548 3924 135576 4100
rect 138284 4091 138296 4137
rect 138348 4128 138354 4140
rect 138348 4100 138384 4128
rect 138290 4088 138296 4091
rect 138348 4088 138354 4100
rect 139854 4088 139860 4140
rect 139912 4128 139918 4140
rect 140314 4128 140320 4140
rect 139912 4100 140320 4128
rect 139912 4088 139918 4100
rect 140314 4088 140320 4100
rect 140372 4128 140378 4140
rect 142816 4128 142844 4168
rect 143350 4156 143356 4168
rect 143408 4156 143414 4208
rect 144779 4205 144807 4236
rect 157242 4224 157248 4236
rect 157300 4224 157306 4276
rect 144764 4199 144822 4205
rect 144764 4165 144776 4199
rect 144810 4165 144822 4199
rect 144764 4159 144822 4165
rect 145558 4156 145564 4208
rect 145616 4196 145622 4208
rect 145653 4199 145711 4205
rect 145653 4196 145665 4199
rect 145616 4168 145665 4196
rect 145616 4156 145622 4168
rect 145653 4165 145665 4168
rect 145699 4165 145711 4199
rect 145653 4159 145711 4165
rect 146662 4156 146668 4208
rect 146720 4196 146726 4208
rect 149238 4196 149244 4208
rect 146720 4168 149244 4196
rect 146720 4156 146726 4168
rect 149238 4156 149244 4168
rect 149296 4156 149302 4208
rect 149640 4199 149698 4205
rect 149640 4165 149652 4199
rect 149686 4196 149698 4199
rect 151814 4196 151820 4208
rect 149686 4168 149836 4196
rect 149686 4165 149698 4168
rect 149640 4159 149698 4165
rect 140372 4100 142844 4128
rect 140372 4088 140378 4100
rect 142890 4088 142896 4140
rect 142948 4137 142954 4140
rect 142948 4128 142960 4137
rect 144178 4128 144184 4140
rect 142948 4100 142993 4128
rect 143184 4100 144184 4128
rect 142948 4091 142960 4100
rect 142948 4088 142954 4091
rect 135714 4020 135720 4072
rect 135772 4060 135778 4072
rect 135901 4063 135959 4069
rect 135901 4060 135913 4063
rect 135772 4032 135913 4060
rect 135772 4020 135778 4032
rect 135901 4029 135913 4032
rect 135947 4029 135959 4063
rect 135901 4023 135959 4029
rect 136082 4020 136088 4072
rect 136140 4060 136146 4072
rect 136453 4063 136511 4069
rect 136453 4060 136465 4063
rect 136140 4032 136465 4060
rect 136140 4020 136146 4032
rect 136453 4029 136465 4032
rect 136499 4060 136511 4063
rect 137830 4060 137836 4072
rect 136499 4032 137836 4060
rect 136499 4029 136511 4032
rect 136453 4023 136511 4029
rect 137830 4020 137836 4032
rect 137888 4060 137894 4072
rect 143184 4069 143212 4100
rect 144178 4088 144184 4100
rect 144236 4128 144242 4140
rect 144860 4128 144914 4134
rect 145009 4131 145067 4137
rect 145009 4128 145021 4131
rect 144236 4100 145021 4128
rect 144236 4088 144242 4100
rect 145009 4097 145021 4100
rect 145055 4097 145067 4131
rect 145009 4091 145067 4097
rect 145190 4088 145196 4140
rect 145248 4128 145254 4140
rect 145837 4131 145895 4137
rect 145837 4128 145849 4131
rect 145248 4100 145849 4128
rect 145248 4088 145254 4100
rect 145837 4097 145849 4100
rect 145883 4097 145895 4131
rect 147214 4128 147220 4140
rect 145837 4091 145895 4097
rect 147048 4100 147220 4128
rect 138017 4063 138075 4069
rect 138017 4060 138029 4063
rect 137888 4032 138029 4060
rect 137888 4020 137894 4032
rect 138017 4029 138029 4032
rect 138063 4029 138075 4063
rect 138017 4023 138075 4029
rect 143169 4063 143227 4069
rect 143169 4029 143181 4063
rect 143215 4029 143227 4063
rect 143169 4023 143227 4029
rect 146021 4063 146079 4069
rect 146021 4029 146033 4063
rect 146067 4060 146079 4063
rect 147048 4060 147076 4100
rect 147214 4088 147220 4100
rect 147272 4088 147278 4140
rect 147789 4131 147847 4137
rect 147789 4097 147801 4131
rect 147835 4128 147847 4131
rect 148778 4128 148784 4140
rect 147835 4100 148784 4128
rect 147835 4097 147847 4100
rect 147789 4091 147847 4097
rect 148778 4088 148784 4100
rect 148836 4088 148842 4140
rect 148042 4060 148048 4072
rect 146067 4032 147076 4060
rect 148003 4032 148048 4060
rect 146067 4029 146079 4032
rect 146021 4023 146079 4029
rect 137005 3995 137063 4001
rect 137005 3961 137017 3995
rect 137051 3992 137063 3995
rect 137557 3995 137615 4001
rect 137557 3992 137569 3995
rect 137051 3964 137569 3992
rect 137051 3961 137063 3964
rect 137005 3955 137063 3961
rect 137557 3961 137569 3964
rect 137603 3992 137615 3995
rect 137646 3992 137652 4004
rect 137603 3964 137652 3992
rect 137603 3961 137615 3964
rect 137557 3955 137615 3961
rect 137646 3952 137652 3964
rect 137704 3952 137710 4004
rect 139394 3992 139400 4004
rect 139355 3964 139400 3992
rect 139394 3952 139400 3964
rect 139452 3952 139458 4004
rect 139946 3992 139952 4004
rect 139859 3964 139952 3992
rect 139946 3952 139952 3964
rect 140004 3992 140010 4004
rect 141050 3992 141056 4004
rect 140004 3964 141056 3992
rect 140004 3952 140010 3964
rect 141050 3952 141056 3964
rect 141108 3952 141114 4004
rect 141786 3992 141792 4004
rect 141747 3964 141792 3992
rect 141786 3952 141792 3964
rect 141844 3952 141850 4004
rect 139762 3924 139768 3936
rect 135548 3896 139768 3924
rect 139762 3884 139768 3896
rect 139820 3884 139826 3936
rect 140038 3884 140044 3936
rect 140096 3924 140102 3936
rect 140498 3924 140504 3936
rect 140096 3896 140504 3924
rect 140096 3884 140102 3896
rect 140498 3884 140504 3896
rect 140556 3884 140562 3936
rect 141418 3884 141424 3936
rect 141476 3924 141482 3936
rect 143184 3924 143212 4023
rect 145558 3952 145564 4004
rect 145616 3992 145622 4004
rect 146036 3992 146064 4023
rect 146938 3992 146944 4004
rect 145616 3964 146064 3992
rect 146496 3964 146944 3992
rect 145616 3952 145622 3964
rect 143626 3924 143632 3936
rect 141476 3896 143212 3924
rect 143587 3896 143632 3924
rect 141476 3884 141482 3896
rect 143626 3884 143632 3896
rect 143684 3924 143690 3936
rect 146496 3924 146524 3964
rect 146938 3952 146944 3964
rect 146996 3952 147002 4004
rect 146662 3924 146668 3936
rect 143684 3896 146524 3924
rect 146623 3896 146668 3924
rect 143684 3884 143690 3896
rect 146662 3884 146668 3896
rect 146720 3884 146726 3936
rect 147048 3924 147076 4032
rect 148042 4020 148048 4032
rect 148100 4020 148106 4072
rect 149808 4060 149836 4168
rect 149900 4168 151820 4196
rect 149900 4140 149928 4168
rect 151814 4156 151820 4168
rect 151872 4156 151878 4208
rect 154424 4199 154482 4205
rect 151933 4168 152228 4196
rect 149882 4088 149888 4140
rect 149940 4128 149946 4140
rect 149940 4100 150033 4128
rect 149940 4088 149946 4100
rect 151538 4088 151544 4140
rect 151596 4128 151602 4140
rect 151933 4128 151961 4168
rect 151596 4100 151961 4128
rect 151596 4088 151602 4100
rect 151998 4088 152004 4140
rect 152056 4137 152062 4140
rect 152056 4128 152068 4137
rect 152200 4128 152228 4168
rect 154424 4165 154436 4199
rect 154470 4196 154482 4199
rect 154666 4196 154672 4208
rect 154470 4168 154672 4196
rect 154470 4165 154482 4168
rect 154424 4159 154482 4165
rect 154666 4156 154672 4168
rect 154724 4156 154730 4208
rect 155144 4168 155448 4196
rect 152734 4128 152740 4140
rect 152056 4100 152101 4128
rect 152200 4100 152596 4128
rect 152695 4100 152740 4128
rect 152056 4091 152068 4100
rect 152056 4088 152062 4091
rect 150066 4060 150072 4072
rect 149808 4032 150072 4060
rect 150066 4020 150072 4032
rect 150124 4060 150130 4072
rect 151262 4060 151268 4072
rect 150124 4032 151268 4060
rect 150124 4020 150130 4032
rect 151262 4020 151268 4032
rect 151320 4020 151326 4072
rect 152277 4063 152335 4069
rect 152277 4029 152289 4063
rect 152323 4060 152335 4063
rect 152458 4060 152464 4072
rect 152323 4032 152464 4060
rect 152323 4029 152335 4032
rect 152277 4023 152335 4029
rect 152458 4020 152464 4032
rect 152516 4020 152522 4072
rect 152568 4060 152596 4100
rect 152734 4088 152740 4100
rect 152792 4088 152798 4140
rect 155144 4128 155172 4168
rect 153580 4100 155172 4128
rect 153580 4060 153608 4100
rect 155218 4088 155224 4140
rect 155276 4128 155282 4140
rect 155313 4131 155371 4137
rect 155313 4128 155325 4131
rect 155276 4100 155325 4128
rect 155276 4088 155282 4100
rect 155313 4097 155325 4100
rect 155359 4097 155371 4131
rect 155420 4128 155448 4168
rect 155957 4131 156015 4137
rect 155957 4128 155969 4131
rect 155420 4100 155969 4128
rect 155313 4091 155371 4097
rect 155957 4097 155969 4100
rect 156003 4097 156015 4131
rect 155957 4091 156015 4097
rect 156141 4131 156199 4137
rect 156141 4097 156153 4131
rect 156187 4097 156199 4131
rect 156141 4091 156199 4097
rect 156325 4131 156383 4137
rect 156325 4097 156337 4131
rect 156371 4128 156383 4131
rect 156414 4128 156420 4140
rect 156371 4100 156420 4128
rect 156371 4097 156383 4100
rect 156325 4091 156383 4097
rect 154666 4060 154672 4072
rect 152568 4032 153608 4060
rect 154627 4032 154672 4060
rect 154666 4020 154672 4032
rect 154724 4020 154730 4072
rect 156156 4060 156184 4091
rect 156414 4088 156420 4100
rect 156472 4088 156478 4140
rect 156506 4088 156512 4140
rect 156564 4128 156570 4140
rect 156969 4131 157027 4137
rect 156969 4128 156981 4131
rect 156564 4100 156981 4128
rect 156564 4088 156570 4100
rect 156969 4097 156981 4100
rect 157015 4097 157027 4131
rect 156969 4091 157027 4097
rect 157613 4131 157671 4137
rect 157613 4097 157625 4131
rect 157659 4128 157671 4131
rect 157702 4128 157708 4140
rect 157659 4100 157708 4128
rect 157659 4097 157671 4100
rect 157613 4091 157671 4097
rect 157702 4088 157708 4100
rect 157760 4088 157766 4140
rect 158254 4128 158260 4140
rect 158215 4100 158260 4128
rect 158254 4088 158260 4100
rect 158312 4088 158318 4140
rect 154776 4032 156184 4060
rect 148060 3964 148640 3992
rect 147674 3924 147680 3936
rect 147048 3896 147680 3924
rect 147674 3884 147680 3896
rect 147732 3884 147738 3936
rect 147858 3884 147864 3936
rect 147916 3924 147922 3936
rect 148060 3924 148088 3964
rect 148502 3924 148508 3936
rect 147916 3896 148088 3924
rect 148463 3896 148508 3924
rect 147916 3884 147922 3896
rect 148502 3884 148508 3896
rect 148560 3884 148566 3936
rect 148612 3924 148640 3964
rect 149900 3964 151032 3992
rect 149900 3924 149928 3964
rect 150894 3924 150900 3936
rect 148612 3896 149928 3924
rect 150855 3896 150900 3924
rect 150894 3884 150900 3896
rect 150952 3884 150958 3936
rect 151004 3924 151032 3964
rect 152292 3964 153424 3992
rect 152292 3924 152320 3964
rect 153286 3924 153292 3936
rect 151004 3896 152320 3924
rect 153247 3896 153292 3924
rect 153286 3884 153292 3896
rect 153344 3884 153350 3936
rect 153396 3924 153424 3964
rect 154776 3924 154804 4032
rect 155126 3992 155132 4004
rect 155087 3964 155132 3992
rect 155126 3952 155132 3964
rect 155184 3952 155190 4004
rect 156046 3952 156052 4004
rect 156104 3992 156110 4004
rect 158073 3995 158131 4001
rect 158073 3992 158085 3995
rect 156104 3964 158085 3992
rect 156104 3952 156110 3964
rect 158073 3961 158085 3964
rect 158119 3961 158131 3995
rect 158073 3955 158131 3961
rect 153396 3896 154804 3924
rect 154942 3884 154948 3936
rect 155000 3924 155006 3936
rect 156414 3924 156420 3936
rect 155000 3896 156420 3924
rect 155000 3884 155006 3896
rect 156414 3884 156420 3896
rect 156472 3884 156478 3936
rect 156782 3924 156788 3936
rect 156743 3896 156788 3924
rect 156782 3884 156788 3896
rect 156840 3884 156846 3936
rect 156874 3884 156880 3936
rect 156932 3924 156938 3936
rect 157429 3927 157487 3933
rect 157429 3924 157441 3927
rect 156932 3896 157441 3924
rect 156932 3884 156938 3896
rect 157429 3893 157441 3896
rect 157475 3893 157487 3927
rect 157429 3887 157487 3893
rect 1104 3834 158884 3856
rect 1104 3782 20672 3834
rect 20724 3782 20736 3834
rect 20788 3782 20800 3834
rect 20852 3782 20864 3834
rect 20916 3782 20928 3834
rect 20980 3782 60117 3834
rect 60169 3782 60181 3834
rect 60233 3782 60245 3834
rect 60297 3782 60309 3834
rect 60361 3782 60373 3834
rect 60425 3782 99562 3834
rect 99614 3782 99626 3834
rect 99678 3782 99690 3834
rect 99742 3782 99754 3834
rect 99806 3782 99818 3834
rect 99870 3782 139007 3834
rect 139059 3782 139071 3834
rect 139123 3782 139135 3834
rect 139187 3782 139199 3834
rect 139251 3782 139263 3834
rect 139315 3782 158884 3834
rect 1104 3760 158884 3782
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 13998 3720 14004 3732
rect 13311 3692 14004 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16172 3692 16681 3720
rect 16172 3680 16178 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 18877 3723 18935 3729
rect 18877 3689 18889 3723
rect 18923 3720 18935 3723
rect 20438 3720 20444 3732
rect 18923 3692 20444 3720
rect 18923 3689 18935 3692
rect 18877 3683 18935 3689
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20809 3723 20867 3729
rect 20809 3689 20821 3723
rect 20855 3720 20867 3723
rect 21818 3720 21824 3732
rect 20855 3692 21824 3720
rect 20855 3689 20867 3692
rect 20809 3683 20867 3689
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 24857 3723 24915 3729
rect 24857 3689 24869 3723
rect 24903 3720 24915 3723
rect 25222 3720 25228 3732
rect 24903 3692 25228 3720
rect 24903 3689 24915 3692
rect 24857 3683 24915 3689
rect 25222 3680 25228 3692
rect 25280 3680 25286 3732
rect 25685 3723 25743 3729
rect 25685 3689 25697 3723
rect 25731 3720 25743 3723
rect 25866 3720 25872 3732
rect 25731 3692 25872 3720
rect 25731 3689 25743 3692
rect 25685 3683 25743 3689
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 30558 3720 30564 3732
rect 30519 3692 30564 3720
rect 30558 3680 30564 3692
rect 30616 3680 30622 3732
rect 32953 3723 33011 3729
rect 32953 3720 32965 3723
rect 30668 3692 32965 3720
rect 16209 3655 16267 3661
rect 16209 3621 16221 3655
rect 16255 3652 16267 3655
rect 16298 3652 16304 3664
rect 16255 3624 16304 3652
rect 16255 3621 16267 3624
rect 16209 3615 16267 3621
rect 16298 3612 16304 3624
rect 16356 3612 16362 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21634 3652 21640 3664
rect 20772 3624 21640 3652
rect 20772 3612 20778 3624
rect 21634 3612 21640 3624
rect 21692 3612 21698 3664
rect 24762 3612 24768 3664
rect 24820 3652 24826 3664
rect 30668 3652 30696 3692
rect 32953 3689 32965 3692
rect 32999 3689 33011 3723
rect 32953 3683 33011 3689
rect 36906 3680 36912 3732
rect 36964 3720 36970 3732
rect 37001 3723 37059 3729
rect 37001 3720 37013 3723
rect 36964 3692 37013 3720
rect 36964 3680 36970 3692
rect 37001 3689 37013 3692
rect 37047 3689 37059 3723
rect 37001 3683 37059 3689
rect 37182 3680 37188 3732
rect 37240 3720 37246 3732
rect 45462 3720 45468 3732
rect 37240 3692 45468 3720
rect 37240 3680 37246 3692
rect 45462 3680 45468 3692
rect 45520 3680 45526 3732
rect 49789 3723 49847 3729
rect 45572 3692 49740 3720
rect 24820 3624 30696 3652
rect 32493 3655 32551 3661
rect 24820 3612 24826 3624
rect 32493 3621 32505 3655
rect 32539 3652 32551 3655
rect 32582 3652 32588 3664
rect 32539 3624 32588 3652
rect 32539 3621 32551 3624
rect 32493 3615 32551 3621
rect 32582 3612 32588 3624
rect 32640 3612 32646 3664
rect 36541 3655 36599 3661
rect 36541 3621 36553 3655
rect 36587 3652 36599 3655
rect 37366 3652 37372 3664
rect 36587 3624 37372 3652
rect 36587 3621 36599 3624
rect 36541 3615 36599 3621
rect 37366 3612 37372 3624
rect 37424 3652 37430 3664
rect 37734 3652 37740 3664
rect 37424 3624 37740 3652
rect 37424 3612 37430 3624
rect 37734 3612 37740 3624
rect 37792 3612 37798 3664
rect 45186 3652 45192 3664
rect 45147 3624 45192 3652
rect 45186 3612 45192 3624
rect 45244 3612 45250 3664
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 31110 3584 31116 3596
rect 13320 3556 17632 3584
rect 13320 3544 13326 3556
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 13998 3408 14004 3460
rect 14056 3448 14062 3460
rect 14568 3448 14596 3479
rect 16666 3476 16672 3528
rect 16724 3516 16730 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16724 3488 16865 3516
rect 16724 3476 16730 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17604 3516 17632 3556
rect 23676 3556 25636 3584
rect 31071 3556 31116 3584
rect 17604 3488 18092 3516
rect 17497 3479 17555 3485
rect 14056 3420 14596 3448
rect 14056 3408 14062 3420
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16960 3448 16988 3479
rect 16356 3420 16988 3448
rect 16356 3408 16362 3420
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14277 3383 14335 3389
rect 14277 3380 14289 3383
rect 13596 3352 14289 3380
rect 13596 3340 13602 3352
rect 14277 3349 14289 3352
rect 14323 3349 14335 3383
rect 15562 3380 15568 3392
rect 15523 3352 15568 3380
rect 14277 3343 14335 3349
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 17512 3380 17540 3479
rect 17586 3408 17592 3460
rect 17644 3448 17650 3460
rect 17742 3451 17800 3457
rect 17742 3448 17754 3451
rect 17644 3420 17754 3448
rect 17644 3408 17650 3420
rect 17742 3417 17754 3420
rect 17788 3417 17800 3451
rect 17742 3411 17800 3417
rect 17954 3380 17960 3392
rect 17512 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18064 3380 18092 3488
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18506 3516 18512 3528
rect 18288 3488 18512 3516
rect 18288 3476 18294 3488
rect 18506 3476 18512 3488
rect 18564 3516 18570 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18564 3488 19441 3516
rect 18564 3476 18570 3488
rect 19429 3485 19441 3488
rect 19475 3516 19487 3519
rect 20070 3516 20076 3528
rect 19475 3488 20076 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 20070 3476 20076 3488
rect 20128 3516 20134 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20128 3488 21281 3516
rect 20128 3476 20134 3488
rect 21269 3485 21281 3488
rect 21315 3516 21327 3519
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21315 3488 21925 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21913 3485 21925 3488
rect 21959 3516 21971 3519
rect 22554 3516 22560 3528
rect 21959 3488 22560 3516
rect 21959 3485 21971 3488
rect 21913 3479 21971 3485
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 19674 3451 19732 3457
rect 19674 3448 19686 3451
rect 18472 3420 19686 3448
rect 18472 3408 18478 3420
rect 19674 3417 19686 3420
rect 19720 3417 19732 3451
rect 19674 3411 19732 3417
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 22158 3451 22216 3457
rect 22158 3448 22170 3451
rect 19944 3420 22170 3448
rect 19944 3408 19950 3420
rect 22158 3417 22170 3420
rect 22204 3417 22216 3451
rect 22158 3411 22216 3417
rect 23676 3380 23704 3556
rect 25222 3476 25228 3528
rect 25280 3516 25286 3528
rect 25317 3519 25375 3525
rect 25317 3516 25329 3519
rect 25280 3488 25329 3516
rect 25280 3476 25286 3488
rect 25317 3485 25329 3488
rect 25363 3485 25375 3519
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 25317 3479 25375 3485
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 25608 3516 25636 3556
rect 31110 3544 31116 3556
rect 31168 3544 31174 3596
rect 45572 3584 45600 3692
rect 49712 3652 49740 3692
rect 49789 3689 49801 3723
rect 49835 3720 49847 3723
rect 50890 3720 50896 3732
rect 49835 3692 50896 3720
rect 49835 3689 49847 3692
rect 49789 3683 49847 3689
rect 50890 3680 50896 3692
rect 50948 3680 50954 3732
rect 62114 3720 62120 3732
rect 59004 3692 62120 3720
rect 49712 3624 50200 3652
rect 34256 3556 45600 3584
rect 34256 3516 34284 3556
rect 25608 3488 34284 3516
rect 34330 3476 34336 3528
rect 34388 3516 34394 3528
rect 34388 3488 34433 3516
rect 34388 3476 34394 3488
rect 37182 3476 37188 3528
rect 37240 3516 37246 3528
rect 37366 3516 37372 3528
rect 37240 3488 37285 3516
rect 37327 3488 37372 3516
rect 37240 3476 37246 3488
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 46566 3516 46572 3528
rect 46527 3488 46572 3516
rect 46566 3476 46572 3488
rect 46624 3476 46630 3528
rect 48409 3519 48467 3525
rect 48409 3485 48421 3519
rect 48455 3516 48467 3519
rect 48455 3488 49832 3516
rect 48455 3485 48467 3488
rect 48409 3479 48467 3485
rect 31369 3451 31427 3457
rect 31369 3448 31381 3451
rect 31312 3420 31381 3448
rect 18064 3352 23704 3380
rect 23845 3383 23903 3389
rect 23845 3349 23857 3383
rect 23891 3380 23903 3383
rect 24394 3380 24400 3392
rect 23891 3352 24400 3380
rect 23891 3349 23903 3352
rect 23845 3343 23903 3349
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 30558 3340 30564 3392
rect 30616 3380 30622 3392
rect 31312 3380 31340 3420
rect 31369 3417 31381 3420
rect 31415 3417 31427 3451
rect 31369 3411 31427 3417
rect 32858 3408 32864 3460
rect 32916 3448 32922 3460
rect 34066 3451 34124 3457
rect 34066 3448 34078 3451
rect 32916 3420 34078 3448
rect 32916 3408 32922 3420
rect 34066 3417 34078 3420
rect 34112 3417 34124 3451
rect 34066 3411 34124 3417
rect 30616 3352 31340 3380
rect 30616 3340 30622 3352
rect 33778 3340 33784 3392
rect 33836 3380 33842 3392
rect 34348 3380 34376 3476
rect 37200 3448 37228 3476
rect 37829 3451 37887 3457
rect 37829 3448 37841 3451
rect 37200 3420 37841 3448
rect 37829 3417 37841 3420
rect 37875 3417 37887 3451
rect 46302 3451 46360 3457
rect 46302 3448 46314 3451
rect 37829 3411 37887 3417
rect 44560 3420 46314 3448
rect 33836 3352 34376 3380
rect 33836 3340 33842 3352
rect 37918 3340 37924 3392
rect 37976 3380 37982 3392
rect 44560 3389 44588 3420
rect 46302 3417 46314 3420
rect 46348 3417 46360 3451
rect 46302 3411 46360 3417
rect 48676 3451 48734 3457
rect 48676 3417 48688 3451
rect 48722 3448 48734 3451
rect 49694 3448 49700 3460
rect 48722 3420 49700 3448
rect 48722 3417 48734 3420
rect 48676 3411 48734 3417
rect 49694 3408 49700 3420
rect 49752 3408 49758 3460
rect 49804 3448 49832 3488
rect 50172 3448 50200 3624
rect 52362 3544 52368 3596
rect 52420 3584 52426 3596
rect 57238 3584 57244 3596
rect 52420 3556 57244 3584
rect 52420 3544 52426 3556
rect 57238 3544 57244 3556
rect 57296 3544 57302 3596
rect 58526 3584 58532 3596
rect 58487 3556 58532 3584
rect 58526 3544 58532 3556
rect 58584 3584 58590 3596
rect 58710 3584 58716 3596
rect 58584 3556 58716 3584
rect 58584 3544 58590 3556
rect 58710 3544 58716 3556
rect 58768 3584 58774 3596
rect 59004 3593 59032 3692
rect 62114 3680 62120 3692
rect 62172 3680 62178 3732
rect 63037 3723 63095 3729
rect 63037 3689 63049 3723
rect 63083 3720 63095 3723
rect 63494 3720 63500 3732
rect 63083 3692 63500 3720
rect 63083 3689 63095 3692
rect 63037 3683 63095 3689
rect 63494 3680 63500 3692
rect 63552 3720 63558 3732
rect 64598 3720 64604 3732
rect 63552 3692 64604 3720
rect 63552 3680 63558 3692
rect 64598 3680 64604 3692
rect 64656 3680 64662 3732
rect 64874 3720 64880 3732
rect 64835 3692 64880 3720
rect 64874 3680 64880 3692
rect 64932 3680 64938 3732
rect 73154 3720 73160 3732
rect 73115 3692 73160 3720
rect 73154 3680 73160 3692
rect 73212 3680 73218 3732
rect 77110 3680 77116 3732
rect 77168 3720 77174 3732
rect 88426 3720 88432 3732
rect 77168 3692 77524 3720
rect 88387 3692 88432 3720
rect 77168 3680 77174 3692
rect 59170 3612 59176 3664
rect 59228 3652 59234 3664
rect 72605 3655 72663 3661
rect 72605 3652 72617 3655
rect 59228 3624 72617 3652
rect 59228 3612 59234 3624
rect 72605 3621 72617 3624
rect 72651 3621 72663 3655
rect 72605 3615 72663 3621
rect 58989 3587 59047 3593
rect 58989 3584 59001 3587
rect 58768 3556 59001 3584
rect 58768 3544 58774 3556
rect 58989 3553 59001 3556
rect 59035 3553 59047 3587
rect 58989 3547 59047 3553
rect 53742 3516 53748 3528
rect 53703 3488 53748 3516
rect 53742 3476 53748 3488
rect 53800 3476 53806 3528
rect 58273 3519 58331 3525
rect 58273 3485 58285 3519
rect 58319 3516 58331 3519
rect 58434 3516 58440 3528
rect 58319 3488 58440 3516
rect 58319 3485 58331 3488
rect 58273 3479 58331 3485
rect 58434 3476 58440 3488
rect 58492 3476 58498 3528
rect 61289 3519 61347 3525
rect 61289 3485 61301 3519
rect 61335 3516 61347 3519
rect 62393 3519 62451 3525
rect 62393 3516 62405 3519
rect 61335 3488 62405 3516
rect 61335 3485 61347 3488
rect 61289 3479 61347 3485
rect 62393 3485 62405 3488
rect 62439 3485 62451 3519
rect 62393 3479 62451 3485
rect 65061 3519 65119 3525
rect 65061 3485 65073 3519
rect 65107 3516 65119 3519
rect 65794 3516 65800 3528
rect 65107 3488 65800 3516
rect 65107 3485 65119 3488
rect 65061 3479 65119 3485
rect 61304 3448 61332 3479
rect 62022 3448 62028 3460
rect 49804 3420 49924 3448
rect 50172 3420 61332 3448
rect 61983 3420 62028 3448
rect 44545 3383 44603 3389
rect 44545 3380 44557 3383
rect 37976 3352 44557 3380
rect 37976 3340 37982 3352
rect 44545 3349 44557 3352
rect 44591 3349 44603 3383
rect 44545 3343 44603 3349
rect 46842 3340 46848 3392
rect 46900 3380 46906 3392
rect 49602 3380 49608 3392
rect 46900 3352 49608 3380
rect 46900 3340 46906 3352
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 49896 3380 49924 3420
rect 62022 3408 62028 3420
rect 62080 3408 62086 3460
rect 62408 3448 62436 3479
rect 65794 3476 65800 3488
rect 65852 3476 65858 3528
rect 72620 3516 72648 3615
rect 77496 3593 77524 3692
rect 88426 3680 88432 3692
rect 88484 3720 88490 3732
rect 94498 3720 94504 3732
rect 88484 3692 90404 3720
rect 94459 3692 94504 3720
rect 88484 3680 88490 3692
rect 80238 3612 80244 3664
rect 80296 3652 80302 3664
rect 88981 3655 89039 3661
rect 88981 3652 88993 3655
rect 80296 3624 88993 3652
rect 80296 3612 80302 3624
rect 88981 3621 88993 3624
rect 89027 3621 89039 3655
rect 88981 3615 89039 3621
rect 90376 3593 90404 3692
rect 94498 3680 94504 3692
rect 94556 3680 94562 3732
rect 96801 3723 96859 3729
rect 96801 3689 96813 3723
rect 96847 3720 96859 3723
rect 101861 3723 101919 3729
rect 96847 3692 101812 3720
rect 96847 3689 96859 3692
rect 96801 3683 96859 3689
rect 77481 3587 77539 3593
rect 77481 3553 77493 3587
rect 77527 3553 77539 3587
rect 77481 3547 77539 3553
rect 90361 3587 90419 3593
rect 90361 3553 90373 3587
rect 90407 3553 90419 3587
rect 96816 3584 96844 3683
rect 98733 3655 98791 3661
rect 98733 3621 98745 3655
rect 98779 3652 98791 3655
rect 99006 3652 99012 3664
rect 98779 3624 99012 3652
rect 98779 3621 98791 3624
rect 98733 3615 98791 3621
rect 99006 3612 99012 3624
rect 99064 3612 99070 3664
rect 101784 3652 101812 3692
rect 101861 3689 101873 3723
rect 101907 3720 101919 3723
rect 102042 3720 102048 3732
rect 101907 3692 102048 3720
rect 101907 3689 101919 3692
rect 101861 3683 101919 3689
rect 102042 3680 102048 3692
rect 102100 3680 102106 3732
rect 108206 3720 108212 3732
rect 102152 3692 108212 3720
rect 102152 3652 102180 3692
rect 108206 3680 108212 3692
rect 108264 3680 108270 3732
rect 113910 3680 113916 3732
rect 113968 3720 113974 3732
rect 115385 3723 115443 3729
rect 115385 3720 115397 3723
rect 113968 3692 115397 3720
rect 113968 3680 113974 3692
rect 115385 3689 115397 3692
rect 115431 3689 115443 3723
rect 115385 3683 115443 3689
rect 117958 3680 117964 3732
rect 118016 3720 118022 3732
rect 119617 3723 119675 3729
rect 119617 3720 119629 3723
rect 118016 3692 119629 3720
rect 118016 3680 118022 3692
rect 119617 3689 119629 3692
rect 119663 3689 119675 3723
rect 121917 3723 121975 3729
rect 119617 3683 119675 3689
rect 119724 3692 121040 3720
rect 101784 3624 102180 3652
rect 90361 3547 90419 3553
rect 95804 3556 96844 3584
rect 103241 3587 103299 3593
rect 74270 3519 74328 3525
rect 74270 3516 74282 3519
rect 72620 3488 74282 3516
rect 74270 3485 74282 3488
rect 74316 3485 74328 3519
rect 74534 3516 74540 3528
rect 74495 3488 74540 3516
rect 74270 3479 74328 3485
rect 74534 3476 74540 3488
rect 74592 3476 74598 3528
rect 90105 3519 90163 3525
rect 90105 3485 90117 3519
rect 90151 3516 90163 3519
rect 90542 3516 90548 3528
rect 90151 3488 90548 3516
rect 90151 3485 90163 3488
rect 90105 3479 90163 3485
rect 90542 3476 90548 3488
rect 90600 3476 90606 3528
rect 95625 3519 95683 3525
rect 95625 3485 95637 3519
rect 95671 3516 95683 3519
rect 95804 3516 95832 3556
rect 103241 3553 103253 3587
rect 103287 3584 103299 3587
rect 105170 3584 105176 3596
rect 103287 3556 105176 3584
rect 103287 3553 103299 3556
rect 103241 3547 103299 3553
rect 105170 3544 105176 3556
rect 105228 3544 105234 3596
rect 110141 3587 110199 3593
rect 110141 3584 110153 3587
rect 109972 3556 110153 3584
rect 95671 3488 95832 3516
rect 95881 3519 95939 3525
rect 95671 3485 95683 3488
rect 95625 3479 95683 3485
rect 95881 3485 95893 3519
rect 95927 3516 95939 3519
rect 96246 3516 96252 3528
rect 95927 3488 96252 3516
rect 95927 3485 95939 3488
rect 95881 3479 95939 3485
rect 96246 3476 96252 3488
rect 96304 3516 96310 3528
rect 100113 3519 100171 3525
rect 100113 3516 100125 3519
rect 96304 3488 100125 3516
rect 96304 3476 96310 3488
rect 100113 3485 100125 3488
rect 100159 3516 100171 3519
rect 100665 3519 100723 3525
rect 100665 3516 100677 3519
rect 100159 3488 100677 3516
rect 100159 3485 100171 3488
rect 100113 3479 100171 3485
rect 100665 3485 100677 3488
rect 100711 3516 100723 3519
rect 109034 3516 109040 3528
rect 100711 3488 109040 3516
rect 100711 3485 100723 3488
rect 100665 3479 100723 3485
rect 109034 3476 109040 3488
rect 109092 3516 109098 3528
rect 109586 3516 109592 3528
rect 109092 3488 109592 3516
rect 109092 3476 109098 3488
rect 109586 3476 109592 3488
rect 109644 3516 109650 3528
rect 109681 3519 109739 3525
rect 109681 3516 109693 3519
rect 109644 3488 109693 3516
rect 109644 3476 109650 3488
rect 109681 3485 109693 3488
rect 109727 3516 109739 3519
rect 109972 3516 110000 3556
rect 110141 3553 110153 3556
rect 110187 3584 110199 3587
rect 110693 3587 110751 3593
rect 110693 3584 110705 3587
rect 110187 3556 110705 3584
rect 110187 3553 110199 3556
rect 110141 3547 110199 3553
rect 110693 3553 110705 3556
rect 110739 3584 110751 3587
rect 110966 3584 110972 3596
rect 110739 3556 110972 3584
rect 110739 3553 110751 3556
rect 110693 3547 110751 3553
rect 110966 3544 110972 3556
rect 111024 3544 111030 3596
rect 116762 3584 116768 3596
rect 116723 3556 116768 3584
rect 116762 3544 116768 3556
rect 116820 3544 116826 3596
rect 119724 3584 119752 3692
rect 121012 3652 121040 3692
rect 121917 3689 121929 3723
rect 121963 3720 121975 3723
rect 126146 3720 126152 3732
rect 121963 3692 126152 3720
rect 121963 3689 121975 3692
rect 121917 3683 121975 3689
rect 126146 3680 126152 3692
rect 126204 3680 126210 3732
rect 126701 3723 126759 3729
rect 126701 3689 126713 3723
rect 126747 3720 126759 3723
rect 126882 3720 126888 3732
rect 126747 3692 126888 3720
rect 126747 3689 126759 3692
rect 126701 3683 126759 3689
rect 126882 3680 126888 3692
rect 126940 3680 126946 3732
rect 127621 3723 127679 3729
rect 127621 3689 127633 3723
rect 127667 3720 127679 3723
rect 127894 3720 127900 3732
rect 127667 3692 127900 3720
rect 127667 3689 127679 3692
rect 127621 3683 127679 3689
rect 127894 3680 127900 3692
rect 127952 3680 127958 3732
rect 127986 3680 127992 3732
rect 128044 3720 128050 3732
rect 138750 3720 138756 3732
rect 128044 3692 138756 3720
rect 128044 3680 128050 3692
rect 138750 3680 138756 3692
rect 138808 3680 138814 3732
rect 140409 3723 140467 3729
rect 138860 3692 139900 3720
rect 123018 3652 123024 3664
rect 121012 3624 123024 3652
rect 123018 3612 123024 3624
rect 123076 3612 123082 3664
rect 125505 3655 125563 3661
rect 125505 3621 125517 3655
rect 125551 3621 125563 3655
rect 125505 3615 125563 3621
rect 120994 3584 121000 3596
rect 118988 3556 119752 3584
rect 120955 3556 121000 3584
rect 109727 3488 110000 3516
rect 109727 3485 109739 3488
rect 109681 3479 109739 3485
rect 110046 3476 110052 3528
rect 110104 3516 110110 3528
rect 117774 3516 117780 3528
rect 110104 3488 117084 3516
rect 117687 3488 117780 3516
rect 110104 3476 110110 3488
rect 67542 3448 67548 3460
rect 62408 3420 67548 3448
rect 67542 3408 67548 3420
rect 67600 3408 67606 3460
rect 74442 3408 74448 3460
rect 74500 3448 74506 3460
rect 77214 3451 77272 3457
rect 77214 3448 77226 3451
rect 74500 3420 77226 3448
rect 74500 3408 74506 3420
rect 77214 3417 77226 3420
rect 77260 3448 77272 3451
rect 77941 3451 77999 3457
rect 77941 3448 77953 3451
rect 77260 3420 77953 3448
rect 77260 3417 77272 3420
rect 77214 3411 77272 3417
rect 77941 3417 77953 3420
rect 77987 3448 77999 3451
rect 84838 3448 84844 3460
rect 77987 3420 84844 3448
rect 77987 3417 77999 3420
rect 77941 3411 77999 3417
rect 84838 3408 84844 3420
rect 84896 3408 84902 3460
rect 99868 3451 99926 3457
rect 99868 3417 99880 3451
rect 99914 3448 99926 3451
rect 99914 3420 102916 3448
rect 99914 3417 99926 3420
rect 99868 3411 99926 3417
rect 51074 3380 51080 3392
rect 49896 3352 51080 3380
rect 51074 3340 51080 3352
rect 51132 3340 51138 3392
rect 53558 3380 53564 3392
rect 53519 3352 53564 3380
rect 53558 3340 53564 3352
rect 53616 3340 53622 3392
rect 57146 3380 57152 3392
rect 57059 3352 57152 3380
rect 57146 3340 57152 3352
rect 57204 3380 57210 3392
rect 57606 3380 57612 3392
rect 57204 3352 57612 3380
rect 57204 3340 57210 3352
rect 57606 3340 57612 3352
rect 57664 3340 57670 3392
rect 66162 3340 66168 3392
rect 66220 3380 66226 3392
rect 69198 3380 69204 3392
rect 66220 3352 69204 3380
rect 66220 3340 66226 3352
rect 69198 3340 69204 3352
rect 69256 3340 69262 3392
rect 76098 3380 76104 3392
rect 76059 3352 76104 3380
rect 76098 3340 76104 3352
rect 76156 3340 76162 3392
rect 102888 3380 102916 3420
rect 102962 3408 102968 3460
rect 103020 3457 103026 3460
rect 103020 3448 103032 3457
rect 109436 3451 109494 3457
rect 103020 3420 103065 3448
rect 103020 3411 103032 3420
rect 109436 3417 109448 3451
rect 109482 3448 109494 3451
rect 110138 3448 110144 3460
rect 109482 3420 110144 3448
rect 109482 3417 109494 3420
rect 109436 3411 109494 3417
rect 103020 3408 103026 3411
rect 110138 3408 110144 3420
rect 110196 3408 110202 3460
rect 116520 3451 116578 3457
rect 116520 3417 116532 3451
rect 116566 3448 116578 3451
rect 116946 3448 116952 3460
rect 116566 3420 116952 3448
rect 116566 3417 116578 3420
rect 116520 3411 116578 3417
rect 116946 3408 116952 3420
rect 117004 3408 117010 3460
rect 117056 3448 117084 3488
rect 117774 3476 117780 3488
rect 117832 3516 117838 3528
rect 118786 3516 118792 3528
rect 117832 3488 118792 3516
rect 117832 3476 117838 3488
rect 118786 3476 118792 3488
rect 118844 3476 118850 3528
rect 117682 3448 117688 3460
rect 117056 3420 117688 3448
rect 117682 3408 117688 3420
rect 117740 3408 117746 3460
rect 118044 3451 118102 3457
rect 118044 3417 118056 3451
rect 118090 3448 118102 3451
rect 118988 3448 119016 3556
rect 120994 3544 121000 3556
rect 121052 3544 121058 3596
rect 122926 3544 122932 3596
rect 122984 3584 122990 3596
rect 123294 3584 123300 3596
rect 122984 3556 123300 3584
rect 122984 3544 122990 3556
rect 123294 3544 123300 3556
rect 123352 3544 123358 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 123938 3584 123944 3596
rect 123536 3556 123944 3584
rect 123536 3544 123542 3556
rect 123938 3544 123944 3556
rect 123996 3544 124002 3596
rect 125520 3584 125548 3615
rect 125594 3612 125600 3664
rect 125652 3652 125658 3664
rect 129458 3652 129464 3664
rect 125652 3624 127848 3652
rect 129419 3624 129464 3652
rect 125652 3612 125658 3624
rect 127710 3584 127716 3596
rect 125520 3556 126836 3584
rect 119890 3476 119896 3528
rect 119948 3516 119954 3528
rect 123573 3519 123631 3525
rect 123573 3516 123585 3519
rect 119948 3488 123585 3516
rect 119948 3476 119954 3488
rect 123573 3485 123585 3488
rect 123619 3485 123631 3519
rect 123573 3479 123631 3485
rect 124125 3519 124183 3525
rect 124125 3485 124137 3519
rect 124171 3516 124183 3519
rect 125318 3516 125324 3528
rect 124171 3488 125324 3516
rect 124171 3485 124183 3488
rect 124125 3479 124183 3485
rect 120730 3451 120788 3457
rect 120730 3448 120742 3451
rect 118090 3420 119016 3448
rect 119172 3420 120742 3448
rect 118090 3417 118102 3420
rect 118044 3411 118102 3417
rect 106458 3380 106464 3392
rect 102888 3352 106464 3380
rect 106458 3340 106464 3352
rect 106516 3340 106522 3392
rect 108298 3380 108304 3392
rect 108259 3352 108304 3380
rect 108298 3340 108304 3352
rect 108356 3340 108362 3392
rect 110046 3340 110052 3392
rect 110104 3380 110110 3392
rect 111610 3380 111616 3392
rect 110104 3352 111616 3380
rect 110104 3340 110110 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 114830 3340 114836 3392
rect 114888 3380 114894 3392
rect 118234 3380 118240 3392
rect 114888 3352 118240 3380
rect 114888 3340 114894 3352
rect 118234 3340 118240 3352
rect 118292 3340 118298 3392
rect 119172 3389 119200 3420
rect 120730 3417 120742 3420
rect 120776 3448 120788 3451
rect 121270 3448 121276 3460
rect 120776 3420 121276 3448
rect 120776 3417 120788 3420
rect 120730 3411 120788 3417
rect 121270 3408 121276 3420
rect 121328 3408 121334 3460
rect 119157 3383 119215 3389
rect 119157 3349 119169 3383
rect 119203 3349 119215 3383
rect 119157 3343 119215 3349
rect 119706 3340 119712 3392
rect 119764 3380 119770 3392
rect 122469 3383 122527 3389
rect 122469 3380 122481 3383
rect 119764 3352 122481 3380
rect 119764 3340 119770 3352
rect 122469 3349 122481 3352
rect 122515 3380 122527 3383
rect 122558 3380 122564 3392
rect 122515 3352 122564 3380
rect 122515 3349 122527 3352
rect 122469 3343 122527 3349
rect 122558 3340 122564 3352
rect 122616 3340 122622 3392
rect 123018 3380 123024 3392
rect 122979 3352 123024 3380
rect 123018 3340 123024 3352
rect 123076 3340 123082 3392
rect 123588 3380 123616 3479
rect 125318 3476 125324 3488
rect 125376 3476 125382 3528
rect 125962 3516 125968 3528
rect 125428 3488 125968 3516
rect 124392 3451 124450 3457
rect 124392 3417 124404 3451
rect 124438 3448 124450 3451
rect 125428 3448 125456 3488
rect 125962 3476 125968 3488
rect 126020 3476 126026 3528
rect 124438 3420 125456 3448
rect 126808 3448 126836 3556
rect 126900 3556 127716 3584
rect 126900 3525 126928 3556
rect 127710 3544 127716 3556
rect 127768 3544 127774 3596
rect 126885 3519 126943 3525
rect 126885 3485 126897 3519
rect 126931 3485 126943 3519
rect 127066 3516 127072 3528
rect 127027 3488 127072 3516
rect 126885 3479 126943 3485
rect 127066 3476 127072 3488
rect 127124 3476 127130 3528
rect 127820 3516 127848 3624
rect 129458 3612 129464 3624
rect 129516 3612 129522 3664
rect 131022 3612 131028 3664
rect 131080 3652 131086 3664
rect 137922 3652 137928 3664
rect 131080 3624 137928 3652
rect 131080 3612 131086 3624
rect 137922 3612 137928 3624
rect 137980 3612 137986 3664
rect 138014 3612 138020 3664
rect 138072 3652 138078 3664
rect 138477 3655 138535 3661
rect 138477 3652 138489 3655
rect 138072 3624 138489 3652
rect 138072 3612 138078 3624
rect 138477 3621 138489 3624
rect 138523 3621 138535 3655
rect 138477 3615 138535 3621
rect 129734 3584 129740 3596
rect 128924 3556 129740 3584
rect 128354 3516 128360 3528
rect 127820 3488 128360 3516
rect 128354 3476 128360 3488
rect 128412 3476 128418 3528
rect 128924 3516 128952 3556
rect 129734 3544 129740 3556
rect 129792 3544 129798 3596
rect 131206 3544 131212 3596
rect 131264 3584 131270 3596
rect 131393 3587 131451 3593
rect 131393 3584 131405 3587
rect 131264 3556 131405 3584
rect 131264 3544 131270 3556
rect 131393 3553 131405 3556
rect 131439 3584 131451 3587
rect 138860 3584 138888 3692
rect 139872 3652 139900 3692
rect 140409 3689 140421 3723
rect 140455 3720 140467 3723
rect 140498 3720 140504 3732
rect 140455 3692 140504 3720
rect 140455 3689 140467 3692
rect 140409 3683 140467 3689
rect 140498 3680 140504 3692
rect 140556 3720 140562 3732
rect 141973 3723 142031 3729
rect 141973 3720 141985 3723
rect 140556 3692 141985 3720
rect 140556 3680 140562 3692
rect 141973 3689 141985 3692
rect 142019 3720 142031 3723
rect 142338 3720 142344 3732
rect 142019 3692 142344 3720
rect 142019 3689 142031 3692
rect 141973 3683 142031 3689
rect 142338 3680 142344 3692
rect 142396 3680 142402 3732
rect 142525 3723 142583 3729
rect 142525 3689 142537 3723
rect 142571 3720 142583 3723
rect 142614 3720 142620 3732
rect 142571 3692 142620 3720
rect 142571 3689 142583 3692
rect 142525 3683 142583 3689
rect 142614 3680 142620 3692
rect 142672 3680 142678 3732
rect 146294 3720 146300 3732
rect 142816 3692 145236 3720
rect 146255 3692 146300 3720
rect 142816 3652 142844 3692
rect 139872 3624 142844 3652
rect 144178 3584 144184 3596
rect 131439 3556 138888 3584
rect 144139 3556 144184 3584
rect 131439 3553 131451 3556
rect 131393 3547 131451 3553
rect 144178 3544 144184 3556
rect 144236 3544 144242 3596
rect 128648 3488 128952 3516
rect 129001 3519 129059 3525
rect 128648 3448 128676 3488
rect 129001 3485 129013 3519
rect 129047 3516 129059 3519
rect 129182 3516 129188 3528
rect 129047 3488 129188 3516
rect 129047 3485 129059 3488
rect 129001 3479 129059 3485
rect 129182 3476 129188 3488
rect 129240 3516 129246 3528
rect 130841 3519 130899 3525
rect 130841 3516 130853 3519
rect 129240 3488 130853 3516
rect 129240 3476 129246 3488
rect 130841 3485 130853 3488
rect 130887 3516 130899 3519
rect 131853 3519 131911 3525
rect 131408 3516 131528 3518
rect 131853 3516 131865 3519
rect 130887 3490 131865 3516
rect 130887 3488 131436 3490
rect 131500 3488 131865 3490
rect 130887 3485 130899 3488
rect 130841 3479 130899 3485
rect 131853 3485 131865 3488
rect 131899 3516 131911 3519
rect 132494 3516 132500 3528
rect 131899 3488 132500 3516
rect 131899 3485 131911 3488
rect 131853 3479 131911 3485
rect 132494 3476 132500 3488
rect 132552 3476 132558 3528
rect 132678 3476 132684 3528
rect 132736 3516 132742 3528
rect 132773 3519 132831 3525
rect 132773 3516 132785 3519
rect 132736 3488 132785 3516
rect 132736 3476 132742 3488
rect 132773 3485 132785 3488
rect 132819 3485 132831 3519
rect 132954 3516 132960 3528
rect 132915 3488 132960 3516
rect 132773 3479 132831 3485
rect 132954 3476 132960 3488
rect 133012 3476 133018 3528
rect 133141 3519 133199 3525
rect 133141 3485 133153 3519
rect 133187 3516 133199 3519
rect 133230 3516 133236 3528
rect 133187 3488 133236 3516
rect 133187 3485 133199 3488
rect 133141 3479 133199 3485
rect 133230 3476 133236 3488
rect 133288 3516 133294 3528
rect 133506 3516 133512 3528
rect 133288 3488 133512 3516
rect 133288 3476 133294 3488
rect 133506 3476 133512 3488
rect 133564 3516 133570 3528
rect 134153 3519 134211 3525
rect 134153 3516 134165 3519
rect 133564 3488 134165 3516
rect 133564 3476 133570 3488
rect 134153 3485 134165 3488
rect 134199 3485 134211 3519
rect 135346 3516 135352 3528
rect 135259 3488 135352 3516
rect 134153 3479 134211 3485
rect 135346 3476 135352 3488
rect 135404 3516 135410 3528
rect 135901 3519 135959 3525
rect 135901 3516 135913 3519
rect 135404 3488 135913 3516
rect 135404 3476 135410 3488
rect 135901 3485 135913 3488
rect 135947 3516 135959 3519
rect 137278 3516 137284 3528
rect 135947 3488 137284 3516
rect 135947 3485 135959 3488
rect 135901 3479 135959 3485
rect 137278 3476 137284 3488
rect 137336 3516 137342 3528
rect 137646 3516 137652 3528
rect 137336 3488 137652 3516
rect 137336 3476 137342 3488
rect 137646 3476 137652 3488
rect 137704 3516 137710 3528
rect 138017 3519 138075 3525
rect 138017 3516 138029 3519
rect 137704 3488 138029 3516
rect 137704 3476 137710 3488
rect 138017 3485 138029 3488
rect 138063 3516 138075 3519
rect 139857 3519 139915 3525
rect 139857 3516 139869 3519
rect 138063 3488 139869 3516
rect 138063 3485 138075 3488
rect 138017 3479 138075 3485
rect 139857 3485 139869 3488
rect 139903 3516 139915 3519
rect 139946 3516 139952 3528
rect 139903 3488 139952 3516
rect 139903 3485 139915 3488
rect 139857 3479 139915 3485
rect 139946 3476 139952 3488
rect 140004 3476 140010 3528
rect 143537 3519 143595 3525
rect 143537 3485 143549 3519
rect 143583 3516 143595 3519
rect 143626 3516 143632 3528
rect 143583 3488 143632 3516
rect 143583 3485 143595 3488
rect 143537 3479 143595 3485
rect 143626 3476 143632 3488
rect 143684 3476 143690 3528
rect 143718 3476 143724 3528
rect 143776 3516 143782 3528
rect 145208 3516 145236 3692
rect 146294 3680 146300 3692
rect 146352 3680 146358 3732
rect 149514 3720 149520 3732
rect 146404 3692 149520 3720
rect 145374 3612 145380 3664
rect 145432 3652 145438 3664
rect 146404 3652 146432 3692
rect 149514 3680 149520 3692
rect 149572 3680 149578 3732
rect 149606 3680 149612 3732
rect 149664 3720 149670 3732
rect 149885 3723 149943 3729
rect 149885 3720 149897 3723
rect 149664 3692 149897 3720
rect 149664 3680 149670 3692
rect 149885 3689 149897 3692
rect 149931 3689 149943 3723
rect 149885 3683 149943 3689
rect 150158 3680 150164 3732
rect 150216 3720 150222 3732
rect 152826 3720 152832 3732
rect 150216 3692 151860 3720
rect 152787 3692 152832 3720
rect 150216 3680 150222 3692
rect 148318 3652 148324 3664
rect 145432 3624 146432 3652
rect 147692 3624 148324 3652
rect 145432 3612 145438 3624
rect 147692 3584 147720 3624
rect 148318 3612 148324 3624
rect 148376 3612 148382 3664
rect 151832 3652 151860 3692
rect 152826 3680 152832 3692
rect 152884 3680 152890 3732
rect 156874 3720 156880 3732
rect 152936 3692 156880 3720
rect 152936 3652 152964 3692
rect 156874 3680 156880 3692
rect 156932 3680 156938 3732
rect 151832 3624 152964 3652
rect 155678 3612 155684 3664
rect 155736 3652 155742 3664
rect 156785 3655 156843 3661
rect 156785 3652 156797 3655
rect 155736 3624 156797 3652
rect 155736 3612 155742 3624
rect 156785 3621 156797 3624
rect 156831 3621 156843 3655
rect 156785 3615 156843 3621
rect 147600 3556 147720 3584
rect 147600 3516 147628 3556
rect 151814 3544 151820 3596
rect 151872 3584 151878 3596
rect 152550 3584 152556 3596
rect 151872 3556 152556 3584
rect 151872 3544 151878 3556
rect 152550 3544 152556 3556
rect 152608 3584 152614 3596
rect 152608 3556 152780 3584
rect 152608 3544 152614 3556
rect 143776 3488 144132 3516
rect 145208 3488 147628 3516
rect 143776 3476 143782 3488
rect 126808 3420 128676 3448
rect 128756 3451 128814 3457
rect 124438 3417 124450 3420
rect 124392 3411 124450 3417
rect 128756 3417 128768 3451
rect 128802 3448 128814 3451
rect 129090 3448 129096 3460
rect 128802 3420 129096 3448
rect 128802 3417 128814 3420
rect 128756 3411 128814 3417
rect 129090 3408 129096 3420
rect 129148 3408 129154 3460
rect 129734 3408 129740 3460
rect 129792 3448 129798 3460
rect 130470 3448 130476 3460
rect 129792 3420 130476 3448
rect 129792 3408 129798 3420
rect 130470 3408 130476 3420
rect 130528 3408 130534 3460
rect 130596 3451 130654 3457
rect 130596 3417 130608 3451
rect 130642 3448 130654 3451
rect 131206 3448 131212 3460
rect 130642 3420 131212 3448
rect 130642 3417 130654 3420
rect 130596 3411 130654 3417
rect 131206 3408 131212 3420
rect 131264 3408 131270 3460
rect 132972 3448 133000 3476
rect 133601 3451 133659 3457
rect 133601 3448 133613 3451
rect 132972 3420 133613 3448
rect 133601 3417 133613 3420
rect 133647 3417 133659 3451
rect 138290 3448 138296 3460
rect 133601 3411 133659 3417
rect 133708 3420 138296 3448
rect 127618 3380 127624 3392
rect 123588 3352 127624 3380
rect 127618 3340 127624 3352
rect 127676 3340 127682 3392
rect 127710 3340 127716 3392
rect 127768 3380 127774 3392
rect 129458 3380 129464 3392
rect 127768 3352 129464 3380
rect 127768 3340 127774 3352
rect 129458 3340 129464 3352
rect 129516 3340 129522 3392
rect 129918 3340 129924 3392
rect 129976 3380 129982 3392
rect 133708 3380 133736 3420
rect 138290 3408 138296 3420
rect 138348 3408 138354 3460
rect 138750 3408 138756 3460
rect 138808 3448 138814 3460
rect 139486 3448 139492 3460
rect 138808 3420 139492 3448
rect 138808 3408 138814 3420
rect 139486 3408 139492 3420
rect 139544 3408 139550 3460
rect 139612 3451 139670 3457
rect 139612 3417 139624 3451
rect 139658 3448 139670 3451
rect 140682 3448 140688 3460
rect 139658 3420 140688 3448
rect 139658 3417 139670 3420
rect 139612 3411 139670 3417
rect 140682 3408 140688 3420
rect 140740 3408 140746 3460
rect 141050 3408 141056 3460
rect 141108 3448 141114 3460
rect 144104 3448 144132 3488
rect 147674 3476 147680 3528
rect 147732 3516 147738 3528
rect 148042 3516 148048 3528
rect 147732 3488 148048 3516
rect 147732 3476 147738 3488
rect 148042 3476 148048 3488
rect 148100 3476 148106 3528
rect 148505 3519 148563 3525
rect 148505 3485 148517 3519
rect 148551 3516 148563 3519
rect 148551 3488 149008 3516
rect 148551 3485 148563 3488
rect 148505 3479 148563 3485
rect 144426 3451 144484 3457
rect 144426 3448 144438 3451
rect 141108 3420 143856 3448
rect 144104 3420 144438 3448
rect 141108 3408 141114 3420
rect 134702 3380 134708 3392
rect 129976 3352 133736 3380
rect 134663 3352 134708 3380
rect 129976 3340 129982 3352
rect 134702 3340 134708 3352
rect 134760 3380 134766 3392
rect 135346 3380 135352 3392
rect 134760 3352 135352 3380
rect 134760 3340 134766 3352
rect 135346 3340 135352 3352
rect 135404 3340 135410 3392
rect 136450 3380 136456 3392
rect 136411 3352 136456 3380
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 136910 3380 136916 3392
rect 136871 3352 136916 3380
rect 136910 3340 136916 3352
rect 136968 3340 136974 3392
rect 137186 3340 137192 3392
rect 137244 3380 137250 3392
rect 139854 3380 139860 3392
rect 137244 3352 139860 3380
rect 137244 3340 137250 3352
rect 139854 3340 139860 3352
rect 139912 3340 139918 3392
rect 140590 3340 140596 3392
rect 140648 3380 140654 3392
rect 140961 3383 141019 3389
rect 140961 3380 140973 3383
rect 140648 3352 140973 3380
rect 140648 3340 140654 3352
rect 140961 3349 140973 3352
rect 141007 3380 141019 3383
rect 142982 3380 142988 3392
rect 141007 3352 142988 3380
rect 141007 3349 141019 3352
rect 140961 3343 141019 3349
rect 142982 3340 142988 3352
rect 143040 3340 143046 3392
rect 143718 3380 143724 3392
rect 143679 3352 143724 3380
rect 143718 3340 143724 3352
rect 143776 3340 143782 3392
rect 143828 3380 143856 3420
rect 144426 3417 144438 3420
rect 144472 3417 144484 3451
rect 144426 3411 144484 3417
rect 145006 3408 145012 3460
rect 145064 3448 145070 3460
rect 147306 3448 147312 3460
rect 145064 3420 147312 3448
rect 145064 3408 145070 3420
rect 147306 3408 147312 3420
rect 147364 3408 147370 3460
rect 147432 3451 147490 3457
rect 147432 3417 147444 3451
rect 147478 3448 147490 3451
rect 147582 3448 147588 3460
rect 147478 3420 147588 3448
rect 147478 3417 147490 3420
rect 147432 3411 147490 3417
rect 147582 3408 147588 3420
rect 147640 3408 147646 3460
rect 148226 3408 148232 3460
rect 148284 3448 148290 3460
rect 148750 3451 148808 3457
rect 148750 3448 148762 3451
rect 148284 3420 148762 3448
rect 148284 3408 148290 3420
rect 148750 3417 148762 3420
rect 148796 3417 148808 3451
rect 148980 3448 149008 3488
rect 149054 3476 149060 3528
rect 149112 3516 149118 3528
rect 152458 3516 152464 3528
rect 149112 3488 151676 3516
rect 152419 3488 152464 3516
rect 149112 3476 149118 3488
rect 149882 3448 149888 3460
rect 148980 3420 149888 3448
rect 148750 3411 148808 3417
rect 149882 3408 149888 3420
rect 149940 3408 149946 3460
rect 149974 3408 149980 3460
rect 150032 3448 150038 3460
rect 150618 3448 150624 3460
rect 150032 3420 150624 3448
rect 150032 3408 150038 3420
rect 150618 3408 150624 3420
rect 150676 3408 150682 3460
rect 151538 3448 151544 3460
rect 151596 3457 151602 3460
rect 151508 3420 151544 3448
rect 151538 3408 151544 3420
rect 151596 3411 151608 3457
rect 151648 3448 151676 3488
rect 152458 3476 152464 3488
rect 152516 3476 152522 3528
rect 152645 3519 152703 3525
rect 152645 3485 152657 3519
rect 152691 3485 152703 3519
rect 152645 3479 152703 3485
rect 152660 3448 152688 3479
rect 151648 3420 152688 3448
rect 152752 3448 152780 3556
rect 153102 3476 153108 3528
rect 153160 3516 153166 3528
rect 154298 3516 154304 3528
rect 153160 3488 154304 3516
rect 153160 3476 153166 3488
rect 154298 3476 154304 3488
rect 154356 3476 154362 3528
rect 155126 3516 155132 3528
rect 155087 3488 155132 3516
rect 155126 3476 155132 3488
rect 155184 3476 155190 3528
rect 155770 3516 155776 3528
rect 155731 3488 155776 3516
rect 155770 3476 155776 3488
rect 155828 3476 155834 3528
rect 155865 3519 155923 3525
rect 155865 3485 155877 3519
rect 155911 3485 155923 3519
rect 156966 3516 156972 3528
rect 156927 3488 156972 3516
rect 155865 3479 155923 3485
rect 154666 3448 154672 3460
rect 152752 3420 154672 3448
rect 151596 3408 151602 3411
rect 154666 3408 154672 3420
rect 154724 3408 154730 3460
rect 154884 3451 154942 3457
rect 154884 3417 154896 3451
rect 154930 3448 154942 3451
rect 155034 3448 155040 3460
rect 154930 3420 155040 3448
rect 154930 3417 154942 3420
rect 154884 3411 154942 3417
rect 155034 3408 155040 3420
rect 155092 3408 155098 3460
rect 155218 3408 155224 3460
rect 155276 3448 155282 3460
rect 155880 3448 155908 3479
rect 156966 3476 156972 3488
rect 157024 3476 157030 3528
rect 157610 3516 157616 3528
rect 157571 3488 157616 3516
rect 157610 3476 157616 3488
rect 157668 3476 157674 3528
rect 155276 3420 155908 3448
rect 155276 3408 155282 3420
rect 145561 3383 145619 3389
rect 145561 3380 145573 3383
rect 143828 3352 145573 3380
rect 145561 3349 145573 3352
rect 145607 3380 145619 3383
rect 146202 3380 146208 3392
rect 145607 3352 146208 3380
rect 145607 3349 145619 3352
rect 145561 3343 145619 3349
rect 146202 3340 146208 3352
rect 146260 3340 146266 3392
rect 146570 3340 146576 3392
rect 146628 3380 146634 3392
rect 149146 3380 149152 3392
rect 146628 3352 149152 3380
rect 146628 3340 146634 3352
rect 149146 3340 149152 3352
rect 149204 3340 149210 3392
rect 149238 3340 149244 3392
rect 149296 3380 149302 3392
rect 150437 3383 150495 3389
rect 150437 3380 150449 3383
rect 149296 3352 150449 3380
rect 149296 3340 149302 3352
rect 150437 3349 150449 3352
rect 150483 3349 150495 3383
rect 150437 3343 150495 3349
rect 151262 3340 151268 3392
rect 151320 3380 151326 3392
rect 153378 3380 153384 3392
rect 151320 3352 153384 3380
rect 151320 3340 151326 3352
rect 153378 3340 153384 3352
rect 153436 3340 153442 3392
rect 153746 3380 153752 3392
rect 153707 3352 153752 3380
rect 153746 3340 153752 3352
rect 153804 3340 153810 3392
rect 153930 3340 153936 3392
rect 153988 3380 153994 3392
rect 155589 3383 155647 3389
rect 155589 3380 155601 3383
rect 153988 3352 155601 3380
rect 153988 3340 153994 3352
rect 155589 3349 155601 3352
rect 155635 3349 155647 3383
rect 157426 3380 157432 3392
rect 157387 3352 157432 3380
rect 155589 3343 155647 3349
rect 157426 3340 157432 3352
rect 157484 3340 157490 3392
rect 1104 3290 159043 3312
rect 1104 3238 40394 3290
rect 40446 3238 40458 3290
rect 40510 3238 40522 3290
rect 40574 3238 40586 3290
rect 40638 3238 40650 3290
rect 40702 3238 79839 3290
rect 79891 3238 79903 3290
rect 79955 3238 79967 3290
rect 80019 3238 80031 3290
rect 80083 3238 80095 3290
rect 80147 3238 119284 3290
rect 119336 3238 119348 3290
rect 119400 3238 119412 3290
rect 119464 3238 119476 3290
rect 119528 3238 119540 3290
rect 119592 3238 158729 3290
rect 158781 3238 158793 3290
rect 158845 3238 158857 3290
rect 158909 3238 158921 3290
rect 158973 3238 158985 3290
rect 159037 3238 159043 3290
rect 1104 3216 159043 3238
rect 11054 3176 11060 3188
rect 11015 3148 11060 3176
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11701 3179 11759 3185
rect 11701 3176 11713 3179
rect 11480 3148 11713 3176
rect 11480 3136 11486 3148
rect 11701 3145 11713 3148
rect 11747 3145 11759 3179
rect 11701 3139 11759 3145
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 13906 3176 13912 3188
rect 13771 3148 13912 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 13998 3136 14004 3188
rect 14056 3176 14062 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 14056 3148 14197 3176
rect 14056 3136 14062 3148
rect 14185 3145 14197 3148
rect 14231 3145 14243 3179
rect 14185 3139 14243 3145
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 18782 3176 18788 3188
rect 17083 3148 18788 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 20070 3176 20076 3188
rect 20031 3148 20076 3176
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 23934 3176 23940 3188
rect 22388 3148 22968 3176
rect 23895 3148 23940 3176
rect 12836 3111 12894 3117
rect 12836 3077 12848 3111
rect 12882 3108 12894 3111
rect 13354 3108 13360 3120
rect 12882 3080 13360 3108
rect 12882 3077 12894 3080
rect 12836 3071 12894 3077
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15381 3111 15439 3117
rect 15381 3108 15393 3111
rect 15160 3080 15393 3108
rect 15160 3068 15166 3080
rect 15381 3077 15393 3080
rect 15427 3108 15439 3111
rect 15427 3080 18276 3108
rect 15427 3077 15439 3080
rect 15381 3071 15439 3077
rect 18248 3052 18276 3080
rect 18322 3068 18328 3120
rect 18380 3108 18386 3120
rect 18478 3111 18536 3117
rect 18478 3108 18490 3111
rect 18380 3080 18490 3108
rect 18380 3068 18386 3080
rect 18478 3077 18490 3080
rect 18524 3077 18536 3111
rect 18478 3071 18536 3077
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 20530 3108 20536 3120
rect 18656 3080 20536 3108
rect 18656 3068 18662 3080
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 22388 3108 22416 3148
rect 20649 3080 22416 3108
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 18230 3040 18236 3052
rect 18191 3012 18236 3040
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 19334 3040 19340 3052
rect 18340 3012 19340 3040
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13814 2972 13820 2984
rect 13127 2944 13820 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14516 2944 14841 2972
rect 14516 2932 14522 2944
rect 14829 2941 14841 2944
rect 14875 2972 14887 2975
rect 18340 2972 18368 3012
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 20649 2972 20677 3080
rect 22462 3068 22468 3120
rect 22520 3108 22526 3120
rect 22802 3111 22860 3117
rect 22802 3108 22814 3111
rect 22520 3080 22814 3108
rect 22520 3068 22526 3080
rect 22802 3077 22814 3080
rect 22848 3077 22860 3111
rect 22940 3108 22968 3148
rect 23934 3136 23940 3148
rect 23992 3136 23998 3188
rect 24394 3136 24400 3188
rect 24452 3176 24458 3188
rect 24489 3179 24547 3185
rect 24489 3176 24501 3179
rect 24452 3148 24501 3176
rect 24452 3136 24458 3148
rect 24489 3145 24501 3148
rect 24535 3176 24547 3179
rect 24670 3176 24676 3188
rect 24535 3148 24676 3176
rect 24535 3145 24547 3148
rect 24489 3139 24547 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 31665 3179 31723 3185
rect 31665 3176 31677 3179
rect 24820 3148 31677 3176
rect 24820 3136 24826 3148
rect 31665 3145 31677 3148
rect 31711 3145 31723 3179
rect 31665 3139 31723 3145
rect 32677 3179 32735 3185
rect 32677 3145 32689 3179
rect 32723 3176 32735 3179
rect 32766 3176 32772 3188
rect 32723 3148 32772 3176
rect 32723 3145 32735 3148
rect 32677 3139 32735 3145
rect 32766 3136 32772 3148
rect 32824 3136 32830 3188
rect 32950 3136 32956 3188
rect 33008 3176 33014 3188
rect 44453 3179 44511 3185
rect 44453 3176 44465 3179
rect 33008 3148 44465 3176
rect 33008 3136 33014 3148
rect 44453 3145 44465 3148
rect 44499 3145 44511 3179
rect 44453 3139 44511 3145
rect 49145 3179 49203 3185
rect 49145 3145 49157 3179
rect 49191 3176 49203 3179
rect 50798 3176 50804 3188
rect 49191 3148 50804 3176
rect 49191 3145 49203 3148
rect 49145 3139 49203 3145
rect 26786 3108 26792 3120
rect 22940 3080 26792 3108
rect 22802 3071 22860 3077
rect 26786 3068 26792 3080
rect 26844 3068 26850 3120
rect 26970 3068 26976 3120
rect 27028 3108 27034 3120
rect 37918 3108 37924 3120
rect 27028 3080 37924 3108
rect 27028 3068 27034 3080
rect 37918 3068 37924 3080
rect 37976 3068 37982 3120
rect 44468 3108 44496 3139
rect 50798 3136 50804 3148
rect 50856 3176 50862 3188
rect 62577 3179 62635 3185
rect 62577 3176 62589 3179
rect 50856 3148 62589 3176
rect 50856 3136 50862 3148
rect 62577 3145 62589 3148
rect 62623 3145 62635 3179
rect 66254 3176 66260 3188
rect 66215 3148 66260 3176
rect 62577 3139 62635 3145
rect 46118 3111 46176 3117
rect 46118 3108 46130 3111
rect 44468 3080 46130 3108
rect 46118 3077 46130 3080
rect 46164 3077 46176 3111
rect 47210 3108 47216 3120
rect 47123 3080 47216 3108
rect 46118 3071 46176 3077
rect 47210 3068 47216 3080
rect 47268 3108 47274 3120
rect 56410 3117 56416 3120
rect 55585 3111 55643 3117
rect 55585 3108 55597 3111
rect 47268 3080 55597 3108
rect 47268 3068 47274 3080
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 20806 3040 20812 3052
rect 20763 3012 20812 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 22554 3040 22560 3052
rect 22515 3012 22560 3040
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 30541 3043 30599 3049
rect 30541 3040 30553 3043
rect 29748 3012 30553 3040
rect 14875 2944 18368 2972
rect 19260 2944 20677 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 15252 2876 18092 2904
rect 15252 2864 15258 2876
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 17954 2836 17960 2848
rect 17635 2808 17960 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18064 2836 18092 2876
rect 19260 2836 19288 2944
rect 23934 2932 23940 2984
rect 23992 2972 23998 2984
rect 29748 2981 29776 3012
rect 30541 3009 30553 3012
rect 30587 3009 30599 3043
rect 30541 3003 30599 3009
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 32493 3043 32551 3049
rect 31076 3012 32352 3040
rect 31076 3000 31082 3012
rect 29733 2975 29791 2981
rect 29733 2972 29745 2975
rect 23992 2944 29745 2972
rect 23992 2932 23998 2944
rect 29733 2941 29745 2944
rect 29779 2941 29791 2975
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 29733 2935 29791 2941
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 32324 2981 32352 3012
rect 32493 3009 32505 3043
rect 32539 3040 32551 3043
rect 33042 3040 33048 3052
rect 32539 3012 33048 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 33042 3000 33048 3012
rect 33100 3040 33106 3052
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 33100 3012 33701 3040
rect 33100 3000 33106 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 41794 3043 41852 3049
rect 41794 3040 41806 3043
rect 33689 3003 33747 3009
rect 40144 3012 41806 3040
rect 32309 2975 32367 2981
rect 32309 2941 32321 2975
rect 32355 2972 32367 2975
rect 33137 2975 33195 2981
rect 33137 2972 33149 2975
rect 32355 2944 33149 2972
rect 32355 2941 32367 2944
rect 32309 2935 32367 2941
rect 33137 2941 33149 2944
rect 33183 2941 33195 2975
rect 33137 2935 33195 2941
rect 19613 2907 19671 2913
rect 19613 2873 19625 2907
rect 19659 2904 19671 2907
rect 20714 2904 20720 2916
rect 19659 2876 20720 2904
rect 19659 2873 19671 2876
rect 19613 2867 19671 2873
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 20901 2907 20959 2913
rect 20901 2873 20913 2907
rect 20947 2904 20959 2907
rect 22462 2904 22468 2916
rect 20947 2876 22468 2904
rect 20947 2873 20959 2876
rect 20901 2867 20959 2873
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 40144 2913 40172 3012
rect 41794 3009 41806 3012
rect 41840 3009 41852 3043
rect 41794 3003 41852 3009
rect 42061 3043 42119 3049
rect 42061 3009 42073 3043
rect 42107 3040 42119 3043
rect 44174 3040 44180 3052
rect 42107 3012 44180 3040
rect 42107 3009 42119 3012
rect 42061 3003 42119 3009
rect 44174 3000 44180 3012
rect 44232 3040 44238 3052
rect 46385 3043 46443 3049
rect 46385 3040 46397 3043
rect 44232 3012 46397 3040
rect 44232 3000 44238 3012
rect 46385 3009 46397 3012
rect 46431 3040 46443 3043
rect 46566 3040 46572 3052
rect 46431 3012 46572 3040
rect 46431 3009 46443 3012
rect 46385 3003 46443 3009
rect 46566 3000 46572 3012
rect 46624 3000 46630 3052
rect 47780 3049 47808 3080
rect 55585 3077 55597 3080
rect 55631 3108 55643 3111
rect 56404 3108 56416 3117
rect 55631 3080 56180 3108
rect 56371 3080 56416 3108
rect 55631 3077 55643 3080
rect 55585 3071 55643 3077
rect 48038 3049 48044 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3009 47823 3043
rect 48032 3040 48044 3049
rect 47999 3012 48044 3040
rect 47765 3003 47823 3009
rect 48032 3003 48044 3012
rect 48038 3000 48044 3003
rect 48096 3000 48102 3052
rect 49786 3000 49792 3052
rect 49844 3040 49850 3052
rect 50718 3043 50776 3049
rect 50718 3040 50730 3043
rect 49844 3012 50730 3040
rect 49844 3000 49850 3012
rect 50718 3009 50730 3012
rect 50764 3009 50776 3043
rect 50718 3003 50776 3009
rect 50985 3043 51043 3049
rect 50985 3009 50997 3043
rect 51031 3040 51043 3043
rect 51074 3040 51080 3052
rect 51031 3012 51080 3040
rect 51031 3009 51043 3012
rect 50985 3003 51043 3009
rect 51074 3000 51080 3012
rect 51132 3000 51138 3052
rect 56152 3049 56180 3080
rect 56404 3071 56416 3080
rect 56410 3068 56416 3071
rect 56468 3068 56474 3120
rect 62592 3108 62620 3139
rect 66254 3136 66260 3148
rect 66312 3136 66318 3188
rect 68465 3179 68523 3185
rect 68465 3145 68477 3179
rect 68511 3176 68523 3179
rect 69106 3176 69112 3188
rect 68511 3148 69112 3176
rect 68511 3145 68523 3148
rect 68465 3139 68523 3145
rect 69106 3136 69112 3148
rect 69164 3136 69170 3188
rect 69198 3136 69204 3188
rect 69256 3176 69262 3188
rect 76098 3176 76104 3188
rect 69256 3148 76104 3176
rect 69256 3136 69262 3148
rect 76098 3136 76104 3148
rect 76156 3136 76162 3188
rect 81158 3136 81164 3188
rect 81216 3176 81222 3188
rect 81253 3179 81311 3185
rect 81253 3176 81265 3179
rect 81216 3148 81265 3176
rect 81216 3136 81222 3148
rect 81253 3145 81265 3148
rect 81299 3176 81311 3179
rect 81342 3176 81348 3188
rect 81299 3148 81348 3176
rect 81299 3145 81311 3148
rect 81253 3139 81311 3145
rect 81342 3136 81348 3148
rect 81400 3136 81406 3188
rect 83090 3136 83096 3188
rect 83148 3176 83154 3188
rect 96246 3176 96252 3188
rect 83148 3148 94544 3176
rect 96207 3148 96252 3176
rect 83148 3136 83154 3148
rect 64334 3111 64392 3117
rect 64334 3108 64346 3111
rect 62592 3080 64346 3108
rect 64334 3077 64346 3080
rect 64380 3077 64392 3111
rect 94516 3108 94544 3148
rect 96246 3136 96252 3148
rect 96304 3136 96310 3188
rect 109310 3136 109316 3188
rect 109368 3176 109374 3188
rect 109589 3179 109647 3185
rect 109589 3176 109601 3179
rect 109368 3148 109601 3176
rect 109368 3136 109374 3148
rect 109589 3145 109601 3148
rect 109635 3145 109647 3179
rect 110138 3176 110144 3188
rect 110099 3148 110144 3176
rect 109589 3139 109647 3145
rect 110138 3136 110144 3148
rect 110196 3136 110202 3188
rect 114830 3176 114836 3188
rect 114791 3148 114836 3176
rect 114830 3136 114836 3148
rect 114888 3136 114894 3188
rect 115658 3176 115664 3188
rect 115619 3148 115664 3176
rect 115658 3136 115664 3148
rect 115716 3136 115722 3188
rect 116946 3176 116952 3188
rect 116859 3148 116952 3176
rect 116946 3136 116952 3148
rect 117004 3176 117010 3188
rect 117004 3148 119108 3176
rect 117004 3136 117010 3148
rect 108298 3108 108304 3120
rect 64334 3071 64392 3077
rect 64432 3080 94452 3108
rect 94516 3080 108304 3108
rect 56137 3043 56195 3049
rect 56137 3009 56149 3043
rect 56183 3009 56195 3043
rect 56137 3003 56195 3009
rect 62022 3000 62028 3052
rect 62080 3040 62086 3052
rect 64432 3040 64460 3080
rect 64598 3040 64604 3052
rect 62080 3012 64460 3040
rect 64559 3012 64604 3040
rect 62080 3000 62086 3012
rect 64598 3000 64604 3012
rect 64656 3000 64662 3052
rect 67370 3043 67428 3049
rect 67370 3040 67382 3043
rect 65720 3012 67382 3040
rect 42886 2932 42892 2984
rect 42944 2972 42950 2984
rect 42944 2944 45416 2972
rect 42944 2932 42950 2944
rect 40129 2907 40187 2913
rect 40129 2904 40141 2907
rect 23860 2876 29868 2904
rect 18064 2808 19288 2836
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 23860 2836 23888 2876
rect 19392 2808 23888 2836
rect 29840 2836 29868 2876
rect 31220 2876 40141 2904
rect 31220 2836 31248 2876
rect 40129 2873 40141 2876
rect 40175 2873 40187 2907
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 40129 2867 40187 2873
rect 40236 2876 40816 2904
rect 29840 2808 31248 2836
rect 19392 2796 19398 2808
rect 38838 2796 38844 2848
rect 38896 2836 38902 2848
rect 40236 2836 40264 2876
rect 38896 2808 40264 2836
rect 38896 2796 38902 2808
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 40681 2839 40739 2845
rect 40681 2836 40693 2839
rect 40368 2808 40693 2836
rect 40368 2796 40374 2808
rect 40681 2805 40693 2808
rect 40727 2805 40739 2839
rect 40788 2836 40816 2876
rect 43180 2876 45017 2904
rect 43180 2836 43208 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45005 2867 45063 2873
rect 40788 2808 43208 2836
rect 45388 2836 45416 2944
rect 49694 2864 49700 2916
rect 49752 2864 49758 2916
rect 57238 2864 57244 2916
rect 57296 2904 57302 2916
rect 63221 2907 63279 2913
rect 63221 2904 63233 2907
rect 57296 2876 63233 2904
rect 57296 2864 57302 2876
rect 63221 2873 63233 2876
rect 63267 2873 63279 2907
rect 63221 2867 63279 2873
rect 49605 2839 49663 2845
rect 49605 2836 49617 2839
rect 45388 2808 49617 2836
rect 40681 2799 40739 2805
rect 49605 2805 49617 2808
rect 49651 2805 49663 2839
rect 49712 2836 49740 2864
rect 51718 2836 51724 2848
rect 49712 2808 51724 2836
rect 49605 2799 49663 2805
rect 51718 2796 51724 2808
rect 51776 2836 51782 2848
rect 57517 2839 57575 2845
rect 57517 2836 57529 2839
rect 51776 2808 57529 2836
rect 51776 2796 51782 2808
rect 57517 2805 57529 2808
rect 57563 2805 57575 2839
rect 57517 2799 57575 2805
rect 57606 2796 57612 2848
rect 57664 2836 57670 2848
rect 65720 2845 65748 3012
rect 67370 3009 67382 3012
rect 67416 3009 67428 3043
rect 67370 3003 67428 3009
rect 67542 3000 67548 3052
rect 67600 3040 67606 3052
rect 94424 3040 94452 3080
rect 108298 3068 108304 3080
rect 108356 3068 108362 3120
rect 108390 3068 108396 3120
rect 108448 3108 108454 3120
rect 118510 3108 118516 3120
rect 108448 3080 118516 3108
rect 108448 3068 108454 3080
rect 118510 3068 118516 3080
rect 118568 3068 118574 3120
rect 119080 3108 119108 3148
rect 119154 3136 119160 3188
rect 119212 3176 119218 3188
rect 126606 3176 126612 3188
rect 119212 3148 126612 3176
rect 119212 3136 119218 3148
rect 126606 3136 126612 3148
rect 126664 3136 126670 3188
rect 126790 3176 126796 3188
rect 126751 3148 126796 3176
rect 126790 3136 126796 3148
rect 126848 3136 126854 3188
rect 127066 3136 127072 3188
rect 127124 3176 127130 3188
rect 127894 3176 127900 3188
rect 127124 3148 127900 3176
rect 127124 3136 127130 3148
rect 127894 3136 127900 3148
rect 127952 3136 127958 3188
rect 129090 3176 129096 3188
rect 129051 3148 129096 3176
rect 129090 3136 129096 3148
rect 129148 3136 129154 3188
rect 131117 3179 131175 3185
rect 131117 3145 131129 3179
rect 131163 3176 131175 3179
rect 131942 3176 131948 3188
rect 131163 3148 131948 3176
rect 131163 3145 131175 3148
rect 131117 3139 131175 3145
rect 131942 3136 131948 3148
rect 132000 3136 132006 3188
rect 132494 3136 132500 3188
rect 132552 3176 132558 3188
rect 132865 3179 132923 3185
rect 132865 3176 132877 3179
rect 132552 3148 132877 3176
rect 132552 3136 132558 3148
rect 132865 3145 132877 3148
rect 132911 3176 132923 3179
rect 134153 3179 134211 3185
rect 134153 3176 134165 3179
rect 132911 3148 134165 3176
rect 132911 3145 132923 3148
rect 132865 3139 132923 3145
rect 134153 3145 134165 3148
rect 134199 3176 134211 3179
rect 134702 3176 134708 3188
rect 134199 3148 134708 3176
rect 134199 3145 134211 3148
rect 134153 3139 134211 3145
rect 134702 3136 134708 3148
rect 134760 3136 134766 3188
rect 135438 3176 135444 3188
rect 135399 3148 135444 3176
rect 135438 3136 135444 3148
rect 135496 3136 135502 3188
rect 136358 3176 136364 3188
rect 135548 3148 136364 3176
rect 121086 3108 121092 3120
rect 119080 3080 121092 3108
rect 121086 3068 121092 3080
rect 121144 3068 121150 3120
rect 122006 3068 122012 3120
rect 122064 3108 122070 3120
rect 125962 3108 125968 3120
rect 122064 3080 125968 3108
rect 122064 3068 122070 3080
rect 125962 3068 125968 3080
rect 126020 3068 126026 3120
rect 126328 3080 131436 3108
rect 96982 3040 96988 3052
rect 67600 3012 80054 3040
rect 94424 3012 96988 3040
rect 67600 3000 67606 3012
rect 67637 2975 67695 2981
rect 67637 2941 67649 2975
rect 67683 2972 67695 2975
rect 69106 2972 69112 2984
rect 67683 2944 69112 2972
rect 67683 2941 67695 2944
rect 67637 2935 67695 2941
rect 69106 2932 69112 2944
rect 69164 2972 69170 2984
rect 72789 2975 72847 2981
rect 72789 2972 72801 2975
rect 69164 2944 72801 2972
rect 69164 2932 69170 2944
rect 72789 2941 72801 2944
rect 72835 2972 72847 2975
rect 74534 2972 74540 2984
rect 72835 2944 74540 2972
rect 72835 2941 72847 2944
rect 72789 2935 72847 2941
rect 74534 2932 74540 2944
rect 74592 2932 74598 2984
rect 80026 2904 80054 3012
rect 96982 3000 96988 3012
rect 97040 3000 97046 3052
rect 107654 3000 107660 3052
rect 107712 3040 107718 3052
rect 114005 3043 114063 3049
rect 114005 3040 114017 3043
rect 107712 3012 114017 3040
rect 107712 3000 107718 3012
rect 114005 3009 114017 3012
rect 114051 3009 114063 3043
rect 114830 3040 114836 3052
rect 114005 3003 114063 3009
rect 114112 3012 114836 3040
rect 88518 2932 88524 2984
rect 88576 2972 88582 2984
rect 88576 2944 104204 2972
rect 88576 2932 88582 2944
rect 100846 2904 100852 2916
rect 80026 2876 100852 2904
rect 100846 2864 100852 2876
rect 100904 2864 100910 2916
rect 104176 2904 104204 2944
rect 106458 2932 106464 2984
rect 106516 2972 106522 2984
rect 113821 2975 113879 2981
rect 106516 2944 110184 2972
rect 106516 2932 106522 2944
rect 110046 2904 110052 2916
rect 104176 2876 110052 2904
rect 110046 2864 110052 2876
rect 110104 2864 110110 2916
rect 65705 2839 65763 2845
rect 65705 2836 65717 2839
rect 57664 2808 65717 2836
rect 57664 2796 57670 2808
rect 65705 2805 65717 2808
rect 65751 2805 65763 2839
rect 82998 2836 83004 2848
rect 82911 2808 83004 2836
rect 65705 2799 65763 2805
rect 82998 2796 83004 2808
rect 83056 2836 83062 2848
rect 98638 2836 98644 2848
rect 83056 2808 98644 2836
rect 83056 2796 83062 2808
rect 98638 2796 98644 2808
rect 98696 2796 98702 2848
rect 110156 2836 110184 2944
rect 113821 2941 113833 2975
rect 113867 2972 113879 2975
rect 114112 2972 114140 3012
rect 114830 3000 114836 3012
rect 114888 3000 114894 3052
rect 115474 3040 115480 3052
rect 115435 3012 115480 3040
rect 115474 3000 115480 3012
rect 115532 3000 115538 3052
rect 118237 3043 118295 3049
rect 118237 3009 118249 3043
rect 118283 3040 118295 3043
rect 118418 3040 118424 3052
rect 118283 3012 118424 3040
rect 118283 3009 118295 3012
rect 118237 3003 118295 3009
rect 118418 3000 118424 3012
rect 118476 3000 118482 3052
rect 126149 3043 126207 3049
rect 126149 3040 126161 3043
rect 118712 3012 126161 3040
rect 113867 2944 114140 2972
rect 114189 2975 114247 2981
rect 113867 2941 113879 2944
rect 113821 2935 113879 2941
rect 114189 2941 114201 2975
rect 114235 2972 114247 2975
rect 118712 2972 118740 3012
rect 126149 3009 126161 3012
rect 126195 3009 126207 3043
rect 126149 3003 126207 3009
rect 120074 2972 120080 2984
rect 114235 2944 118740 2972
rect 120035 2944 120080 2972
rect 114235 2941 114247 2944
rect 114189 2935 114247 2941
rect 120074 2932 120080 2944
rect 120132 2932 120138 2984
rect 120626 2972 120632 2984
rect 120587 2944 120632 2972
rect 120626 2932 120632 2944
rect 120684 2932 120690 2984
rect 120902 2932 120908 2984
rect 120960 2972 120966 2984
rect 121641 2975 121699 2981
rect 121641 2972 121653 2975
rect 120960 2944 121653 2972
rect 120960 2932 120966 2944
rect 121641 2941 121653 2944
rect 121687 2972 121699 2975
rect 122190 2972 122196 2984
rect 121687 2944 122196 2972
rect 121687 2941 121699 2944
rect 121641 2935 121699 2941
rect 122190 2932 122196 2944
rect 122248 2932 122254 2984
rect 122837 2975 122895 2981
rect 122837 2941 122849 2975
rect 122883 2972 122895 2975
rect 125594 2972 125600 2984
rect 122883 2944 125600 2972
rect 122883 2941 122895 2944
rect 122837 2935 122895 2941
rect 125594 2932 125600 2944
rect 125652 2932 125658 2984
rect 125962 2932 125968 2984
rect 126020 2972 126026 2984
rect 126328 2972 126356 3080
rect 131408 3064 131436 3080
rect 131574 3068 131580 3120
rect 131632 3108 131638 3120
rect 131632 3080 131677 3108
rect 131632 3068 131638 3080
rect 131850 3068 131856 3120
rect 131908 3108 131914 3120
rect 135548 3108 135576 3148
rect 136358 3136 136364 3148
rect 136416 3136 136422 3188
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 138661 3179 138719 3185
rect 136508 3148 138014 3176
rect 136508 3136 136514 3148
rect 137554 3117 137560 3120
rect 137548 3108 137560 3117
rect 131908 3080 135576 3108
rect 137515 3080 137560 3108
rect 131908 3068 131914 3080
rect 137548 3071 137560 3080
rect 137554 3068 137560 3071
rect 137612 3068 137618 3120
rect 137986 3108 138014 3148
rect 138661 3145 138673 3179
rect 138707 3176 138719 3179
rect 139670 3176 139676 3188
rect 138707 3148 139676 3176
rect 138707 3145 138719 3148
rect 138661 3139 138719 3145
rect 139670 3136 139676 3148
rect 139728 3136 139734 3188
rect 139854 3176 139860 3188
rect 139815 3148 139860 3176
rect 139854 3136 139860 3148
rect 139912 3136 139918 3188
rect 139946 3136 139952 3188
rect 140004 3176 140010 3188
rect 140593 3179 140651 3185
rect 140593 3176 140605 3179
rect 140004 3148 140605 3176
rect 140004 3136 140010 3148
rect 140593 3145 140605 3148
rect 140639 3176 140651 3179
rect 141418 3176 141424 3188
rect 140639 3148 141424 3176
rect 140639 3145 140651 3148
rect 140593 3139 140651 3145
rect 141418 3136 141424 3148
rect 141476 3176 141482 3188
rect 141970 3176 141976 3188
rect 141476 3148 141976 3176
rect 141476 3136 141482 3148
rect 141970 3136 141976 3148
rect 142028 3136 142034 3188
rect 142525 3179 142583 3185
rect 142525 3145 142537 3179
rect 142571 3176 142583 3179
rect 142614 3176 142620 3188
rect 142571 3148 142620 3176
rect 142571 3145 142583 3148
rect 142525 3139 142583 3145
rect 141694 3108 141700 3120
rect 137986 3080 141700 3108
rect 141694 3068 141700 3080
rect 141752 3068 141758 3120
rect 141881 3111 141939 3117
rect 141881 3077 141893 3111
rect 141927 3108 141939 3111
rect 142540 3108 142568 3139
rect 142614 3136 142620 3148
rect 142672 3136 142678 3188
rect 142890 3136 142896 3188
rect 142948 3176 142954 3188
rect 146478 3176 146484 3188
rect 142948 3148 146484 3176
rect 142948 3136 142954 3148
rect 146478 3136 146484 3148
rect 146536 3136 146542 3188
rect 147030 3176 147036 3188
rect 146991 3148 147036 3176
rect 147030 3136 147036 3148
rect 147088 3136 147094 3188
rect 147674 3176 147680 3188
rect 147508 3148 147680 3176
rect 141927 3080 142568 3108
rect 141927 3077 141939 3080
rect 141881 3071 141939 3077
rect 127437 3043 127495 3049
rect 127437 3009 127449 3043
rect 127483 3040 127495 3043
rect 127526 3040 127532 3052
rect 127483 3012 127532 3040
rect 127483 3009 127495 3012
rect 127437 3003 127495 3009
rect 127526 3000 127532 3012
rect 127584 3000 127590 3052
rect 128633 3043 128691 3049
rect 128633 3040 128645 3043
rect 127636 3012 128645 3040
rect 126020 2944 126356 2972
rect 126020 2932 126026 2944
rect 126606 2932 126612 2984
rect 126664 2972 126670 2984
rect 127636 2972 127664 3012
rect 128633 3009 128645 3012
rect 128679 3040 128691 3043
rect 129366 3040 129372 3052
rect 128679 3012 129372 3040
rect 128679 3009 128691 3012
rect 128633 3003 128691 3009
rect 129366 3000 129372 3012
rect 129424 3000 129430 3052
rect 130194 3000 130200 3052
rect 130252 3040 130258 3052
rect 130933 3043 130991 3049
rect 130933 3040 130945 3043
rect 130252 3012 130945 3040
rect 130252 3000 130258 3012
rect 130933 3009 130945 3012
rect 130979 3009 130991 3043
rect 131408 3040 131508 3064
rect 136554 3043 136612 3049
rect 136554 3040 136566 3043
rect 131408 3036 136566 3040
rect 131480 3012 136566 3036
rect 130933 3003 130991 3009
rect 136554 3009 136566 3012
rect 136600 3040 136612 3043
rect 136910 3040 136916 3052
rect 136600 3012 136916 3040
rect 136600 3009 136612 3012
rect 136554 3003 136612 3009
rect 136910 3000 136916 3012
rect 136968 3000 136974 3052
rect 137278 3040 137284 3052
rect 137239 3012 137284 3040
rect 137278 3000 137284 3012
rect 137336 3000 137342 3052
rect 139397 3043 139455 3049
rect 137388 3012 139348 3040
rect 126664 2944 127664 2972
rect 126664 2932 126670 2944
rect 127802 2932 127808 2984
rect 127860 2972 127866 2984
rect 130749 2975 130807 2981
rect 130749 2972 130761 2975
rect 127860 2944 130056 2972
rect 127860 2932 127866 2944
rect 110322 2864 110328 2916
rect 110380 2904 110386 2916
rect 118053 2907 118111 2913
rect 118053 2904 118065 2907
rect 110380 2876 118065 2904
rect 110380 2864 110386 2876
rect 118053 2873 118065 2876
rect 118099 2873 118111 2907
rect 118053 2867 118111 2873
rect 118789 2907 118847 2913
rect 118789 2873 118801 2907
rect 118835 2904 118847 2907
rect 129918 2904 129924 2916
rect 118835 2876 129924 2904
rect 118835 2873 118847 2876
rect 118789 2867 118847 2873
rect 129918 2864 129924 2876
rect 129976 2864 129982 2916
rect 111518 2836 111524 2848
rect 110156 2808 111524 2836
rect 111518 2796 111524 2808
rect 111576 2796 111582 2848
rect 117590 2836 117596 2848
rect 117551 2808 117596 2836
rect 117590 2796 117596 2808
rect 117648 2796 117654 2848
rect 117682 2796 117688 2848
rect 117740 2836 117746 2848
rect 119154 2836 119160 2848
rect 117740 2808 119160 2836
rect 117740 2796 117746 2808
rect 119154 2796 119160 2808
rect 119212 2796 119218 2848
rect 119338 2836 119344 2848
rect 119299 2808 119344 2836
rect 119338 2796 119344 2808
rect 119396 2796 119402 2848
rect 123386 2836 123392 2848
rect 123347 2808 123392 2836
rect 123386 2796 123392 2808
rect 123444 2796 123450 2848
rect 123846 2836 123852 2848
rect 123807 2808 123852 2836
rect 123846 2796 123852 2808
rect 123904 2796 123910 2848
rect 123938 2796 123944 2848
rect 123996 2836 124002 2848
rect 124401 2839 124459 2845
rect 124401 2836 124413 2839
rect 123996 2808 124413 2836
rect 123996 2796 124002 2808
rect 124401 2805 124413 2808
rect 124447 2805 124459 2839
rect 124401 2799 124459 2805
rect 125137 2839 125195 2845
rect 125137 2805 125149 2839
rect 125183 2836 125195 2839
rect 125226 2836 125232 2848
rect 125183 2808 125232 2836
rect 125183 2805 125195 2808
rect 125137 2799 125195 2805
rect 125226 2796 125232 2808
rect 125284 2796 125290 2848
rect 125870 2796 125876 2848
rect 125928 2836 125934 2848
rect 125965 2839 126023 2845
rect 125965 2836 125977 2839
rect 125928 2808 125977 2836
rect 125928 2796 125934 2808
rect 125965 2805 125977 2808
rect 126011 2805 126023 2839
rect 125965 2799 126023 2805
rect 126054 2796 126060 2848
rect 126112 2836 126118 2848
rect 127253 2839 127311 2845
rect 127253 2836 127265 2839
rect 126112 2808 127265 2836
rect 126112 2796 126118 2808
rect 127253 2805 127265 2808
rect 127299 2805 127311 2839
rect 127253 2799 127311 2805
rect 127894 2796 127900 2848
rect 127952 2836 127958 2848
rect 128814 2836 128820 2848
rect 127952 2808 128820 2836
rect 127952 2796 127958 2808
rect 128814 2796 128820 2808
rect 128872 2796 128878 2848
rect 130028 2836 130056 2944
rect 130396 2944 130761 2972
rect 130194 2904 130200 2916
rect 130155 2876 130200 2904
rect 130194 2864 130200 2876
rect 130252 2864 130258 2916
rect 130396 2836 130424 2944
rect 130749 2941 130761 2944
rect 130795 2941 130807 2975
rect 130749 2935 130807 2941
rect 136821 2975 136879 2981
rect 136821 2941 136833 2975
rect 136867 2941 136879 2975
rect 136928 2972 136956 3000
rect 137388 2972 137416 3012
rect 136928 2944 137416 2972
rect 139320 2972 139348 3012
rect 139397 3009 139409 3043
rect 139443 3040 139455 3043
rect 142908 3040 142936 3136
rect 142982 3068 142988 3120
rect 143040 3108 143046 3120
rect 144764 3111 144822 3117
rect 143040 3080 144132 3108
rect 143040 3068 143046 3080
rect 139443 3012 142936 3040
rect 143169 3043 143227 3049
rect 139443 3009 139455 3012
rect 139397 3003 139455 3009
rect 143169 3009 143181 3043
rect 143215 3040 143227 3043
rect 144104 3040 144132 3080
rect 144764 3077 144776 3111
rect 144810 3108 144822 3111
rect 145466 3108 145472 3120
rect 144810 3080 145472 3108
rect 144810 3077 144822 3080
rect 144764 3071 144822 3077
rect 145466 3068 145472 3080
rect 145524 3068 145530 3120
rect 147508 3108 147536 3148
rect 147674 3136 147680 3148
rect 147732 3136 147738 3188
rect 150158 3176 150164 3188
rect 147784 3148 150164 3176
rect 145668 3080 147536 3108
rect 145558 3040 145564 3052
rect 143215 3012 144040 3040
rect 144104 3012 145564 3040
rect 143215 3009 143227 3012
rect 143169 3003 143227 3009
rect 143810 2972 143816 2984
rect 139320 2944 143816 2972
rect 136821 2935 136879 2941
rect 131114 2836 131120 2848
rect 130028 2808 131120 2836
rect 131114 2796 131120 2808
rect 131172 2796 131178 2848
rect 133138 2796 133144 2848
rect 133196 2836 133202 2848
rect 136836 2836 136864 2935
rect 143810 2932 143816 2944
rect 143868 2932 143874 2984
rect 143629 2907 143687 2913
rect 143629 2904 143641 2907
rect 138584 2876 143641 2904
rect 133196 2808 136864 2836
rect 133196 2796 133202 2808
rect 136910 2796 136916 2848
rect 136968 2836 136974 2848
rect 138584 2836 138612 2876
rect 143629 2873 143641 2876
rect 143675 2873 143687 2907
rect 143629 2867 143687 2873
rect 136968 2808 138612 2836
rect 136968 2796 136974 2808
rect 140682 2796 140688 2848
rect 140740 2836 140746 2848
rect 142985 2839 143043 2845
rect 142985 2836 142997 2839
rect 140740 2808 142997 2836
rect 140740 2796 140746 2808
rect 142985 2805 142997 2808
rect 143031 2805 143043 2839
rect 144012 2836 144040 3012
rect 145558 3000 145564 3012
rect 145616 3000 145622 3052
rect 145668 2984 145696 3080
rect 147508 3049 147536 3080
rect 147582 3068 147588 3120
rect 147640 3108 147646 3120
rect 147784 3108 147812 3148
rect 150158 3136 150164 3148
rect 150216 3136 150222 3188
rect 150710 3136 150716 3188
rect 150768 3176 150774 3188
rect 150805 3179 150863 3185
rect 150805 3176 150817 3179
rect 150768 3148 150817 3176
rect 150768 3136 150774 3148
rect 150805 3145 150817 3148
rect 150851 3145 150863 3179
rect 150805 3139 150863 3145
rect 150912 3148 154252 3176
rect 147640 3080 147812 3108
rect 147640 3068 147646 3080
rect 147858 3068 147864 3120
rect 147916 3108 147922 3120
rect 150912 3108 150940 3148
rect 151446 3108 151452 3120
rect 147916 3080 150940 3108
rect 151096 3080 151452 3108
rect 147916 3068 147922 3080
rect 145920 3043 145978 3049
rect 145920 3009 145932 3043
rect 145966 3040 145978 3043
rect 147493 3043 147551 3049
rect 145966 3012 147444 3040
rect 145966 3009 145978 3012
rect 145920 3003 145978 3009
rect 145009 2975 145067 2981
rect 145009 2941 145021 2975
rect 145055 2972 145067 2975
rect 145282 2972 145288 2984
rect 145055 2944 145288 2972
rect 145055 2941 145067 2944
rect 145009 2935 145067 2941
rect 145282 2932 145288 2944
rect 145340 2932 145346 2984
rect 145650 2972 145656 2984
rect 145611 2944 145656 2972
rect 145650 2932 145656 2944
rect 145708 2932 145714 2984
rect 146938 2836 146944 2848
rect 144012 2808 146944 2836
rect 142985 2799 143043 2805
rect 146938 2796 146944 2808
rect 146996 2796 147002 2848
rect 147416 2836 147444 3012
rect 147493 3009 147505 3043
rect 147539 3009 147551 3043
rect 147493 3003 147551 3009
rect 147760 3043 147818 3049
rect 147760 3009 147772 3043
rect 147806 3040 147818 3043
rect 149422 3040 149428 3052
rect 147806 3012 149428 3040
rect 147806 3009 147818 3012
rect 147760 3003 147818 3009
rect 149422 3000 149428 3012
rect 149480 3000 149486 3052
rect 149514 3000 149520 3052
rect 149572 3040 149578 3052
rect 149701 3043 149759 3049
rect 149572 3012 149617 3040
rect 149572 3000 149578 3012
rect 149701 3009 149713 3043
rect 149747 3040 149759 3043
rect 150526 3040 150532 3052
rect 149747 3012 150532 3040
rect 149747 3009 149759 3012
rect 149701 3003 149759 3009
rect 150526 3000 150532 3012
rect 150584 3000 150590 3052
rect 150618 3000 150624 3052
rect 150676 3040 150682 3052
rect 150989 3043 151047 3049
rect 150989 3040 151001 3043
rect 150676 3012 151001 3040
rect 150676 3000 150682 3012
rect 150989 3009 151001 3012
rect 151035 3009 151047 3043
rect 150989 3003 151047 3009
rect 149146 2932 149152 2984
rect 149204 2972 149210 2984
rect 149333 2975 149391 2981
rect 149333 2972 149345 2975
rect 149204 2944 149345 2972
rect 149204 2932 149210 2944
rect 149333 2941 149345 2944
rect 149379 2941 149391 2975
rect 149333 2935 149391 2941
rect 150253 2975 150311 2981
rect 150253 2941 150265 2975
rect 150299 2972 150311 2975
rect 151096 2972 151124 3080
rect 151446 3068 151452 3080
rect 151504 3068 151510 3120
rect 151998 3108 152004 3120
rect 151959 3080 152004 3108
rect 151998 3068 152004 3080
rect 152056 3068 152062 3120
rect 152185 3111 152243 3117
rect 152185 3077 152197 3111
rect 152231 3108 152243 3111
rect 152274 3108 152280 3120
rect 152231 3080 152280 3108
rect 152231 3077 152243 3080
rect 152185 3071 152243 3077
rect 152274 3068 152280 3080
rect 152332 3068 152338 3120
rect 151354 3000 151360 3052
rect 151412 3040 151418 3052
rect 153657 3043 153715 3049
rect 151412 3012 153148 3040
rect 151412 3000 151418 3012
rect 150299 2944 151124 2972
rect 151173 2975 151231 2981
rect 150299 2941 150311 2944
rect 150253 2935 150311 2941
rect 151173 2941 151185 2975
rect 151219 2972 151231 2975
rect 151814 2972 151820 2984
rect 151219 2944 151820 2972
rect 151219 2941 151231 2944
rect 151173 2935 151231 2941
rect 151814 2932 151820 2944
rect 151872 2932 151878 2984
rect 151906 2932 151912 2984
rect 151964 2972 151970 2984
rect 152737 2975 152795 2981
rect 152737 2972 152749 2975
rect 151964 2944 152749 2972
rect 151964 2932 151970 2944
rect 152737 2941 152749 2944
rect 152783 2972 152795 2975
rect 153010 2972 153016 2984
rect 152783 2944 153016 2972
rect 152783 2941 152795 2944
rect 152737 2935 152795 2941
rect 153010 2932 153016 2944
rect 153068 2932 153074 2984
rect 153120 2972 153148 3012
rect 153657 3009 153669 3043
rect 153703 3040 153715 3043
rect 153838 3040 153844 3052
rect 153703 3012 153844 3040
rect 153703 3009 153715 3012
rect 153657 3003 153715 3009
rect 153838 3000 153844 3012
rect 153896 3000 153902 3052
rect 154224 3044 154252 3148
rect 154390 3136 154396 3188
rect 154448 3136 154454 3188
rect 154574 3176 154580 3188
rect 154535 3148 154580 3176
rect 154574 3136 154580 3148
rect 154632 3136 154638 3188
rect 155405 3179 155463 3185
rect 155405 3145 155417 3179
rect 155451 3176 155463 3179
rect 156598 3176 156604 3188
rect 155451 3148 156604 3176
rect 155451 3145 155463 3148
rect 155405 3139 155463 3145
rect 156598 3136 156604 3148
rect 156656 3136 156662 3188
rect 157245 3179 157303 3185
rect 157245 3145 157257 3179
rect 157291 3176 157303 3179
rect 158162 3176 158168 3188
rect 157291 3148 158168 3176
rect 157291 3145 157303 3148
rect 157245 3139 157303 3145
rect 158162 3136 158168 3148
rect 158220 3136 158226 3188
rect 154408 3108 154436 3136
rect 154408 3080 156644 3108
rect 154393 3044 154451 3049
rect 154224 3043 154451 3044
rect 154224 3016 154405 3043
rect 154393 3009 154405 3016
rect 154439 3009 154451 3043
rect 154393 3003 154451 3009
rect 154482 3000 154488 3052
rect 154540 3040 154546 3052
rect 155126 3040 155132 3052
rect 154540 3012 155132 3040
rect 154540 3000 154546 3012
rect 155126 3000 155132 3012
rect 155184 3000 155190 3052
rect 155221 3043 155279 3049
rect 155221 3009 155233 3043
rect 155267 3040 155279 3043
rect 155402 3040 155408 3052
rect 155267 3012 155408 3040
rect 155267 3009 155279 3012
rect 155221 3003 155279 3009
rect 155402 3000 155408 3012
rect 155460 3000 155466 3052
rect 156616 3049 156644 3080
rect 156601 3043 156659 3049
rect 156601 3009 156613 3043
rect 156647 3009 156659 3043
rect 157058 3040 157064 3052
rect 157019 3012 157064 3040
rect 156601 3003 156659 3009
rect 157058 3000 157064 3012
rect 157116 3000 157122 3052
rect 158257 3043 158315 3049
rect 158257 3040 158269 3043
rect 157306 3012 158269 3040
rect 153120 2944 153884 2972
rect 148594 2864 148600 2916
rect 148652 2904 148658 2916
rect 148873 2907 148931 2913
rect 148652 2876 148824 2904
rect 148652 2864 148658 2876
rect 148686 2836 148692 2848
rect 147416 2808 148692 2836
rect 148686 2796 148692 2808
rect 148744 2796 148750 2848
rect 148796 2836 148824 2876
rect 148873 2873 148885 2907
rect 148919 2904 148931 2907
rect 151262 2904 151268 2916
rect 148919 2876 151268 2904
rect 148919 2873 148931 2876
rect 148873 2867 148931 2873
rect 151262 2864 151268 2876
rect 151320 2864 151326 2916
rect 153194 2904 153200 2916
rect 151832 2876 153200 2904
rect 151832 2836 151860 2876
rect 153194 2864 153200 2876
rect 153252 2864 153258 2916
rect 153470 2904 153476 2916
rect 153431 2876 153476 2904
rect 153470 2864 153476 2876
rect 153528 2864 153534 2916
rect 153856 2904 153884 2944
rect 154022 2932 154028 2984
rect 154080 2972 154086 2984
rect 154209 2975 154267 2981
rect 154209 2972 154221 2975
rect 154080 2944 154221 2972
rect 154080 2932 154086 2944
rect 154209 2941 154221 2944
rect 154255 2972 154267 2975
rect 154942 2972 154948 2984
rect 154255 2944 154948 2972
rect 154255 2941 154267 2944
rect 154209 2935 154267 2941
rect 154942 2932 154948 2944
rect 155000 2932 155006 2984
rect 155037 2975 155095 2981
rect 155037 2941 155049 2975
rect 155083 2972 155095 2975
rect 156230 2972 156236 2984
rect 155083 2944 156236 2972
rect 155083 2941 155095 2944
rect 155037 2935 155095 2941
rect 156230 2932 156236 2944
rect 156288 2932 156294 2984
rect 156322 2932 156328 2984
rect 156380 2972 156386 2984
rect 157306 2972 157334 3012
rect 158257 3009 158269 3012
rect 158303 3009 158315 3043
rect 158257 3003 158315 3009
rect 156380 2944 157334 2972
rect 156380 2932 156386 2944
rect 155586 2904 155592 2916
rect 153856 2876 155592 2904
rect 155586 2864 155592 2876
rect 155644 2864 155650 2916
rect 155954 2864 155960 2916
rect 156012 2904 156018 2916
rect 158073 2907 158131 2913
rect 158073 2904 158085 2907
rect 156012 2876 158085 2904
rect 156012 2864 156018 2876
rect 158073 2873 158085 2876
rect 158119 2873 158131 2907
rect 158073 2867 158131 2873
rect 148796 2808 151860 2836
rect 154206 2796 154212 2848
rect 154264 2836 154270 2848
rect 155770 2836 155776 2848
rect 154264 2808 155776 2836
rect 154264 2796 154270 2808
rect 155770 2796 155776 2808
rect 155828 2796 155834 2848
rect 156414 2836 156420 2848
rect 156375 2808 156420 2836
rect 156414 2796 156420 2808
rect 156472 2796 156478 2848
rect 156506 2796 156512 2848
rect 156564 2836 156570 2848
rect 157150 2836 157156 2848
rect 156564 2808 157156 2836
rect 156564 2796 156570 2808
rect 157150 2796 157156 2808
rect 157208 2796 157214 2848
rect 1104 2746 158884 2768
rect 1104 2694 20672 2746
rect 20724 2694 20736 2746
rect 20788 2694 20800 2746
rect 20852 2694 20864 2746
rect 20916 2694 20928 2746
rect 20980 2694 60117 2746
rect 60169 2694 60181 2746
rect 60233 2694 60245 2746
rect 60297 2694 60309 2746
rect 60361 2694 60373 2746
rect 60425 2694 99562 2746
rect 99614 2694 99626 2746
rect 99678 2694 99690 2746
rect 99742 2694 99754 2746
rect 99806 2694 99818 2746
rect 99870 2694 139007 2746
rect 139059 2694 139071 2746
rect 139123 2694 139135 2746
rect 139187 2694 139199 2746
rect 139251 2694 139263 2746
rect 139315 2694 158884 2746
rect 1104 2672 158884 2694
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 4764 2604 5273 2632
rect 4764 2592 4770 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 5261 2595 5319 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13814 2632 13820 2644
rect 13311 2604 13820 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 18012 2604 18245 2632
rect 18012 2592 18018 2604
rect 18233 2601 18245 2604
rect 18279 2632 18291 2635
rect 18782 2632 18788 2644
rect 18279 2604 18788 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 19610 2592 19616 2644
rect 19668 2632 19674 2644
rect 19797 2635 19855 2641
rect 19797 2632 19809 2635
rect 19668 2604 19809 2632
rect 19668 2592 19674 2604
rect 19797 2601 19809 2604
rect 19843 2601 19855 2635
rect 26421 2635 26479 2641
rect 26421 2632 26433 2635
rect 19797 2595 19855 2601
rect 24596 2604 26433 2632
rect 13630 2564 13636 2576
rect 6886 2536 13636 2564
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 5460 2468 6561 2496
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 5460 2437 5488 2468
rect 6549 2465 6561 2468
rect 6595 2496 6607 2499
rect 6886 2496 6914 2536
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 18877 2567 18935 2573
rect 18877 2533 18889 2567
rect 18923 2564 18935 2567
rect 19886 2564 19892 2576
rect 18923 2536 19892 2564
rect 18923 2533 18935 2536
rect 18877 2527 18935 2533
rect 19886 2524 19892 2536
rect 19944 2524 19950 2576
rect 11146 2496 11152 2508
rect 6595 2468 6914 2496
rect 9784 2468 11152 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5810 2428 5816 2440
rect 5675 2400 5816 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 5810 2388 5816 2400
rect 5868 2428 5874 2440
rect 9784 2428 9812 2468
rect 11146 2456 11152 2468
rect 11204 2496 11210 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11204 2468 12265 2496
rect 11204 2456 11210 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 12253 2459 12311 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 24596 2505 24624 2604
rect 26421 2601 26433 2604
rect 26467 2601 26479 2635
rect 26421 2595 26479 2601
rect 41322 2592 41328 2644
rect 41380 2632 41386 2644
rect 45373 2635 45431 2641
rect 45373 2632 45385 2635
rect 41380 2604 45385 2632
rect 41380 2592 41386 2604
rect 45373 2601 45385 2604
rect 45419 2601 45431 2635
rect 45373 2595 45431 2601
rect 49513 2635 49571 2641
rect 49513 2601 49525 2635
rect 49559 2632 49571 2635
rect 49694 2632 49700 2644
rect 49559 2604 49700 2632
rect 49559 2601 49571 2604
rect 49513 2595 49571 2601
rect 49694 2592 49700 2604
rect 49752 2592 49758 2644
rect 59814 2592 59820 2644
rect 59872 2632 59878 2644
rect 60093 2635 60151 2641
rect 60093 2632 60105 2635
rect 59872 2604 60105 2632
rect 59872 2592 59878 2604
rect 60093 2601 60105 2604
rect 60139 2601 60151 2635
rect 60093 2595 60151 2601
rect 60737 2635 60795 2641
rect 60737 2601 60749 2635
rect 60783 2632 60795 2635
rect 63310 2632 63316 2644
rect 60783 2604 63316 2632
rect 60783 2601 60795 2604
rect 60737 2595 60795 2601
rect 63310 2592 63316 2604
rect 63368 2632 63374 2644
rect 65797 2635 65855 2641
rect 65797 2632 65809 2635
rect 63368 2604 65809 2632
rect 63368 2592 63374 2604
rect 25958 2564 25964 2576
rect 25919 2536 25964 2564
rect 25958 2524 25964 2536
rect 26016 2524 26022 2576
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24452 2468 24593 2496
rect 24452 2456 24458 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 33778 2496 33784 2508
rect 33739 2468 33784 2496
rect 24581 2459 24639 2465
rect 33778 2456 33784 2468
rect 33836 2456 33842 2508
rect 46201 2499 46259 2505
rect 46201 2496 46213 2499
rect 45572 2468 46213 2496
rect 5868 2400 9812 2428
rect 5868 2388 5874 2400
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11112 2400 12081 2428
rect 11112 2388 11118 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 17460 2400 18705 2428
rect 17460 2388 17466 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 20921 2431 20979 2437
rect 20921 2397 20933 2431
rect 20967 2428 20979 2431
rect 21082 2428 21088 2440
rect 20967 2400 21088 2428
rect 20967 2397 20979 2400
rect 20921 2391 20979 2397
rect 21082 2388 21088 2400
rect 21140 2388 21146 2440
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 45572 2437 45600 2468
rect 46201 2465 46213 2468
rect 46247 2496 46259 2499
rect 47302 2496 47308 2508
rect 46247 2468 47308 2496
rect 46247 2465 46259 2468
rect 46201 2459 46259 2465
rect 47302 2456 47308 2468
rect 47360 2456 47366 2508
rect 58710 2496 58716 2508
rect 58671 2468 58716 2496
rect 58710 2456 58716 2468
rect 58768 2456 58774 2508
rect 63512 2505 63540 2604
rect 65797 2601 65809 2604
rect 65843 2601 65855 2635
rect 65797 2595 65855 2601
rect 71038 2592 71044 2644
rect 71096 2632 71102 2644
rect 74169 2635 74227 2641
rect 74169 2632 74181 2635
rect 71096 2604 74181 2632
rect 71096 2592 71102 2604
rect 74169 2601 74181 2604
rect 74215 2601 74227 2635
rect 81434 2632 81440 2644
rect 81395 2604 81440 2632
rect 74169 2595 74227 2601
rect 81434 2592 81440 2604
rect 81492 2592 81498 2644
rect 107286 2592 107292 2644
rect 107344 2632 107350 2644
rect 107565 2635 107623 2641
rect 107565 2632 107577 2635
rect 107344 2604 107577 2632
rect 107344 2592 107350 2604
rect 107565 2601 107577 2604
rect 107611 2601 107623 2635
rect 109586 2632 109592 2644
rect 109547 2604 109592 2632
rect 107565 2595 107623 2601
rect 109586 2592 109592 2604
rect 109644 2592 109650 2644
rect 112714 2592 112720 2644
rect 112772 2632 112778 2644
rect 113177 2635 113235 2641
rect 113177 2632 113189 2635
rect 112772 2604 113189 2632
rect 112772 2592 112778 2604
rect 113177 2601 113189 2604
rect 113223 2601 113235 2635
rect 113634 2632 113640 2644
rect 113595 2604 113640 2632
rect 113177 2595 113235 2601
rect 64877 2567 64935 2573
rect 64877 2533 64889 2567
rect 64923 2564 64935 2567
rect 65978 2564 65984 2576
rect 64923 2536 65984 2564
rect 64923 2533 64935 2536
rect 64877 2527 64935 2533
rect 65978 2524 65984 2536
rect 66036 2524 66042 2576
rect 63497 2499 63555 2505
rect 63497 2465 63509 2499
rect 63543 2465 63555 2499
rect 63497 2459 63555 2465
rect 108945 2499 109003 2505
rect 108945 2465 108957 2499
rect 108991 2496 109003 2499
rect 109604 2496 109632 2592
rect 108991 2468 109632 2496
rect 108991 2465 109003 2468
rect 108945 2459 109003 2465
rect 24837 2431 24895 2437
rect 24837 2428 24849 2431
rect 23624 2400 24849 2428
rect 23624 2388 23630 2400
rect 24837 2397 24849 2400
rect 24883 2397 24895 2431
rect 24837 2391 24895 2397
rect 45557 2431 45615 2437
rect 45557 2397 45569 2431
rect 45603 2397 45615 2431
rect 45557 2391 45615 2397
rect 45649 2431 45707 2437
rect 45649 2397 45661 2431
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2360 2283 2363
rect 11698 2360 11704 2372
rect 2271 2332 11704 2360
rect 2271 2329 2283 2332
rect 2225 2323 2283 2329
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 33514 2363 33572 2369
rect 33514 2360 33526 2363
rect 31772 2332 33526 2360
rect 31772 2304 31800 2332
rect 33514 2329 33526 2332
rect 33560 2329 33572 2363
rect 33514 2323 33572 2329
rect 44637 2363 44695 2369
rect 44637 2329 44649 2363
rect 44683 2360 44695 2363
rect 45370 2360 45376 2372
rect 44683 2332 45376 2360
rect 44683 2329 44695 2332
rect 44637 2323 44695 2329
rect 45370 2320 45376 2332
rect 45428 2360 45434 2372
rect 45664 2360 45692 2391
rect 56594 2388 56600 2440
rect 56652 2428 56658 2440
rect 58969 2431 59027 2437
rect 58969 2428 58981 2431
rect 56652 2400 58981 2428
rect 56652 2388 56658 2400
rect 58969 2397 58981 2400
rect 59015 2397 59027 2431
rect 58969 2391 59027 2397
rect 59262 2388 59268 2440
rect 59320 2428 59326 2440
rect 63753 2431 63811 2437
rect 63753 2428 63765 2431
rect 59320 2400 63765 2428
rect 59320 2388 59326 2400
rect 63753 2397 63765 2400
rect 63799 2397 63811 2431
rect 63753 2391 63811 2397
rect 73709 2431 73767 2437
rect 73709 2397 73721 2431
rect 73755 2428 73767 2431
rect 74534 2428 74540 2440
rect 73755 2400 74540 2428
rect 73755 2397 73767 2400
rect 73709 2391 73767 2397
rect 74534 2388 74540 2400
rect 74592 2428 74598 2440
rect 75549 2431 75607 2437
rect 75549 2428 75561 2431
rect 74592 2400 75561 2428
rect 74592 2388 74598 2400
rect 75549 2397 75561 2400
rect 75595 2397 75607 2431
rect 75549 2391 75607 2397
rect 81342 2388 81348 2440
rect 81400 2428 81406 2440
rect 82817 2431 82875 2437
rect 82817 2428 82829 2431
rect 81400 2400 82829 2428
rect 81400 2388 81406 2400
rect 82817 2397 82829 2400
rect 82863 2397 82875 2431
rect 82817 2391 82875 2397
rect 108689 2431 108747 2437
rect 108689 2397 108701 2431
rect 108735 2428 108747 2431
rect 111242 2428 111248 2440
rect 108735 2400 111248 2428
rect 108735 2397 108747 2400
rect 108689 2391 108747 2397
rect 111242 2388 111248 2400
rect 111300 2388 111306 2440
rect 113192 2428 113220 2595
rect 113634 2592 113640 2604
rect 113692 2592 113698 2644
rect 114462 2592 114468 2644
rect 114520 2632 114526 2644
rect 114741 2635 114799 2641
rect 114741 2632 114753 2635
rect 114520 2604 114753 2632
rect 114520 2592 114526 2604
rect 114741 2601 114753 2604
rect 114787 2601 114799 2635
rect 114741 2595 114799 2601
rect 122837 2635 122895 2641
rect 122837 2601 122849 2635
rect 122883 2632 122895 2635
rect 123294 2632 123300 2644
rect 122883 2604 123300 2632
rect 122883 2601 122895 2604
rect 122837 2595 122895 2601
rect 123294 2592 123300 2604
rect 123352 2592 123358 2644
rect 123389 2635 123447 2641
rect 123389 2601 123401 2635
rect 123435 2632 123447 2635
rect 125134 2632 125140 2644
rect 123435 2604 125140 2632
rect 123435 2601 123447 2604
rect 123389 2595 123447 2601
rect 125134 2592 125140 2604
rect 125192 2592 125198 2644
rect 125965 2635 126023 2641
rect 125965 2601 125977 2635
rect 126011 2632 126023 2635
rect 126330 2632 126336 2644
rect 126011 2604 126336 2632
rect 126011 2601 126023 2604
rect 125965 2595 126023 2601
rect 126330 2592 126336 2604
rect 126388 2592 126394 2644
rect 127066 2632 127072 2644
rect 127027 2604 127072 2632
rect 127066 2592 127072 2604
rect 127124 2592 127130 2644
rect 130194 2632 130200 2644
rect 130155 2604 130200 2632
rect 130194 2592 130200 2604
rect 130252 2592 130258 2644
rect 131574 2592 131580 2644
rect 131632 2632 131638 2644
rect 132129 2635 132187 2641
rect 132129 2632 132141 2635
rect 131632 2604 132141 2632
rect 131632 2592 131638 2604
rect 132129 2601 132141 2604
rect 132175 2601 132187 2635
rect 134610 2632 134616 2644
rect 132129 2595 132187 2601
rect 132466 2604 134472 2632
rect 134571 2604 134616 2632
rect 114005 2499 114063 2505
rect 114005 2465 114017 2499
rect 114051 2496 114063 2499
rect 114480 2496 114508 2592
rect 122190 2524 122196 2576
rect 122248 2564 122254 2576
rect 126422 2564 126428 2576
rect 122248 2536 126428 2564
rect 122248 2524 122254 2536
rect 126422 2524 126428 2536
rect 126480 2524 126486 2576
rect 132466 2564 132494 2604
rect 128326 2536 132494 2564
rect 134444 2564 134472 2604
rect 134610 2592 134616 2604
rect 134668 2592 134674 2644
rect 137278 2632 137284 2644
rect 134720 2604 137048 2632
rect 137239 2604 137284 2632
rect 134720 2564 134748 2604
rect 134444 2536 134748 2564
rect 137020 2564 137048 2604
rect 137278 2592 137284 2604
rect 137336 2592 137342 2644
rect 138658 2592 138664 2644
rect 138716 2632 138722 2644
rect 139489 2635 139547 2641
rect 139489 2632 139501 2635
rect 138716 2604 139501 2632
rect 138716 2592 138722 2604
rect 139489 2601 139501 2604
rect 139535 2632 139547 2635
rect 139762 2632 139768 2644
rect 139535 2604 139768 2632
rect 139535 2601 139547 2604
rect 139489 2595 139547 2601
rect 139762 2592 139768 2604
rect 139820 2592 139826 2644
rect 141602 2632 141608 2644
rect 139872 2604 141608 2632
rect 139872 2564 139900 2604
rect 141602 2592 141608 2604
rect 141660 2592 141666 2644
rect 142522 2632 142528 2644
rect 142483 2604 142528 2632
rect 142522 2592 142528 2604
rect 142580 2632 142586 2644
rect 143077 2635 143135 2641
rect 143077 2632 143089 2635
rect 142580 2604 143089 2632
rect 142580 2592 142586 2604
rect 143077 2601 143089 2604
rect 143123 2601 143135 2635
rect 143077 2595 143135 2601
rect 144178 2592 144184 2644
rect 144236 2632 144242 2644
rect 147033 2635 147091 2641
rect 144236 2604 145144 2632
rect 144236 2592 144242 2604
rect 143718 2564 143724 2576
rect 137020 2536 139900 2564
rect 143679 2536 143724 2564
rect 119341 2499 119399 2505
rect 119341 2496 119353 2499
rect 114051 2468 114508 2496
rect 118712 2468 119353 2496
rect 114051 2465 114063 2468
rect 114005 2459 114063 2465
rect 113821 2431 113879 2437
rect 113821 2428 113833 2431
rect 113192 2400 113833 2428
rect 113821 2397 113833 2400
rect 113867 2397 113879 2431
rect 113821 2391 113879 2397
rect 118533 2431 118591 2437
rect 118533 2397 118545 2431
rect 118579 2428 118591 2431
rect 118712 2428 118740 2468
rect 119341 2465 119353 2468
rect 119387 2496 119399 2499
rect 128326 2496 128354 2536
rect 143718 2524 143724 2536
rect 143776 2524 143782 2576
rect 129550 2496 129556 2508
rect 119387 2468 128354 2496
rect 129511 2468 129556 2496
rect 119387 2465 119399 2468
rect 119341 2459 119399 2465
rect 129550 2456 129556 2468
rect 129608 2496 129614 2508
rect 129608 2468 130424 2496
rect 129608 2456 129614 2468
rect 118579 2400 118740 2428
rect 118579 2397 118591 2400
rect 118533 2391 118591 2397
rect 118786 2388 118792 2440
rect 118844 2428 118850 2440
rect 118844 2400 118937 2428
rect 118844 2388 118850 2400
rect 120534 2388 120540 2440
rect 120592 2428 120598 2440
rect 121917 2431 121975 2437
rect 121917 2428 121929 2431
rect 120592 2400 121929 2428
rect 120592 2388 120598 2400
rect 121917 2397 121929 2400
rect 121963 2428 121975 2431
rect 126330 2428 126336 2440
rect 121963 2400 126336 2428
rect 121963 2397 121975 2400
rect 121917 2391 121975 2397
rect 126330 2388 126336 2400
rect 126388 2388 126394 2440
rect 130396 2437 130424 2468
rect 131114 2456 131120 2508
rect 131172 2496 131178 2508
rect 131577 2499 131635 2505
rect 131577 2496 131589 2499
rect 131172 2468 131589 2496
rect 131172 2456 131178 2468
rect 131577 2465 131589 2468
rect 131623 2465 131635 2499
rect 131577 2459 131635 2465
rect 133138 2456 133144 2508
rect 133196 2496 133202 2508
rect 133233 2499 133291 2505
rect 133233 2496 133245 2499
rect 133196 2468 133245 2496
rect 133196 2456 133202 2468
rect 133233 2465 133245 2468
rect 133279 2465 133291 2499
rect 135346 2496 135352 2508
rect 135307 2468 135352 2496
rect 133233 2459 133291 2465
rect 135346 2456 135352 2468
rect 135404 2456 135410 2508
rect 138474 2496 138480 2508
rect 137848 2468 138480 2496
rect 135622 2437 135628 2440
rect 130381 2431 130439 2437
rect 130381 2397 130393 2431
rect 130427 2397 130439 2431
rect 130381 2391 130439 2397
rect 130565 2431 130623 2437
rect 130565 2397 130577 2431
rect 130611 2397 130623 2431
rect 130565 2391 130623 2397
rect 135616 2391 135628 2437
rect 135680 2428 135686 2440
rect 135680 2400 135716 2428
rect 45428 2332 45692 2360
rect 75304 2363 75362 2369
rect 45428 2320 45434 2332
rect 75304 2329 75316 2363
rect 75350 2360 75362 2363
rect 75454 2360 75460 2372
rect 75350 2332 75460 2360
rect 75350 2329 75362 2332
rect 75304 2323 75362 2329
rect 75454 2320 75460 2332
rect 75512 2320 75518 2372
rect 82572 2363 82630 2369
rect 82572 2329 82584 2363
rect 82618 2360 82630 2363
rect 82998 2360 83004 2372
rect 82618 2332 83004 2360
rect 82618 2329 82630 2332
rect 82572 2323 82630 2329
rect 82998 2320 83004 2332
rect 83056 2320 83062 2372
rect 118804 2360 118832 2388
rect 119338 2360 119344 2372
rect 118804 2332 119344 2360
rect 119338 2320 119344 2332
rect 119396 2360 119402 2372
rect 119985 2363 120043 2369
rect 119985 2360 119997 2363
rect 119396 2332 119997 2360
rect 119396 2320 119402 2332
rect 119985 2329 119997 2332
rect 120031 2360 120043 2363
rect 127989 2363 128047 2369
rect 127989 2360 128001 2363
rect 120031 2332 128001 2360
rect 120031 2329 120043 2332
rect 119985 2323 120043 2329
rect 127989 2329 128001 2332
rect 128035 2360 128047 2363
rect 128998 2360 129004 2372
rect 128035 2332 129004 2360
rect 128035 2329 128047 2332
rect 127989 2323 128047 2329
rect 128998 2320 129004 2332
rect 129056 2320 129062 2372
rect 130580 2360 130608 2391
rect 135622 2388 135628 2391
rect 135680 2388 135686 2400
rect 131117 2363 131175 2369
rect 131117 2360 131129 2363
rect 130580 2332 131129 2360
rect 131117 2329 131129 2332
rect 131163 2360 131175 2363
rect 133138 2360 133144 2372
rect 131163 2332 133144 2360
rect 131163 2329 131175 2332
rect 131117 2323 131175 2329
rect 133138 2320 133144 2332
rect 133196 2320 133202 2372
rect 133500 2363 133558 2369
rect 133500 2329 133512 2363
rect 133546 2360 133558 2363
rect 137848 2360 137876 2468
rect 138474 2456 138480 2468
rect 138532 2456 138538 2508
rect 141970 2496 141976 2508
rect 141931 2468 141976 2496
rect 141970 2456 141976 2468
rect 142028 2456 142034 2508
rect 145116 2505 145144 2604
rect 147033 2601 147045 2635
rect 147079 2632 147091 2635
rect 148870 2632 148876 2644
rect 147079 2604 148876 2632
rect 147079 2601 147091 2604
rect 147033 2595 147091 2601
rect 148870 2592 148876 2604
rect 148928 2592 148934 2644
rect 148962 2592 148968 2644
rect 149020 2632 149026 2644
rect 151633 2635 151691 2641
rect 151633 2632 151645 2635
rect 149020 2604 151645 2632
rect 149020 2592 149026 2604
rect 151633 2601 151645 2604
rect 151679 2601 151691 2635
rect 152182 2632 152188 2644
rect 152143 2604 152188 2632
rect 151633 2595 151691 2601
rect 152182 2592 152188 2604
rect 152240 2592 152246 2644
rect 152734 2632 152740 2644
rect 152695 2604 152740 2632
rect 152734 2592 152740 2604
rect 152792 2592 152798 2644
rect 154485 2635 154543 2641
rect 154485 2601 154497 2635
rect 154531 2632 154543 2635
rect 159082 2632 159088 2644
rect 154531 2604 159088 2632
rect 154531 2601 154543 2604
rect 154485 2595 154543 2601
rect 159082 2592 159088 2604
rect 159140 2592 159146 2644
rect 149422 2524 149428 2576
rect 149480 2564 149486 2576
rect 150250 2564 150256 2576
rect 149480 2536 150256 2564
rect 149480 2524 149486 2536
rect 150250 2524 150256 2536
rect 150308 2524 150314 2576
rect 150434 2524 150440 2576
rect 150492 2564 150498 2576
rect 153381 2567 153439 2573
rect 153381 2564 153393 2567
rect 150492 2536 153393 2564
rect 150492 2524 150498 2536
rect 153381 2533 153393 2536
rect 153427 2533 153439 2567
rect 155770 2564 155776 2576
rect 153381 2527 153439 2533
rect 153488 2536 155776 2564
rect 145101 2499 145159 2505
rect 145101 2465 145113 2499
rect 145147 2496 145159 2499
rect 145650 2496 145656 2508
rect 145147 2468 145656 2496
rect 145147 2465 145159 2468
rect 145101 2459 145159 2465
rect 145650 2456 145656 2468
rect 145708 2456 145714 2508
rect 146938 2456 146944 2508
rect 146996 2496 147002 2508
rect 146996 2468 147996 2496
rect 146996 2456 147002 2468
rect 138658 2428 138664 2440
rect 138619 2400 138664 2428
rect 138658 2388 138664 2400
rect 138716 2388 138722 2440
rect 138753 2431 138811 2437
rect 138753 2397 138765 2431
rect 138799 2397 138811 2431
rect 138753 2391 138811 2397
rect 138937 2431 138995 2437
rect 138937 2397 138949 2431
rect 138983 2428 138995 2431
rect 141878 2428 141884 2440
rect 138983 2400 141884 2428
rect 138983 2397 138995 2400
rect 138937 2391 138995 2397
rect 133546 2332 137876 2360
rect 133546 2329 133558 2332
rect 133500 2323 133558 2329
rect 138014 2320 138020 2372
rect 138072 2360 138078 2372
rect 138768 2360 138796 2391
rect 141878 2388 141884 2400
rect 141936 2388 141942 2440
rect 144845 2431 144903 2437
rect 144845 2397 144857 2431
rect 144891 2428 144903 2431
rect 144891 2400 147536 2428
rect 144891 2397 144903 2400
rect 144845 2391 144903 2397
rect 140866 2360 140872 2372
rect 138072 2332 138796 2360
rect 139412 2332 140872 2360
rect 138072 2320 138078 2332
rect 31754 2292 31760 2304
rect 31715 2264 31760 2292
rect 31754 2252 31760 2264
rect 31812 2252 31818 2304
rect 32398 2292 32404 2304
rect 32359 2264 32404 2292
rect 32398 2252 32404 2264
rect 32456 2252 32462 2304
rect 117406 2292 117412 2304
rect 117367 2264 117412 2292
rect 117406 2252 117412 2264
rect 117464 2252 117470 2304
rect 120810 2292 120816 2304
rect 120771 2264 120816 2292
rect 120810 2252 120816 2264
rect 120868 2252 120874 2304
rect 121362 2292 121368 2304
rect 121323 2264 121368 2292
rect 121362 2252 121368 2264
rect 121420 2252 121426 2304
rect 123846 2292 123852 2304
rect 123807 2264 123852 2292
rect 123846 2252 123852 2264
rect 123904 2252 123910 2304
rect 124398 2292 124404 2304
rect 124359 2264 124404 2292
rect 124398 2252 124404 2264
rect 124456 2252 124462 2304
rect 125318 2292 125324 2304
rect 125279 2264 125324 2292
rect 125318 2252 125324 2264
rect 125376 2252 125382 2304
rect 128538 2292 128544 2304
rect 128499 2264 128544 2292
rect 128538 2252 128544 2264
rect 128596 2252 128602 2304
rect 135254 2252 135260 2304
rect 135312 2292 135318 2304
rect 136729 2295 136787 2301
rect 136729 2292 136741 2295
rect 135312 2264 136741 2292
rect 135312 2252 135318 2264
rect 136729 2261 136741 2264
rect 136775 2292 136787 2295
rect 139412 2292 139440 2332
rect 140866 2320 140872 2332
rect 140924 2320 140930 2372
rect 141694 2360 141700 2372
rect 141752 2369 141758 2372
rect 141752 2363 141786 2369
rect 141638 2332 141700 2360
rect 141694 2320 141700 2332
rect 141774 2360 141786 2363
rect 141970 2360 141976 2372
rect 141774 2332 141976 2360
rect 141774 2329 141786 2332
rect 141752 2323 141786 2329
rect 141752 2320 141758 2323
rect 141970 2320 141976 2332
rect 142028 2320 142034 2372
rect 145926 2369 145932 2372
rect 145920 2360 145932 2369
rect 145887 2332 145932 2360
rect 145920 2323 145932 2332
rect 145926 2320 145932 2323
rect 145984 2320 145990 2372
rect 147508 2360 147536 2400
rect 147674 2388 147680 2440
rect 147732 2428 147738 2440
rect 147732 2400 147777 2428
rect 147732 2388 147738 2400
rect 147508 2332 147674 2360
rect 140590 2292 140596 2304
rect 136775 2264 139440 2292
rect 140551 2264 140596 2292
rect 136775 2261 136787 2264
rect 136729 2255 136787 2261
rect 140590 2252 140596 2264
rect 140648 2252 140654 2304
rect 147490 2292 147496 2304
rect 147451 2264 147496 2292
rect 147490 2252 147496 2264
rect 147548 2252 147554 2304
rect 147646 2292 147674 2332
rect 147858 2292 147864 2304
rect 147646 2264 147864 2292
rect 147858 2252 147864 2264
rect 147916 2252 147922 2304
rect 147968 2292 147996 2468
rect 148042 2456 148048 2508
rect 148100 2496 148106 2508
rect 148229 2499 148287 2505
rect 148229 2496 148241 2499
rect 148100 2468 148241 2496
rect 148100 2456 148106 2468
rect 148229 2465 148241 2468
rect 148275 2465 148287 2499
rect 148229 2459 148287 2465
rect 149698 2456 149704 2508
rect 149756 2496 149762 2508
rect 151173 2499 151231 2505
rect 151173 2496 151185 2499
rect 149756 2468 151185 2496
rect 149756 2456 149762 2468
rect 151173 2465 151185 2468
rect 151219 2496 151231 2499
rect 153488 2496 153516 2536
rect 154114 2496 154120 2508
rect 151219 2468 153516 2496
rect 154075 2468 154120 2496
rect 151219 2465 151231 2468
rect 151173 2459 151231 2465
rect 154114 2456 154120 2468
rect 154172 2456 154178 2508
rect 155328 2505 155356 2536
rect 155770 2524 155776 2536
rect 155828 2524 155834 2576
rect 155954 2524 155960 2576
rect 156012 2564 156018 2576
rect 157426 2564 157432 2576
rect 156012 2536 157432 2564
rect 156012 2524 156018 2536
rect 157426 2524 157432 2536
rect 157484 2524 157490 2576
rect 155313 2499 155371 2505
rect 155313 2465 155325 2499
rect 155359 2465 155371 2499
rect 155313 2459 155371 2465
rect 157150 2456 157156 2508
rect 157208 2496 157214 2508
rect 157245 2499 157303 2505
rect 157245 2496 157257 2499
rect 157208 2468 157257 2496
rect 157208 2456 157214 2468
rect 157245 2465 157257 2468
rect 157291 2465 157303 2499
rect 157245 2459 157303 2465
rect 148778 2388 148784 2440
rect 148836 2428 148842 2440
rect 150069 2431 150127 2437
rect 150069 2428 150081 2431
rect 148836 2400 150081 2428
rect 148836 2388 148842 2400
rect 150069 2397 150081 2400
rect 150115 2397 150127 2431
rect 150069 2391 150127 2397
rect 150342 2388 150348 2440
rect 150400 2428 150406 2440
rect 150989 2431 151047 2437
rect 150989 2428 151001 2431
rect 150400 2400 151001 2428
rect 150400 2388 150406 2400
rect 150989 2397 151001 2400
rect 151035 2397 151047 2431
rect 154298 2428 154304 2440
rect 154259 2400 154304 2428
rect 150989 2391 151047 2397
rect 154298 2388 154304 2400
rect 154356 2388 154362 2440
rect 155126 2428 155132 2440
rect 155087 2400 155132 2428
rect 155126 2388 155132 2400
rect 155184 2388 155190 2440
rect 155862 2388 155868 2440
rect 155920 2428 155926 2440
rect 156141 2431 156199 2437
rect 156141 2428 156153 2431
rect 155920 2400 156153 2428
rect 155920 2388 155926 2400
rect 156141 2397 156153 2400
rect 156187 2397 156199 2431
rect 156141 2391 156199 2397
rect 156785 2431 156843 2437
rect 156785 2397 156797 2431
rect 156831 2397 156843 2431
rect 156785 2391 156843 2397
rect 148496 2363 148554 2369
rect 148496 2329 148508 2363
rect 148542 2360 148554 2363
rect 149146 2360 149152 2372
rect 148542 2332 149152 2360
rect 148542 2329 148554 2332
rect 148496 2323 148554 2329
rect 149146 2320 149152 2332
rect 149204 2320 149210 2372
rect 150805 2363 150863 2369
rect 150805 2360 150817 2363
rect 149256 2332 150817 2360
rect 149256 2292 149284 2332
rect 150805 2329 150817 2332
rect 150851 2329 150863 2363
rect 150805 2323 150863 2329
rect 151078 2320 151084 2372
rect 151136 2360 151142 2372
rect 154945 2363 155003 2369
rect 154945 2360 154957 2363
rect 151136 2332 154957 2360
rect 151136 2320 151142 2332
rect 154945 2329 154957 2332
rect 154991 2329 155003 2363
rect 156800 2360 156828 2391
rect 154945 2323 155003 2329
rect 155052 2332 156828 2360
rect 149606 2292 149612 2304
rect 147968 2264 149284 2292
rect 149567 2264 149612 2292
rect 149606 2252 149612 2264
rect 149664 2252 149670 2304
rect 151722 2252 151728 2304
rect 151780 2292 151786 2304
rect 155052 2292 155080 2332
rect 151780 2264 155080 2292
rect 151780 2252 151786 2264
rect 155862 2252 155868 2304
rect 155920 2292 155926 2304
rect 155957 2295 156015 2301
rect 155957 2292 155969 2295
rect 155920 2264 155969 2292
rect 155920 2252 155926 2264
rect 155957 2261 155969 2264
rect 156003 2261 156015 2295
rect 156598 2292 156604 2304
rect 156559 2264 156604 2292
rect 155957 2255 156015 2261
rect 156598 2252 156604 2264
rect 156656 2252 156662 2304
rect 157794 2292 157800 2304
rect 157755 2264 157800 2292
rect 157794 2252 157800 2264
rect 157852 2252 157858 2304
rect 1104 2202 159043 2224
rect 1104 2150 40394 2202
rect 40446 2150 40458 2202
rect 40510 2150 40522 2202
rect 40574 2150 40586 2202
rect 40638 2150 40650 2202
rect 40702 2150 79839 2202
rect 79891 2150 79903 2202
rect 79955 2150 79967 2202
rect 80019 2150 80031 2202
rect 80083 2150 80095 2202
rect 80147 2150 119284 2202
rect 119336 2150 119348 2202
rect 119400 2150 119412 2202
rect 119464 2150 119476 2202
rect 119528 2150 119540 2202
rect 119592 2150 158729 2202
rect 158781 2150 158793 2202
rect 158845 2150 158857 2202
rect 158909 2150 158921 2202
rect 158973 2150 158985 2202
rect 159037 2150 159043 2202
rect 1104 2128 159043 2150
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 32398 2088 32404 2100
rect 11020 2060 32404 2088
rect 11020 2048 11026 2060
rect 32398 2048 32404 2060
rect 32456 2048 32462 2100
rect 120166 2048 120172 2100
rect 120224 2088 120230 2100
rect 124398 2088 124404 2100
rect 120224 2060 124404 2088
rect 120224 2048 120230 2060
rect 124398 2048 124404 2060
rect 124456 2048 124462 2100
rect 128538 2048 128544 2100
rect 128596 2088 128602 2100
rect 145926 2088 145932 2100
rect 128596 2060 145932 2088
rect 128596 2048 128602 2060
rect 145926 2048 145932 2060
rect 145984 2048 145990 2100
rect 146662 2048 146668 2100
rect 146720 2088 146726 2100
rect 149054 2088 149060 2100
rect 146720 2060 149060 2088
rect 146720 2048 146726 2060
rect 149054 2048 149060 2060
rect 149112 2048 149118 2100
rect 150250 2048 150256 2100
rect 150308 2088 150314 2100
rect 156598 2088 156604 2100
rect 150308 2060 156604 2088
rect 150308 2048 150314 2060
rect 156598 2048 156604 2060
rect 156656 2048 156662 2100
rect 15562 1980 15568 2032
rect 15620 2020 15626 2032
rect 31754 2020 31760 2032
rect 15620 1992 31760 2020
rect 15620 1980 15626 1992
rect 31754 1980 31760 1992
rect 31812 1980 31818 2032
rect 121362 1980 121368 2032
rect 121420 2020 121426 2032
rect 134058 2020 134064 2032
rect 121420 1992 134064 2020
rect 121420 1980 121426 1992
rect 134058 1980 134064 1992
rect 134116 1980 134122 2032
rect 136634 1980 136640 2032
rect 136692 2020 136698 2032
rect 150342 2020 150348 2032
rect 136692 1992 150348 2020
rect 136692 1980 136698 1992
rect 150342 1980 150348 1992
rect 150400 1980 150406 2032
rect 106550 1912 106556 1964
rect 106608 1952 106614 1964
rect 123846 1952 123852 1964
rect 106608 1924 123852 1952
rect 106608 1912 106614 1924
rect 123846 1912 123852 1924
rect 123904 1912 123910 1964
rect 124858 1912 124864 1964
rect 124916 1952 124922 1964
rect 147490 1952 147496 1964
rect 124916 1924 147496 1952
rect 124916 1912 124922 1924
rect 147490 1912 147496 1924
rect 147548 1912 147554 1964
rect 149146 1912 149152 1964
rect 149204 1952 149210 1964
rect 159174 1952 159180 1964
rect 149204 1924 159180 1952
rect 149204 1912 149210 1924
rect 159174 1912 159180 1924
rect 159232 1912 159238 1964
rect 123864 1884 123892 1912
rect 146110 1884 146116 1896
rect 123864 1856 146116 1884
rect 146110 1844 146116 1856
rect 146168 1884 146174 1896
rect 146662 1884 146668 1896
rect 146168 1856 146668 1884
rect 146168 1844 146174 1856
rect 146662 1844 146668 1856
rect 146720 1844 146726 1896
rect 114462 1776 114468 1828
rect 114520 1816 114526 1828
rect 114520 1788 120672 1816
rect 114520 1776 114526 1788
rect 115566 1640 115572 1692
rect 115624 1680 115630 1692
rect 115624 1652 118694 1680
rect 115624 1640 115630 1652
rect 118666 1476 118694 1652
rect 120644 1544 120672 1788
rect 124398 1776 124404 1828
rect 124456 1816 124462 1828
rect 130838 1816 130844 1828
rect 124456 1788 130844 1816
rect 124456 1776 124462 1788
rect 130838 1776 130844 1788
rect 130896 1776 130902 1828
rect 141970 1776 141976 1828
rect 142028 1816 142034 1828
rect 147766 1816 147772 1828
rect 142028 1788 147772 1816
rect 142028 1776 142034 1788
rect 147766 1776 147772 1788
rect 147824 1776 147830 1828
rect 147858 1776 147864 1828
rect 147916 1816 147922 1828
rect 156046 1816 156052 1828
rect 147916 1788 156052 1816
rect 147916 1776 147922 1788
rect 156046 1776 156052 1788
rect 156104 1776 156110 1828
rect 123018 1708 123024 1760
rect 123076 1748 123082 1760
rect 140590 1748 140596 1760
rect 123076 1720 140596 1748
rect 123076 1708 123082 1720
rect 140590 1708 140596 1720
rect 140648 1708 140654 1760
rect 143626 1708 143632 1760
rect 143684 1748 143690 1760
rect 154942 1748 154948 1760
rect 143684 1720 154948 1748
rect 143684 1708 143690 1720
rect 154942 1708 154948 1720
rect 155000 1708 155006 1760
rect 125318 1640 125324 1692
rect 125376 1680 125382 1692
rect 142798 1680 142804 1692
rect 125376 1652 142804 1680
rect 125376 1640 125382 1652
rect 142798 1640 142804 1652
rect 142856 1640 142862 1692
rect 146202 1640 146208 1692
rect 146260 1680 146266 1692
rect 155126 1680 155132 1692
rect 146260 1652 155132 1680
rect 146260 1640 146266 1652
rect 155126 1640 155132 1652
rect 155184 1640 155190 1692
rect 120810 1572 120816 1624
rect 120868 1612 120874 1624
rect 136082 1612 136088 1624
rect 120868 1584 136088 1612
rect 120868 1572 120874 1584
rect 136082 1572 136088 1584
rect 136140 1572 136146 1624
rect 143994 1572 144000 1624
rect 144052 1612 144058 1624
rect 155954 1612 155960 1624
rect 144052 1584 155960 1612
rect 144052 1572 144058 1584
rect 155954 1572 155960 1584
rect 156012 1572 156018 1624
rect 126974 1544 126980 1556
rect 120644 1516 126980 1544
rect 126974 1504 126980 1516
rect 127032 1504 127038 1556
rect 147766 1504 147772 1556
rect 147824 1544 147830 1556
rect 156966 1544 156972 1556
rect 147824 1516 156972 1544
rect 147824 1504 147830 1516
rect 156966 1504 156972 1516
rect 157024 1504 157030 1556
rect 125318 1476 125324 1488
rect 118666 1448 125324 1476
rect 125318 1436 125324 1448
rect 125376 1436 125382 1488
rect 110230 1300 110236 1352
rect 110288 1340 110294 1352
rect 151998 1340 152004 1352
rect 110288 1312 152004 1340
rect 110288 1300 110294 1312
rect 151998 1300 152004 1312
rect 152056 1300 152062 1352
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 150894 1272 150900 1284
rect 115256 1244 150900 1272
rect 115256 1232 115262 1244
rect 150894 1232 150900 1244
rect 150952 1232 150958 1284
rect 121178 1164 121184 1216
rect 121236 1204 121242 1216
rect 155402 1204 155408 1216
rect 121236 1176 155408 1204
rect 121236 1164 121242 1176
rect 155402 1164 155408 1176
rect 155460 1164 155466 1216
rect 119798 1096 119804 1148
rect 119856 1136 119862 1148
rect 150802 1136 150808 1148
rect 119856 1108 150808 1136
rect 119856 1096 119862 1108
rect 150802 1096 150808 1108
rect 150860 1096 150866 1148
rect 101950 1028 101956 1080
rect 102008 1068 102014 1080
rect 128446 1068 128452 1080
rect 102008 1040 128452 1068
rect 102008 1028 102014 1040
rect 128446 1028 128452 1040
rect 128504 1028 128510 1080
rect 129182 1028 129188 1080
rect 129240 1068 129246 1080
rect 151170 1068 151176 1080
rect 129240 1040 151176 1068
rect 129240 1028 129246 1040
rect 151170 1028 151176 1040
rect 151228 1028 151234 1080
rect 113542 960 113548 1012
rect 113600 1000 113606 1012
rect 138106 1000 138112 1012
rect 113600 972 138112 1000
rect 113600 960 113606 972
rect 138106 960 138112 972
rect 138164 960 138170 1012
<< via1 >>
rect 146484 15036 146536 15088
rect 154396 15036 154448 15088
rect 145932 14968 145984 15020
rect 154304 14968 154356 15020
rect 96436 14900 96488 14952
rect 149336 14900 149388 14952
rect 118056 14832 118108 14884
rect 150716 14832 150768 14884
rect 109316 14764 109368 14816
rect 141884 14764 141936 14816
rect 146024 14764 146076 14816
rect 152464 14764 152516 14816
rect 114192 14696 114244 14748
rect 157432 14696 157484 14748
rect 119068 14628 119120 14680
rect 152648 14628 152700 14680
rect 130660 14560 130712 14612
rect 156696 14560 156748 14612
rect 134616 14492 134668 14544
rect 149520 14492 149572 14544
rect 149980 14492 150032 14544
rect 154948 14492 155000 14544
rect 129096 14424 129148 14476
rect 150808 14424 150860 14476
rect 107476 14356 107528 14408
rect 132960 14356 133012 14408
rect 134524 14356 134576 14408
rect 154856 14356 154908 14408
rect 125876 14288 125928 14340
rect 153384 14288 153436 14340
rect 124312 14220 124364 14272
rect 152556 14220 152608 14272
rect 129188 14152 129240 14204
rect 156052 14152 156104 14204
rect 129556 14084 129608 14136
rect 153200 14084 153252 14136
rect 51080 14016 51132 14068
rect 53748 14016 53800 14068
rect 138480 14016 138532 14068
rect 155960 14016 156012 14068
rect 10048 13948 10100 14000
rect 11244 13948 11296 14000
rect 12532 13880 12584 13932
rect 15292 13880 15344 13932
rect 4068 13812 4120 13864
rect 43904 13880 43956 13932
rect 47124 13880 47176 13932
rect 50712 13880 50764 13932
rect 10416 13744 10468 13796
rect 15200 13744 15252 13796
rect 15292 13744 15344 13796
rect 19616 13744 19668 13796
rect 7840 13676 7892 13728
rect 12716 13676 12768 13728
rect 17408 13676 17460 13728
rect 24584 13744 24636 13796
rect 24768 13744 24820 13796
rect 28264 13744 28316 13796
rect 36268 13744 36320 13796
rect 41328 13744 41380 13796
rect 41420 13744 41472 13796
rect 22376 13676 22428 13728
rect 27896 13676 27948 13728
rect 36176 13676 36228 13728
rect 42340 13676 42392 13728
rect 42524 13744 42576 13796
rect 43168 13744 43220 13796
rect 45100 13744 45152 13796
rect 46664 13744 46716 13796
rect 46940 13744 46992 13796
rect 50620 13744 50672 13796
rect 45560 13676 45612 13728
rect 46112 13676 46164 13728
rect 48136 13676 48188 13728
rect 50712 13676 50764 13728
rect 65524 13880 65576 13932
rect 60556 13744 60608 13796
rect 61384 13744 61436 13796
rect 65892 13744 65944 13796
rect 100760 13948 100812 14000
rect 128912 13948 128964 14000
rect 129004 13948 129056 14000
rect 104256 13880 104308 13932
rect 133052 13880 133104 13932
rect 80612 13812 80664 13864
rect 94044 13744 94096 13796
rect 95792 13744 95844 13796
rect 95884 13744 95936 13796
rect 98736 13744 98788 13796
rect 102324 13744 102376 13796
rect 104348 13744 104400 13796
rect 106648 13744 106700 13796
rect 106832 13744 106884 13796
rect 115664 13744 115716 13796
rect 123024 13812 123076 13864
rect 66628 13676 66680 13728
rect 73988 13676 74040 13728
rect 82084 13676 82136 13728
rect 82176 13676 82228 13728
rect 87880 13676 87932 13728
rect 88064 13676 88116 13728
rect 89720 13676 89772 13728
rect 90824 13676 90876 13728
rect 94872 13676 94924 13728
rect 104164 13676 104216 13728
rect 109592 13676 109644 13728
rect 109684 13676 109736 13728
rect 122104 13744 122156 13796
rect 127348 13744 127400 13796
rect 138756 13948 138808 14000
rect 157616 13948 157668 14000
rect 138020 13880 138072 13932
rect 140596 13744 140648 13796
rect 141148 13744 141200 13796
rect 146944 13812 146996 13864
rect 148416 13880 148468 13932
rect 149980 13812 150032 13864
rect 150072 13812 150124 13864
rect 152280 13812 152332 13864
rect 152464 13880 152516 13932
rect 158076 13880 158128 13932
rect 145380 13744 145432 13796
rect 153568 13744 153620 13796
rect 156144 13744 156196 13796
rect 120172 13676 120224 13728
rect 127532 13676 127584 13728
rect 139584 13676 139636 13728
rect 146208 13676 146260 13728
rect 149244 13676 149296 13728
rect 153292 13676 153344 13728
rect 20672 13574 20724 13626
rect 20736 13574 20788 13626
rect 20800 13574 20852 13626
rect 20864 13574 20916 13626
rect 20928 13574 20980 13626
rect 60117 13574 60169 13626
rect 60181 13574 60233 13626
rect 60245 13574 60297 13626
rect 60309 13574 60361 13626
rect 60373 13574 60425 13626
rect 99562 13574 99614 13626
rect 99626 13574 99678 13626
rect 99690 13574 99742 13626
rect 99754 13574 99806 13626
rect 99818 13574 99870 13626
rect 139007 13574 139059 13626
rect 139071 13574 139123 13626
rect 139135 13574 139187 13626
rect 139199 13574 139251 13626
rect 139263 13574 139315 13626
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 9220 13472 9272 13524
rect 12348 13472 12400 13524
rect 10048 13404 10100 13456
rect 15660 13472 15712 13524
rect 17868 13472 17920 13524
rect 18420 13472 18472 13524
rect 19524 13472 19576 13524
rect 21732 13472 21784 13524
rect 14556 13404 14608 13456
rect 21180 13404 21232 13456
rect 21640 13404 21692 13456
rect 12532 13336 12584 13388
rect 22192 13472 22244 13524
rect 23940 13472 23992 13524
rect 24584 13472 24636 13524
rect 27436 13472 27488 13524
rect 28080 13472 28132 13524
rect 28908 13472 28960 13524
rect 30564 13472 30616 13524
rect 32772 13515 32824 13524
rect 32772 13481 32781 13515
rect 32781 13481 32815 13515
rect 32815 13481 32824 13515
rect 32772 13472 32824 13481
rect 34428 13472 34480 13524
rect 22008 13404 22060 13456
rect 22284 13404 22336 13456
rect 25228 13404 25280 13456
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 10232 13268 10284 13320
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11888 13268 11940 13320
rect 12164 13268 12216 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 15752 13268 15804 13320
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 18604 13268 18656 13320
rect 10784 13132 10836 13184
rect 13912 13200 13964 13252
rect 15108 13200 15160 13252
rect 15292 13200 15344 13252
rect 17684 13200 17736 13252
rect 19892 13268 19944 13320
rect 20352 13268 20404 13320
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 24952 13336 25004 13388
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 21364 13200 21416 13252
rect 22192 13200 22244 13252
rect 25044 13268 25096 13320
rect 25136 13268 25188 13320
rect 25780 13268 25832 13320
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 16396 13132 16448 13184
rect 21548 13132 21600 13184
rect 29276 13404 29328 13456
rect 35532 13472 35584 13524
rect 39396 13472 39448 13524
rect 39856 13472 39908 13524
rect 42984 13472 43036 13524
rect 26792 13336 26844 13388
rect 27528 13268 27580 13320
rect 27712 13336 27764 13388
rect 30104 13336 30156 13388
rect 28264 13268 28316 13320
rect 29000 13268 29052 13320
rect 32588 13311 32640 13320
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 24952 13132 25004 13184
rect 26516 13132 26568 13184
rect 30472 13243 30524 13252
rect 30472 13209 30506 13243
rect 30506 13209 30524 13243
rect 30472 13200 30524 13209
rect 26700 13132 26752 13184
rect 32588 13277 32597 13311
rect 32597 13277 32631 13311
rect 32631 13277 32640 13311
rect 32588 13268 32640 13277
rect 34796 13268 34848 13320
rect 36176 13268 36228 13320
rect 43076 13404 43128 13456
rect 38752 13311 38804 13320
rect 34060 13200 34112 13252
rect 34428 13200 34480 13252
rect 38752 13277 38761 13311
rect 38761 13277 38795 13311
rect 38795 13277 38804 13311
rect 38752 13268 38804 13277
rect 35440 13132 35492 13184
rect 36544 13132 36596 13184
rect 37832 13132 37884 13184
rect 41052 13336 41104 13388
rect 50896 13472 50948 13524
rect 45560 13404 45612 13456
rect 46664 13404 46716 13456
rect 49792 13404 49844 13456
rect 39488 13311 39540 13320
rect 39488 13277 39497 13311
rect 39497 13277 39531 13311
rect 39531 13277 39540 13311
rect 39488 13268 39540 13277
rect 40316 13268 40368 13320
rect 41144 13268 41196 13320
rect 52920 13336 52972 13388
rect 55864 13404 55916 13456
rect 60648 13404 60700 13456
rect 41328 13268 41380 13320
rect 41512 13268 41564 13320
rect 41880 13311 41932 13320
rect 41880 13277 41889 13311
rect 41889 13277 41923 13311
rect 41923 13277 41932 13311
rect 41880 13268 41932 13277
rect 42708 13268 42760 13320
rect 45928 13268 45980 13320
rect 42432 13200 42484 13252
rect 40132 13132 40184 13184
rect 43168 13200 43220 13252
rect 43720 13200 43772 13252
rect 43812 13200 43864 13252
rect 42800 13175 42852 13184
rect 42800 13141 42809 13175
rect 42809 13141 42843 13175
rect 42843 13141 42852 13175
rect 42800 13132 42852 13141
rect 43628 13132 43680 13184
rect 45560 13132 45612 13184
rect 47216 13268 47268 13320
rect 49700 13268 49752 13320
rect 49884 13268 49936 13320
rect 48320 13200 48372 13252
rect 53564 13311 53616 13320
rect 53564 13277 53573 13311
rect 53573 13277 53607 13311
rect 53607 13277 53616 13311
rect 53564 13268 53616 13277
rect 49792 13132 49844 13184
rect 50712 13132 50764 13184
rect 50804 13132 50856 13184
rect 55404 13268 55456 13320
rect 55588 13268 55640 13320
rect 56692 13268 56744 13320
rect 58624 13268 58676 13320
rect 56048 13200 56100 13252
rect 53012 13132 53064 13184
rect 60372 13200 60424 13252
rect 60648 13268 60700 13320
rect 60740 13268 60792 13320
rect 60832 13311 60884 13320
rect 60832 13277 60841 13311
rect 60841 13277 60875 13311
rect 60875 13277 60884 13311
rect 63408 13311 63460 13320
rect 60832 13268 60884 13277
rect 63408 13277 63417 13311
rect 63417 13277 63451 13311
rect 63451 13277 63460 13311
rect 63408 13268 63460 13277
rect 61108 13243 61160 13252
rect 61108 13209 61142 13243
rect 61142 13209 61160 13243
rect 63592 13268 63644 13320
rect 65524 13268 65576 13320
rect 65616 13268 65668 13320
rect 61108 13200 61160 13209
rect 57520 13175 57572 13184
rect 57520 13141 57529 13175
rect 57529 13141 57563 13175
rect 57563 13141 57572 13175
rect 57520 13132 57572 13141
rect 58808 13132 58860 13184
rect 60648 13132 60700 13184
rect 65156 13243 65208 13252
rect 65156 13209 65165 13243
rect 65165 13209 65199 13243
rect 65199 13209 65208 13243
rect 65156 13200 65208 13209
rect 66444 13472 66496 13524
rect 66628 13515 66680 13524
rect 66628 13481 66637 13515
rect 66637 13481 66671 13515
rect 66671 13481 66680 13515
rect 66628 13472 66680 13481
rect 68100 13472 68152 13524
rect 69204 13472 69256 13524
rect 69940 13472 69992 13524
rect 70860 13472 70912 13524
rect 71320 13515 71372 13524
rect 71320 13481 71329 13515
rect 71329 13481 71363 13515
rect 71363 13481 71372 13515
rect 71320 13472 71372 13481
rect 72056 13515 72108 13524
rect 72056 13481 72065 13515
rect 72065 13481 72099 13515
rect 72099 13481 72108 13515
rect 72056 13472 72108 13481
rect 72792 13515 72844 13524
rect 72792 13481 72801 13515
rect 72801 13481 72835 13515
rect 72835 13481 72844 13515
rect 72792 13472 72844 13481
rect 73896 13515 73948 13524
rect 73896 13481 73905 13515
rect 73905 13481 73939 13515
rect 73939 13481 73948 13515
rect 73896 13472 73948 13481
rect 74632 13515 74684 13524
rect 74632 13481 74641 13515
rect 74641 13481 74675 13515
rect 74675 13481 74684 13515
rect 74632 13472 74684 13481
rect 75460 13515 75512 13524
rect 75460 13481 75469 13515
rect 75469 13481 75503 13515
rect 75503 13481 75512 13515
rect 75460 13472 75512 13481
rect 76932 13472 76984 13524
rect 78036 13515 78088 13524
rect 78036 13481 78045 13515
rect 78045 13481 78079 13515
rect 78079 13481 78088 13515
rect 78036 13472 78088 13481
rect 79140 13472 79192 13524
rect 79784 13515 79836 13524
rect 79784 13481 79793 13515
rect 79793 13481 79827 13515
rect 79827 13481 79836 13515
rect 79784 13472 79836 13481
rect 80244 13472 80296 13524
rect 80796 13472 80848 13524
rect 81900 13472 81952 13524
rect 83004 13472 83056 13524
rect 84108 13472 84160 13524
rect 84568 13472 84620 13524
rect 84660 13472 84712 13524
rect 65892 13404 65944 13456
rect 73988 13336 74040 13388
rect 66904 13243 66956 13252
rect 66904 13209 66913 13243
rect 66913 13209 66947 13243
rect 66947 13209 66956 13243
rect 66904 13200 66956 13209
rect 68836 13268 68888 13320
rect 69664 13311 69716 13320
rect 69664 13277 69673 13311
rect 69673 13277 69707 13311
rect 69707 13277 69716 13311
rect 69664 13268 69716 13277
rect 71136 13268 71188 13320
rect 71688 13268 71740 13320
rect 70952 13200 71004 13252
rect 73896 13268 73948 13320
rect 79968 13336 80020 13388
rect 81348 13404 81400 13456
rect 83188 13404 83240 13456
rect 88708 13472 88760 13524
rect 88800 13472 88852 13524
rect 91008 13472 91060 13524
rect 95148 13472 95200 13524
rect 98000 13472 98052 13524
rect 102876 13472 102928 13524
rect 104808 13472 104860 13524
rect 106648 13472 106700 13524
rect 107660 13472 107712 13524
rect 107844 13472 107896 13524
rect 88616 13404 88668 13456
rect 91100 13404 91152 13456
rect 93216 13404 93268 13456
rect 95792 13404 95844 13456
rect 97080 13404 97132 13456
rect 98460 13404 98512 13456
rect 101220 13404 101272 13456
rect 103520 13404 103572 13456
rect 108948 13472 109000 13524
rect 110604 13472 110656 13524
rect 112812 13472 112864 13524
rect 113916 13472 113968 13524
rect 115572 13472 115624 13524
rect 109776 13404 109828 13456
rect 111432 13404 111484 13456
rect 114468 13404 114520 13456
rect 116676 13472 116728 13524
rect 118332 13472 118384 13524
rect 120540 13472 120592 13524
rect 122748 13472 122800 13524
rect 125508 13472 125560 13524
rect 126888 13472 126940 13524
rect 75092 13268 75144 13320
rect 75368 13268 75420 13320
rect 77116 13268 77168 13320
rect 77208 13311 77260 13320
rect 77208 13277 77235 13311
rect 77235 13277 77260 13311
rect 77208 13268 77260 13277
rect 75736 13200 75788 13252
rect 75828 13200 75880 13252
rect 64144 13132 64196 13184
rect 65892 13132 65944 13184
rect 65984 13132 66036 13184
rect 79140 13311 79192 13320
rect 79140 13277 79149 13311
rect 79149 13277 79183 13311
rect 79183 13277 79192 13311
rect 79140 13268 79192 13277
rect 77576 13132 77628 13184
rect 81072 13268 81124 13320
rect 81164 13268 81216 13320
rect 82268 13311 82320 13320
rect 82268 13277 82277 13311
rect 82277 13277 82311 13311
rect 82311 13277 82320 13311
rect 82268 13268 82320 13277
rect 84016 13268 84068 13320
rect 84292 13268 84344 13320
rect 88432 13311 88484 13320
rect 88432 13277 88441 13311
rect 88441 13277 88475 13311
rect 88475 13277 88484 13311
rect 88432 13268 88484 13277
rect 89444 13268 89496 13320
rect 89720 13268 89772 13320
rect 90548 13268 90600 13320
rect 90824 13311 90876 13320
rect 90824 13277 90833 13311
rect 90833 13277 90867 13311
rect 90867 13277 90876 13311
rect 90824 13268 90876 13277
rect 91376 13268 91428 13320
rect 84568 13132 84620 13184
rect 85488 13132 85540 13184
rect 88064 13200 88116 13252
rect 88616 13200 88668 13252
rect 89260 13200 89312 13252
rect 92480 13200 92532 13252
rect 95056 13336 95108 13388
rect 94412 13311 94464 13320
rect 94412 13277 94421 13311
rect 94421 13277 94455 13311
rect 94455 13277 94464 13311
rect 94412 13268 94464 13277
rect 95424 13268 95476 13320
rect 95608 13268 95660 13320
rect 104164 13336 104216 13388
rect 95884 13311 95936 13320
rect 95884 13277 95893 13311
rect 95893 13277 95927 13311
rect 95927 13277 95936 13311
rect 95884 13268 95936 13277
rect 96988 13311 97040 13320
rect 96988 13277 96997 13311
rect 96997 13277 97031 13311
rect 97031 13277 97040 13311
rect 96988 13268 97040 13277
rect 97724 13311 97776 13320
rect 97724 13277 97733 13311
rect 97733 13277 97767 13311
rect 97767 13277 97776 13311
rect 97724 13268 97776 13277
rect 96620 13200 96672 13252
rect 96896 13200 96948 13252
rect 99472 13268 99524 13320
rect 100024 13311 100076 13320
rect 100024 13277 100033 13311
rect 100033 13277 100067 13311
rect 100067 13277 100076 13311
rect 100024 13268 100076 13277
rect 101864 13268 101916 13320
rect 102324 13311 102376 13320
rect 102324 13277 102333 13311
rect 102333 13277 102367 13311
rect 102367 13277 102376 13311
rect 102324 13268 102376 13277
rect 102508 13268 102560 13320
rect 103060 13268 103112 13320
rect 104072 13268 104124 13320
rect 110512 13336 110564 13388
rect 86684 13132 86736 13184
rect 88892 13132 88944 13184
rect 88984 13175 89036 13184
rect 88984 13141 88993 13175
rect 88993 13141 89027 13175
rect 89027 13141 89036 13175
rect 88984 13132 89036 13141
rect 91284 13132 91336 13184
rect 95056 13132 95108 13184
rect 96712 13132 96764 13184
rect 96804 13132 96856 13184
rect 99012 13132 99064 13184
rect 102968 13132 103020 13184
rect 103060 13132 103112 13184
rect 107016 13268 107068 13320
rect 109040 13268 109092 13320
rect 109684 13268 109736 13320
rect 110052 13268 110104 13320
rect 111340 13311 111392 13320
rect 108580 13200 108632 13252
rect 106372 13132 106424 13184
rect 110420 13132 110472 13184
rect 111340 13277 111349 13311
rect 111349 13277 111383 13311
rect 111383 13277 111392 13311
rect 111340 13268 111392 13277
rect 112444 13311 112496 13320
rect 112444 13277 112453 13311
rect 112453 13277 112487 13311
rect 112487 13277 112496 13311
rect 112444 13268 112496 13277
rect 112996 13336 113048 13388
rect 114468 13268 114520 13320
rect 114652 13268 114704 13320
rect 115664 13268 115716 13320
rect 117228 13336 117280 13388
rect 119160 13404 119212 13456
rect 117964 13336 118016 13388
rect 121368 13336 121420 13388
rect 122012 13336 122064 13388
rect 116584 13268 116636 13320
rect 112628 13200 112680 13252
rect 112996 13200 113048 13252
rect 113088 13200 113140 13252
rect 117136 13200 117188 13252
rect 117320 13311 117372 13320
rect 117320 13277 117329 13311
rect 117329 13277 117363 13311
rect 117363 13277 117372 13311
rect 117320 13268 117372 13277
rect 119896 13268 119948 13320
rect 120816 13268 120868 13320
rect 120908 13311 120960 13320
rect 120908 13277 120917 13311
rect 120917 13277 120951 13311
rect 120951 13277 120960 13311
rect 120908 13268 120960 13277
rect 122104 13268 122156 13320
rect 113180 13132 113232 13184
rect 114744 13132 114796 13184
rect 117320 13132 117372 13184
rect 119160 13132 119212 13184
rect 123484 13200 123536 13252
rect 124680 13404 124732 13456
rect 126060 13404 126112 13456
rect 127992 13472 128044 13524
rect 129924 13472 129976 13524
rect 131120 13472 131172 13524
rect 132500 13472 132552 13524
rect 133236 13472 133288 13524
rect 128820 13404 128872 13456
rect 124772 13336 124824 13388
rect 125600 13336 125652 13388
rect 125324 13311 125376 13320
rect 125324 13277 125333 13311
rect 125333 13277 125367 13311
rect 125367 13277 125376 13311
rect 125324 13268 125376 13277
rect 127440 13336 127492 13388
rect 127532 13336 127584 13388
rect 130384 13336 130436 13388
rect 127716 13268 127768 13320
rect 127900 13311 127952 13320
rect 127900 13277 127909 13311
rect 127909 13277 127943 13311
rect 127943 13277 127952 13311
rect 127900 13268 127952 13277
rect 128728 13268 128780 13320
rect 130108 13268 130160 13320
rect 132684 13404 132736 13456
rect 134340 13472 134392 13524
rect 135720 13472 135772 13524
rect 136364 13472 136416 13524
rect 137100 13472 137152 13524
rect 138204 13472 138256 13524
rect 138848 13472 138900 13524
rect 139860 13472 139912 13524
rect 140688 13472 140740 13524
rect 141516 13472 141568 13524
rect 138388 13404 138440 13456
rect 138572 13404 138624 13456
rect 141148 13404 141200 13456
rect 141240 13404 141292 13456
rect 142528 13472 142580 13524
rect 148048 13472 148100 13524
rect 148600 13472 148652 13524
rect 149888 13472 149940 13524
rect 131948 13311 132000 13320
rect 131948 13277 131957 13311
rect 131957 13277 131991 13311
rect 131991 13277 132000 13311
rect 135352 13336 135404 13388
rect 131948 13268 132000 13277
rect 132408 13268 132460 13320
rect 124312 13175 124364 13184
rect 124312 13141 124321 13175
rect 124321 13141 124355 13175
rect 124355 13141 124364 13175
rect 124312 13132 124364 13141
rect 124404 13132 124456 13184
rect 128636 13132 128688 13184
rect 128820 13132 128872 13184
rect 129096 13132 129148 13184
rect 131212 13132 131264 13184
rect 133880 13268 133932 13320
rect 135628 13311 135680 13320
rect 135628 13277 135637 13311
rect 135637 13277 135671 13311
rect 135671 13277 135680 13311
rect 135628 13268 135680 13277
rect 136088 13311 136140 13320
rect 136088 13277 136097 13311
rect 136097 13277 136131 13311
rect 136131 13277 136140 13311
rect 136088 13268 136140 13277
rect 136732 13336 136784 13388
rect 138112 13268 138164 13320
rect 139400 13311 139452 13320
rect 139400 13277 139409 13311
rect 139409 13277 139443 13311
rect 139443 13277 139452 13311
rect 139400 13268 139452 13277
rect 140780 13311 140832 13320
rect 140780 13277 140789 13311
rect 140789 13277 140823 13311
rect 140823 13277 140832 13311
rect 140780 13268 140832 13277
rect 140872 13268 140924 13320
rect 133604 13200 133656 13252
rect 139584 13200 139636 13252
rect 139676 13200 139728 13252
rect 147404 13404 147456 13456
rect 146944 13336 146996 13388
rect 148140 13404 148192 13456
rect 151268 13472 151320 13524
rect 151820 13472 151872 13524
rect 150808 13447 150860 13456
rect 149244 13336 149296 13388
rect 150808 13413 150817 13447
rect 150817 13413 150851 13447
rect 150851 13413 150860 13447
rect 150808 13404 150860 13413
rect 153568 13515 153620 13524
rect 153568 13481 153577 13515
rect 153577 13481 153611 13515
rect 153611 13481 153620 13515
rect 154304 13515 154356 13524
rect 153568 13472 153620 13481
rect 154304 13481 154313 13515
rect 154313 13481 154347 13515
rect 154347 13481 154356 13515
rect 154304 13472 154356 13481
rect 155868 13472 155920 13524
rect 155684 13404 155736 13456
rect 155776 13404 155828 13456
rect 152372 13336 152424 13388
rect 156788 13336 156840 13388
rect 143356 13268 143408 13320
rect 147496 13268 147548 13320
rect 144000 13243 144052 13252
rect 144000 13209 144034 13243
rect 144034 13209 144052 13243
rect 144000 13200 144052 13209
rect 133144 13132 133196 13184
rect 135168 13132 135220 13184
rect 135536 13132 135588 13184
rect 142712 13132 142764 13184
rect 143816 13132 143868 13184
rect 145840 13200 145892 13252
rect 146208 13243 146260 13252
rect 146208 13209 146242 13243
rect 146242 13209 146260 13243
rect 146208 13200 146260 13209
rect 146484 13200 146536 13252
rect 145104 13175 145156 13184
rect 145104 13141 145113 13175
rect 145113 13141 145147 13175
rect 145147 13141 145156 13175
rect 145104 13132 145156 13141
rect 148600 13200 148652 13252
rect 149244 13200 149296 13252
rect 150900 13268 150952 13320
rect 152464 13268 152516 13320
rect 152832 13311 152884 13320
rect 152832 13277 152841 13311
rect 152841 13277 152875 13311
rect 152875 13277 152884 13311
rect 152832 13268 152884 13277
rect 153384 13311 153436 13320
rect 153384 13277 153393 13311
rect 153393 13277 153427 13311
rect 153427 13277 153436 13311
rect 153384 13268 153436 13277
rect 153476 13268 153528 13320
rect 154856 13311 154908 13320
rect 154856 13277 154865 13311
rect 154865 13277 154899 13311
rect 154899 13277 154908 13311
rect 154856 13268 154908 13277
rect 155960 13311 156012 13320
rect 155960 13277 155969 13311
rect 155969 13277 156003 13311
rect 156003 13277 156012 13311
rect 155960 13268 156012 13277
rect 156696 13311 156748 13320
rect 156696 13277 156705 13311
rect 156705 13277 156739 13311
rect 156739 13277 156748 13311
rect 156696 13268 156748 13277
rect 157432 13311 157484 13320
rect 157432 13277 157441 13311
rect 157441 13277 157475 13311
rect 157475 13277 157484 13311
rect 157432 13268 157484 13277
rect 149152 13132 149204 13184
rect 151820 13132 151872 13184
rect 152740 13200 152792 13252
rect 153292 13200 153344 13252
rect 152372 13132 152424 13184
rect 153200 13132 153252 13184
rect 153752 13132 153804 13184
rect 154212 13132 154264 13184
rect 154396 13132 154448 13184
rect 40394 13030 40446 13082
rect 40458 13030 40510 13082
rect 40522 13030 40574 13082
rect 40586 13030 40638 13082
rect 40650 13030 40702 13082
rect 79839 13030 79891 13082
rect 79903 13030 79955 13082
rect 79967 13030 80019 13082
rect 80031 13030 80083 13082
rect 80095 13030 80147 13082
rect 119284 13030 119336 13082
rect 119348 13030 119400 13082
rect 119412 13030 119464 13082
rect 119476 13030 119528 13082
rect 119540 13030 119592 13082
rect 158729 13030 158781 13082
rect 158793 13030 158845 13082
rect 158857 13030 158909 13082
rect 158921 13030 158973 13082
rect 158985 13030 159037 13082
rect 9404 12928 9456 12980
rect 10140 12928 10192 12980
rect 11796 12928 11848 12980
rect 11980 12928 12032 12980
rect 13912 12928 13964 12980
rect 15016 12928 15068 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 15752 12928 15804 12980
rect 16764 12928 16816 12980
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 18696 12971 18748 12980
rect 18696 12937 18705 12971
rect 18705 12937 18739 12971
rect 18739 12937 18748 12971
rect 18696 12928 18748 12937
rect 20076 12928 20128 12980
rect 20168 12928 20220 12980
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 11980 12792 12032 12844
rect 10784 12724 10836 12776
rect 10968 12724 11020 12776
rect 15844 12860 15896 12912
rect 23388 12928 23440 12980
rect 24768 12928 24820 12980
rect 25044 12928 25096 12980
rect 26240 12928 26292 12980
rect 26424 12971 26476 12980
rect 26424 12937 26433 12971
rect 26433 12937 26467 12971
rect 26467 12937 26476 12971
rect 26424 12928 26476 12937
rect 26792 12928 26844 12980
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 15016 12767 15068 12776
rect 10048 12656 10100 12708
rect 13452 12656 13504 12708
rect 11888 12588 11940 12640
rect 12348 12588 12400 12640
rect 13084 12588 13136 12640
rect 13360 12588 13412 12640
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 17224 12724 17276 12776
rect 19156 12724 19208 12776
rect 22192 12792 22244 12844
rect 22744 12792 22796 12844
rect 23020 12792 23072 12844
rect 19800 12724 19852 12776
rect 21456 12767 21508 12776
rect 21456 12733 21465 12767
rect 21465 12733 21499 12767
rect 21499 12733 21508 12767
rect 21456 12724 21508 12733
rect 22100 12724 22152 12776
rect 25688 12792 25740 12844
rect 31392 12928 31444 12980
rect 25412 12767 25464 12776
rect 25412 12733 25421 12767
rect 25421 12733 25455 12767
rect 25455 12733 25464 12767
rect 25412 12724 25464 12733
rect 26148 12724 26200 12776
rect 22376 12656 22428 12708
rect 24032 12699 24084 12708
rect 24032 12665 24041 12699
rect 24041 12665 24075 12699
rect 24075 12665 24084 12699
rect 24032 12656 24084 12665
rect 25596 12656 25648 12708
rect 23756 12588 23808 12640
rect 27436 12588 27488 12640
rect 27712 12656 27764 12708
rect 28816 12860 28868 12912
rect 32312 12928 32364 12980
rect 32496 12971 32548 12980
rect 32496 12937 32505 12971
rect 32505 12937 32539 12971
rect 32539 12937 32548 12971
rect 32496 12928 32548 12937
rect 33508 12971 33560 12980
rect 33508 12937 33517 12971
rect 33517 12937 33551 12971
rect 33551 12937 33560 12971
rect 33508 12928 33560 12937
rect 29000 12792 29052 12844
rect 31760 12860 31812 12912
rect 32036 12724 32088 12776
rect 33692 12835 33744 12844
rect 33692 12801 33701 12835
rect 33701 12801 33735 12835
rect 33735 12801 33744 12835
rect 33692 12792 33744 12801
rect 36544 12928 36596 12980
rect 36636 12928 36688 12980
rect 37740 12928 37792 12980
rect 38844 12928 38896 12980
rect 41604 12928 41656 12980
rect 34152 12860 34204 12912
rect 35440 12860 35492 12912
rect 29736 12656 29788 12708
rect 29828 12631 29880 12640
rect 29828 12597 29837 12631
rect 29837 12597 29871 12631
rect 29871 12597 29880 12631
rect 29828 12588 29880 12597
rect 31392 12588 31444 12640
rect 36728 12792 36780 12844
rect 37832 12792 37884 12844
rect 35348 12724 35400 12776
rect 38384 12656 38436 12708
rect 34428 12588 34480 12640
rect 36268 12588 36320 12640
rect 39856 12724 39908 12776
rect 40224 12835 40276 12844
rect 40224 12801 40233 12835
rect 40233 12801 40267 12835
rect 40267 12801 40276 12835
rect 40224 12792 40276 12801
rect 41696 12860 41748 12912
rect 43812 12928 43864 12980
rect 43996 12971 44048 12980
rect 43996 12937 44005 12971
rect 44005 12937 44039 12971
rect 44039 12937 44048 12971
rect 43996 12928 44048 12937
rect 42248 12860 42300 12912
rect 43720 12860 43772 12912
rect 48964 12928 49016 12980
rect 54300 12928 54352 12980
rect 54392 12928 54444 12980
rect 57428 12928 57480 12980
rect 42708 12792 42760 12844
rect 53472 12860 53524 12912
rect 47860 12792 47912 12844
rect 48044 12835 48096 12844
rect 48044 12801 48078 12835
rect 48078 12801 48096 12835
rect 50528 12835 50580 12844
rect 48044 12792 48096 12801
rect 41788 12588 41840 12640
rect 44272 12724 44324 12776
rect 45560 12767 45612 12776
rect 45560 12733 45569 12767
rect 45569 12733 45603 12767
rect 45603 12733 45612 12767
rect 45560 12724 45612 12733
rect 47216 12724 47268 12776
rect 50528 12801 50537 12835
rect 50537 12801 50571 12835
rect 50571 12801 50580 12835
rect 50528 12792 50580 12801
rect 51172 12792 51224 12844
rect 53196 12792 53248 12844
rect 50804 12724 50856 12776
rect 52368 12767 52420 12776
rect 52368 12733 52377 12767
rect 52377 12733 52411 12767
rect 52411 12733 52420 12767
rect 52368 12724 52420 12733
rect 53656 12792 53708 12844
rect 55680 12860 55732 12912
rect 54116 12792 54168 12844
rect 54760 12792 54812 12844
rect 56968 12860 57020 12912
rect 61476 12928 61528 12980
rect 63868 12971 63920 12980
rect 63868 12937 63877 12971
rect 63877 12937 63911 12971
rect 63911 12937 63920 12971
rect 63868 12928 63920 12937
rect 65432 12971 65484 12980
rect 46940 12699 46992 12708
rect 46940 12665 46949 12699
rect 46949 12665 46983 12699
rect 46983 12665 46992 12699
rect 46940 12656 46992 12665
rect 42892 12588 42944 12640
rect 49608 12656 49660 12708
rect 53012 12656 53064 12708
rect 54024 12656 54076 12708
rect 49148 12631 49200 12640
rect 49148 12597 49157 12631
rect 49157 12597 49191 12631
rect 49191 12597 49200 12631
rect 49148 12588 49200 12597
rect 50896 12588 50948 12640
rect 51632 12588 51684 12640
rect 54300 12588 54352 12640
rect 54392 12588 54444 12640
rect 56048 12792 56100 12844
rect 56876 12792 56928 12844
rect 58256 12835 58308 12844
rect 55680 12724 55732 12776
rect 58256 12801 58265 12835
rect 58265 12801 58299 12835
rect 58299 12801 58308 12835
rect 58256 12792 58308 12801
rect 60556 12835 60608 12844
rect 60556 12801 60574 12835
rect 60574 12801 60608 12835
rect 60832 12835 60884 12844
rect 60556 12792 60608 12801
rect 60832 12801 60841 12835
rect 60841 12801 60875 12835
rect 60875 12801 60884 12835
rect 60832 12792 60884 12801
rect 63408 12860 63460 12912
rect 65432 12937 65441 12971
rect 65441 12937 65475 12971
rect 65475 12937 65484 12971
rect 65432 12928 65484 12937
rect 66076 12971 66128 12980
rect 66076 12937 66085 12971
rect 66085 12937 66119 12971
rect 66119 12937 66128 12971
rect 66076 12928 66128 12937
rect 66996 12971 67048 12980
rect 66996 12937 67005 12971
rect 67005 12937 67039 12971
rect 67039 12937 67048 12971
rect 66996 12928 67048 12937
rect 67548 12928 67600 12980
rect 61384 12792 61436 12844
rect 58808 12724 58860 12776
rect 59176 12724 59228 12776
rect 59544 12724 59596 12776
rect 61016 12724 61068 12776
rect 57980 12588 58032 12640
rect 58164 12588 58216 12640
rect 61936 12588 61988 12640
rect 62764 12588 62816 12640
rect 64420 12792 64472 12844
rect 65156 12860 65208 12912
rect 66904 12860 66956 12912
rect 66260 12835 66312 12844
rect 64052 12656 64104 12708
rect 66260 12801 66269 12835
rect 66269 12801 66303 12835
rect 66303 12801 66312 12835
rect 66260 12792 66312 12801
rect 66812 12835 66864 12844
rect 66812 12801 66821 12835
rect 66821 12801 66855 12835
rect 66855 12801 66864 12835
rect 66812 12792 66864 12801
rect 66904 12724 66956 12776
rect 71780 12928 71832 12980
rect 72516 12928 72568 12980
rect 73620 12928 73672 12980
rect 75276 12928 75328 12980
rect 76380 12928 76432 12980
rect 76656 12928 76708 12980
rect 77208 12928 77260 12980
rect 77392 12928 77444 12980
rect 77760 12928 77812 12980
rect 78772 12971 78824 12980
rect 78772 12937 78781 12971
rect 78781 12937 78815 12971
rect 78815 12937 78824 12971
rect 78772 12928 78824 12937
rect 79508 12971 79560 12980
rect 79508 12937 79517 12971
rect 79517 12937 79551 12971
rect 79551 12937 79560 12971
rect 79508 12928 79560 12937
rect 80244 12928 80296 12980
rect 77576 12860 77628 12912
rect 82452 12928 82504 12980
rect 83556 12928 83608 12980
rect 84016 12928 84068 12980
rect 86592 12928 86644 12980
rect 69480 12835 69532 12844
rect 69480 12801 69498 12835
rect 69498 12801 69532 12835
rect 69480 12792 69532 12801
rect 72332 12792 72384 12844
rect 69940 12724 69992 12776
rect 73068 12792 73120 12844
rect 74632 12792 74684 12844
rect 74816 12835 74868 12844
rect 74816 12801 74825 12835
rect 74825 12801 74859 12835
rect 74859 12801 74868 12835
rect 74816 12792 74868 12801
rect 74172 12724 74224 12776
rect 75000 12724 75052 12776
rect 66444 12656 66496 12708
rect 67640 12588 67692 12640
rect 73344 12656 73396 12708
rect 74632 12656 74684 12708
rect 76656 12724 76708 12776
rect 76840 12792 76892 12844
rect 77392 12792 77444 12844
rect 87328 12860 87380 12912
rect 87420 12860 87472 12912
rect 77300 12724 77352 12776
rect 75736 12656 75788 12708
rect 78956 12835 79008 12844
rect 78956 12801 78965 12835
rect 78965 12801 78999 12835
rect 78999 12801 79008 12835
rect 78956 12792 79008 12801
rect 81348 12835 81400 12844
rect 81348 12801 81382 12835
rect 81382 12801 81400 12835
rect 81348 12792 81400 12801
rect 83188 12835 83240 12844
rect 83188 12801 83197 12835
rect 83197 12801 83231 12835
rect 83231 12801 83240 12835
rect 83188 12792 83240 12801
rect 84108 12835 84160 12844
rect 84108 12801 84117 12835
rect 84117 12801 84151 12835
rect 84151 12801 84160 12835
rect 84108 12792 84160 12801
rect 84476 12792 84528 12844
rect 87880 12835 87932 12844
rect 87880 12801 87889 12835
rect 87889 12801 87923 12835
rect 87923 12801 87932 12835
rect 87880 12792 87932 12801
rect 88156 12792 88208 12844
rect 89444 12860 89496 12912
rect 92388 12928 92440 12980
rect 94320 12928 94372 12980
rect 96804 12928 96856 12980
rect 74264 12588 74316 12640
rect 75644 12588 75696 12640
rect 77484 12588 77536 12640
rect 80244 12588 80296 12640
rect 82084 12724 82136 12776
rect 85396 12724 85448 12776
rect 85488 12767 85540 12776
rect 85488 12733 85497 12767
rect 85497 12733 85531 12767
rect 85531 12733 85540 12767
rect 85488 12724 85540 12733
rect 80520 12699 80572 12708
rect 80520 12665 80529 12699
rect 80529 12665 80563 12699
rect 80563 12665 80572 12699
rect 80520 12656 80572 12665
rect 82452 12631 82504 12640
rect 82452 12597 82461 12631
rect 82461 12597 82495 12631
rect 82495 12597 82504 12631
rect 82452 12588 82504 12597
rect 84660 12588 84712 12640
rect 86776 12588 86828 12640
rect 88432 12724 88484 12776
rect 89352 12792 89404 12844
rect 89812 12724 89864 12776
rect 91652 12860 91704 12912
rect 91376 12792 91428 12844
rect 93400 12835 93452 12844
rect 93400 12801 93409 12835
rect 93409 12801 93443 12835
rect 93443 12801 93452 12835
rect 95332 12860 95384 12912
rect 95976 12860 96028 12912
rect 97632 12928 97684 12980
rect 98552 12928 98604 12980
rect 100024 12928 100076 12980
rect 100116 12928 100168 12980
rect 101772 12928 101824 12980
rect 102600 12928 102652 12980
rect 103980 12928 104032 12980
rect 104808 12928 104860 12980
rect 107016 12928 107068 12980
rect 107292 12928 107344 12980
rect 108396 12928 108448 12980
rect 112260 12928 112312 12980
rect 113640 12971 113692 12980
rect 113640 12937 113649 12971
rect 113649 12937 113683 12971
rect 113683 12937 113692 12971
rect 113640 12928 113692 12937
rect 93400 12792 93452 12801
rect 95516 12792 95568 12844
rect 98460 12860 98512 12912
rect 98000 12835 98052 12844
rect 87972 12656 88024 12708
rect 94228 12724 94280 12776
rect 90548 12656 90600 12708
rect 94320 12656 94372 12708
rect 88892 12588 88944 12640
rect 89536 12588 89588 12640
rect 92388 12588 92440 12640
rect 93216 12631 93268 12640
rect 93216 12597 93225 12631
rect 93225 12597 93259 12631
rect 93259 12597 93268 12631
rect 93216 12588 93268 12597
rect 93400 12588 93452 12640
rect 95240 12724 95292 12776
rect 98000 12801 98009 12835
rect 98009 12801 98043 12835
rect 98043 12801 98052 12835
rect 98000 12792 98052 12801
rect 100392 12860 100444 12912
rect 100116 12835 100168 12844
rect 100116 12801 100125 12835
rect 100125 12801 100159 12835
rect 100159 12801 100168 12835
rect 100116 12792 100168 12801
rect 101312 12792 101364 12844
rect 103888 12860 103940 12912
rect 104072 12860 104124 12912
rect 99380 12724 99432 12776
rect 100208 12724 100260 12776
rect 103612 12724 103664 12776
rect 103888 12767 103940 12776
rect 103888 12733 103897 12767
rect 103897 12733 103931 12767
rect 103931 12733 103940 12767
rect 103888 12724 103940 12733
rect 104900 12792 104952 12844
rect 109408 12860 109460 12912
rect 113272 12860 113324 12912
rect 106924 12792 106976 12844
rect 108120 12792 108172 12844
rect 105728 12724 105780 12776
rect 107016 12767 107068 12776
rect 107016 12733 107025 12767
rect 107025 12733 107059 12767
rect 107059 12733 107068 12767
rect 107016 12724 107068 12733
rect 109040 12835 109092 12844
rect 109040 12801 109049 12835
rect 109049 12801 109083 12835
rect 109083 12801 109092 12835
rect 109040 12792 109092 12801
rect 94688 12656 94740 12708
rect 94872 12631 94924 12640
rect 94872 12597 94881 12631
rect 94881 12597 94915 12631
rect 94915 12597 94924 12631
rect 94872 12588 94924 12597
rect 96896 12656 96948 12708
rect 96988 12656 97040 12708
rect 98000 12588 98052 12640
rect 99288 12631 99340 12640
rect 99288 12597 99297 12631
rect 99297 12597 99331 12631
rect 99331 12597 99340 12631
rect 99288 12588 99340 12597
rect 99564 12656 99616 12708
rect 100668 12656 100720 12708
rect 108948 12656 109000 12708
rect 112444 12724 112496 12776
rect 117688 12928 117740 12980
rect 117780 12928 117832 12980
rect 119712 12928 119764 12980
rect 120080 12928 120132 12980
rect 121092 12928 121144 12980
rect 120632 12860 120684 12912
rect 115756 12792 115808 12844
rect 115848 12792 115900 12844
rect 116584 12835 116636 12844
rect 116584 12801 116593 12835
rect 116593 12801 116627 12835
rect 116627 12801 116636 12835
rect 116584 12792 116636 12801
rect 113548 12724 113600 12776
rect 114744 12767 114796 12776
rect 114744 12733 114753 12767
rect 114753 12733 114787 12767
rect 114787 12733 114796 12767
rect 114744 12724 114796 12733
rect 110328 12656 110380 12708
rect 114468 12656 114520 12708
rect 117964 12699 118016 12708
rect 103796 12588 103848 12640
rect 104808 12588 104860 12640
rect 106280 12588 106332 12640
rect 107660 12588 107712 12640
rect 109132 12588 109184 12640
rect 109408 12588 109460 12640
rect 110420 12631 110472 12640
rect 110420 12597 110429 12631
rect 110429 12597 110463 12631
rect 110463 12597 110472 12631
rect 110420 12588 110472 12597
rect 110972 12631 111024 12640
rect 110972 12597 110981 12631
rect 110981 12597 111015 12631
rect 111015 12597 111024 12631
rect 110972 12588 111024 12597
rect 111340 12588 111392 12640
rect 114560 12588 114612 12640
rect 116124 12631 116176 12640
rect 116124 12597 116133 12631
rect 116133 12597 116167 12631
rect 116167 12597 116176 12631
rect 116124 12588 116176 12597
rect 117964 12665 117973 12699
rect 117973 12665 118007 12699
rect 118007 12665 118016 12699
rect 117964 12656 118016 12665
rect 118792 12792 118844 12844
rect 119252 12792 119304 12844
rect 120172 12835 120224 12844
rect 120172 12801 120181 12835
rect 120181 12801 120215 12835
rect 120215 12801 120224 12835
rect 120172 12792 120224 12801
rect 121460 12792 121512 12844
rect 123208 12928 123260 12980
rect 123300 12928 123352 12980
rect 125324 12928 125376 12980
rect 126888 12928 126940 12980
rect 128268 12928 128320 12980
rect 129556 12971 129608 12980
rect 129556 12937 129565 12971
rect 129565 12937 129599 12971
rect 129599 12937 129608 12971
rect 129556 12928 129608 12937
rect 129740 12928 129792 12980
rect 130476 12928 130528 12980
rect 123392 12860 123444 12912
rect 125968 12860 126020 12912
rect 124312 12835 124364 12844
rect 124312 12801 124321 12835
rect 124321 12801 124355 12835
rect 124355 12801 124364 12835
rect 124312 12792 124364 12801
rect 126980 12860 127032 12912
rect 127348 12860 127400 12912
rect 127440 12860 127492 12912
rect 130016 12860 130068 12912
rect 131212 12928 131264 12980
rect 131856 12971 131908 12980
rect 131856 12937 131865 12971
rect 131865 12937 131899 12971
rect 131899 12937 131908 12971
rect 131856 12928 131908 12937
rect 131948 12928 132000 12980
rect 133604 12928 133656 12980
rect 133788 12928 133840 12980
rect 134892 12928 134944 12980
rect 136548 12928 136600 12980
rect 137928 12971 137980 12980
rect 137928 12937 137937 12971
rect 137937 12937 137971 12971
rect 137971 12937 137980 12971
rect 137928 12928 137980 12937
rect 139492 12928 139544 12980
rect 140596 12928 140648 12980
rect 142160 12928 142212 12980
rect 122012 12724 122064 12776
rect 128820 12792 128872 12844
rect 129004 12835 129056 12844
rect 129004 12801 129013 12835
rect 129013 12801 129047 12835
rect 129047 12801 129056 12835
rect 129004 12792 129056 12801
rect 126888 12767 126940 12776
rect 126888 12733 126897 12767
rect 126897 12733 126931 12767
rect 126931 12733 126940 12767
rect 126888 12724 126940 12733
rect 127992 12724 128044 12776
rect 129924 12792 129976 12844
rect 130476 12835 130528 12844
rect 130476 12801 130485 12835
rect 130485 12801 130519 12835
rect 130519 12801 130528 12835
rect 130476 12792 130528 12801
rect 133144 12860 133196 12912
rect 138572 12860 138624 12912
rect 146300 12928 146352 12980
rect 120172 12656 120224 12708
rect 130568 12724 130620 12776
rect 134156 12792 134208 12844
rect 134340 12835 134392 12844
rect 134340 12801 134349 12835
rect 134349 12801 134383 12835
rect 134383 12801 134392 12835
rect 134340 12792 134392 12801
rect 136640 12835 136692 12844
rect 132776 12767 132828 12776
rect 132776 12733 132785 12767
rect 132785 12733 132819 12767
rect 132819 12733 132828 12767
rect 132776 12724 132828 12733
rect 133052 12767 133104 12776
rect 133052 12733 133061 12767
rect 133061 12733 133095 12767
rect 133095 12733 133104 12767
rect 133052 12724 133104 12733
rect 136640 12801 136649 12835
rect 136649 12801 136683 12835
rect 136683 12801 136692 12835
rect 136640 12792 136692 12801
rect 137744 12835 137796 12844
rect 137744 12801 137753 12835
rect 137753 12801 137787 12835
rect 137787 12801 137796 12835
rect 137744 12792 137796 12801
rect 143356 12860 143408 12912
rect 135720 12724 135772 12776
rect 136180 12724 136232 12776
rect 139584 12792 139636 12844
rect 141516 12792 141568 12844
rect 142528 12792 142580 12844
rect 142712 12835 142764 12844
rect 142712 12801 142721 12835
rect 142721 12801 142755 12835
rect 142755 12801 142764 12835
rect 142712 12792 142764 12801
rect 148508 12860 148560 12912
rect 148784 12860 148836 12912
rect 150900 12928 150952 12980
rect 152004 12928 152056 12980
rect 152924 12928 152976 12980
rect 153476 12928 153528 12980
rect 156144 12971 156196 12980
rect 156144 12937 156153 12971
rect 156153 12937 156187 12971
rect 156187 12937 156196 12971
rect 156144 12928 156196 12937
rect 156788 12928 156840 12980
rect 158076 12971 158128 12980
rect 158076 12937 158085 12971
rect 158085 12937 158119 12971
rect 158119 12937 158128 12971
rect 158076 12928 158128 12937
rect 151360 12860 151412 12912
rect 147496 12835 147548 12844
rect 147496 12801 147505 12835
rect 147505 12801 147539 12835
rect 147539 12801 147548 12835
rect 147496 12792 147548 12801
rect 148876 12792 148928 12844
rect 149520 12792 149572 12844
rect 149704 12792 149756 12844
rect 152464 12860 152516 12912
rect 118148 12588 118200 12640
rect 119160 12631 119212 12640
rect 119160 12597 119169 12631
rect 119169 12597 119203 12631
rect 119203 12597 119212 12631
rect 119160 12588 119212 12597
rect 119252 12588 119304 12640
rect 122380 12588 122432 12640
rect 122472 12588 122524 12640
rect 125232 12588 125284 12640
rect 125968 12588 126020 12640
rect 126704 12588 126756 12640
rect 142344 12656 142396 12708
rect 143908 12656 143960 12708
rect 129924 12588 129976 12640
rect 135352 12588 135404 12640
rect 142620 12588 142672 12640
rect 145840 12724 145892 12776
rect 149152 12656 149204 12708
rect 150072 12699 150124 12708
rect 144736 12588 144788 12640
rect 145564 12588 145616 12640
rect 147036 12588 147088 12640
rect 150072 12665 150081 12699
rect 150081 12665 150115 12699
rect 150115 12665 150124 12699
rect 150072 12656 150124 12665
rect 150808 12699 150860 12708
rect 150808 12665 150817 12699
rect 150817 12665 150851 12699
rect 150851 12665 150860 12699
rect 150808 12656 150860 12665
rect 150348 12588 150400 12640
rect 153384 12792 153436 12844
rect 153752 12835 153804 12844
rect 155408 12860 155460 12912
rect 155592 12860 155644 12912
rect 153752 12801 153770 12835
rect 153770 12801 153804 12835
rect 153752 12792 153804 12801
rect 154120 12724 154172 12776
rect 156052 12792 156104 12844
rect 156696 12835 156748 12844
rect 156696 12801 156705 12835
rect 156705 12801 156739 12835
rect 156739 12801 156748 12835
rect 156696 12792 156748 12801
rect 152648 12699 152700 12708
rect 152648 12665 152657 12699
rect 152657 12665 152691 12699
rect 152691 12665 152700 12699
rect 152648 12656 152700 12665
rect 152740 12588 152792 12640
rect 154304 12588 154356 12640
rect 158352 12724 158404 12776
rect 158168 12656 158220 12708
rect 20672 12486 20724 12538
rect 20736 12486 20788 12538
rect 20800 12486 20852 12538
rect 20864 12486 20916 12538
rect 20928 12486 20980 12538
rect 60117 12486 60169 12538
rect 60181 12486 60233 12538
rect 60245 12486 60297 12538
rect 60309 12486 60361 12538
rect 60373 12486 60425 12538
rect 99562 12486 99614 12538
rect 99626 12486 99678 12538
rect 99690 12486 99742 12538
rect 99754 12486 99806 12538
rect 99818 12486 99870 12538
rect 139007 12486 139059 12538
rect 139071 12486 139123 12538
rect 139135 12486 139187 12538
rect 139199 12486 139251 12538
rect 139263 12486 139315 12538
rect 10508 12427 10560 12436
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 12072 12384 12124 12436
rect 14004 12384 14056 12436
rect 14096 12384 14148 12436
rect 10048 12248 10100 12300
rect 10968 12248 11020 12300
rect 4436 12180 4488 12232
rect 5724 12180 5776 12232
rect 9864 12223 9916 12232
rect 6828 12112 6880 12164
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11704 12112 11756 12164
rect 19892 12316 19944 12368
rect 20628 12316 20680 12368
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 22836 12384 22888 12436
rect 24492 12384 24544 12436
rect 27252 12427 27304 12436
rect 24400 12316 24452 12368
rect 26148 12316 26200 12368
rect 27252 12393 27261 12427
rect 27261 12393 27295 12427
rect 27295 12393 27304 12427
rect 27252 12384 27304 12393
rect 27804 12384 27856 12436
rect 29460 12384 29512 12436
rect 30656 12427 30708 12436
rect 30656 12393 30665 12427
rect 30665 12393 30699 12427
rect 30699 12393 30708 12427
rect 30656 12384 30708 12393
rect 31300 12384 31352 12436
rect 31668 12384 31720 12436
rect 33876 12384 33928 12436
rect 35164 12427 35216 12436
rect 35164 12393 35173 12427
rect 35173 12393 35207 12427
rect 35207 12393 35216 12427
rect 35164 12384 35216 12393
rect 36084 12384 36136 12436
rect 37188 12384 37240 12436
rect 38292 12384 38344 12436
rect 39948 12384 40000 12436
rect 32036 12291 32088 12300
rect 13176 12180 13228 12232
rect 13544 12180 13596 12232
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 16212 12180 16264 12232
rect 19432 12180 19484 12232
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 21456 12180 21508 12232
rect 24584 12223 24636 12232
rect 14464 12112 14516 12164
rect 15660 12112 15712 12164
rect 16304 12112 16356 12164
rect 4160 12044 4212 12096
rect 9588 12044 9640 12096
rect 14924 12044 14976 12096
rect 16120 12044 16172 12096
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 17224 12044 17276 12096
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 27344 12180 27396 12232
rect 28172 12223 28224 12232
rect 24860 12155 24912 12164
rect 24860 12121 24894 12155
rect 24894 12121 24912 12155
rect 26608 12155 26660 12164
rect 24860 12112 24912 12121
rect 18880 12044 18932 12096
rect 19248 12044 19300 12096
rect 20720 12044 20772 12096
rect 24124 12044 24176 12096
rect 25780 12044 25832 12096
rect 26608 12121 26617 12155
rect 26617 12121 26651 12155
rect 26651 12121 26660 12155
rect 26608 12112 26660 12121
rect 26976 12112 27028 12164
rect 28172 12189 28181 12223
rect 28181 12189 28215 12223
rect 28215 12189 28224 12223
rect 28172 12180 28224 12189
rect 28356 12180 28408 12232
rect 32036 12257 32045 12291
rect 32045 12257 32079 12291
rect 32079 12257 32088 12291
rect 32036 12248 32088 12257
rect 38108 12316 38160 12368
rect 38200 12316 38252 12368
rect 41696 12384 41748 12436
rect 44272 12384 44324 12436
rect 45560 12384 45612 12436
rect 47032 12384 47084 12436
rect 48780 12384 48832 12436
rect 42156 12316 42208 12368
rect 43536 12316 43588 12368
rect 43904 12316 43956 12368
rect 35348 12223 35400 12232
rect 28540 12112 28592 12164
rect 29184 12087 29236 12096
rect 29184 12053 29193 12087
rect 29193 12053 29227 12087
rect 29227 12053 29236 12087
rect 29184 12044 29236 12053
rect 30656 12044 30708 12096
rect 30932 12044 30984 12096
rect 35348 12189 35357 12223
rect 35357 12189 35391 12223
rect 35391 12189 35400 12223
rect 35348 12180 35400 12189
rect 36176 12223 36228 12232
rect 36176 12189 36185 12223
rect 36185 12189 36219 12223
rect 36219 12189 36228 12223
rect 36176 12180 36228 12189
rect 36360 12180 36412 12232
rect 38200 12180 38252 12232
rect 38384 12223 38436 12232
rect 38384 12189 38393 12223
rect 38393 12189 38427 12223
rect 38427 12189 38436 12223
rect 38384 12180 38436 12189
rect 39212 12223 39264 12232
rect 39212 12189 39221 12223
rect 39221 12189 39255 12223
rect 39255 12189 39264 12223
rect 39212 12180 39264 12189
rect 40224 12223 40276 12232
rect 40224 12189 40233 12223
rect 40233 12189 40267 12223
rect 40267 12189 40276 12223
rect 40224 12180 40276 12189
rect 41236 12248 41288 12300
rect 41420 12180 41472 12232
rect 42064 12223 42116 12232
rect 42064 12189 42073 12223
rect 42073 12189 42107 12223
rect 42107 12189 42116 12223
rect 42064 12180 42116 12189
rect 43996 12248 44048 12300
rect 51448 12316 51500 12368
rect 51080 12248 51132 12300
rect 34336 12112 34388 12164
rect 37648 12112 37700 12164
rect 38108 12112 38160 12164
rect 39856 12112 39908 12164
rect 40316 12112 40368 12164
rect 45008 12180 45060 12232
rect 45468 12223 45520 12232
rect 45468 12189 45477 12223
rect 45477 12189 45511 12223
rect 45511 12189 45520 12223
rect 45468 12180 45520 12189
rect 45928 12223 45980 12232
rect 45928 12189 45937 12223
rect 45937 12189 45971 12223
rect 45971 12189 45980 12223
rect 45928 12180 45980 12189
rect 49700 12180 49752 12232
rect 49792 12180 49844 12232
rect 50252 12180 50304 12232
rect 51632 12223 51684 12232
rect 51632 12189 51641 12223
rect 51641 12189 51675 12223
rect 51675 12189 51684 12223
rect 51632 12180 51684 12189
rect 51724 12180 51776 12232
rect 52368 12384 52420 12436
rect 55588 12384 55640 12436
rect 56140 12384 56192 12436
rect 56784 12384 56836 12436
rect 57888 12384 57940 12436
rect 54300 12316 54352 12368
rect 57244 12316 57296 12368
rect 58256 12384 58308 12436
rect 63224 12427 63276 12436
rect 63224 12393 63233 12427
rect 63233 12393 63267 12427
rect 63267 12393 63276 12427
rect 63224 12384 63276 12393
rect 63776 12384 63828 12436
rect 64788 12384 64840 12436
rect 68652 12384 68704 12436
rect 69756 12384 69808 12436
rect 71780 12384 71832 12436
rect 73068 12384 73120 12436
rect 75368 12427 75420 12436
rect 61016 12316 61068 12368
rect 66168 12316 66220 12368
rect 69112 12316 69164 12368
rect 69940 12316 69992 12368
rect 56692 12248 56744 12300
rect 57152 12248 57204 12300
rect 67916 12248 67968 12300
rect 54300 12180 54352 12232
rect 33692 12044 33744 12096
rect 33968 12044 34020 12096
rect 34888 12044 34940 12096
rect 48780 12112 48832 12164
rect 50160 12112 50212 12164
rect 42156 12044 42208 12096
rect 42708 12044 42760 12096
rect 42892 12044 42944 12096
rect 44088 12044 44140 12096
rect 46664 12044 46716 12096
rect 47308 12087 47360 12096
rect 47308 12053 47317 12087
rect 47317 12053 47351 12087
rect 47351 12053 47360 12087
rect 47308 12044 47360 12053
rect 47768 12087 47820 12096
rect 47768 12053 47777 12087
rect 47777 12053 47811 12087
rect 47811 12053 47820 12087
rect 52000 12112 52052 12164
rect 53012 12112 53064 12164
rect 54852 12180 54904 12232
rect 55680 12223 55732 12232
rect 55680 12189 55689 12223
rect 55689 12189 55723 12223
rect 55723 12189 55732 12223
rect 55680 12180 55732 12189
rect 55956 12180 56008 12232
rect 56048 12180 56100 12232
rect 56324 12180 56376 12232
rect 57060 12180 57112 12232
rect 57244 12223 57296 12232
rect 57244 12189 57253 12223
rect 57253 12189 57287 12223
rect 57287 12189 57296 12223
rect 57244 12180 57296 12189
rect 57336 12180 57388 12232
rect 59544 12223 59596 12232
rect 59544 12189 59553 12223
rect 59553 12189 59587 12223
rect 59587 12189 59596 12223
rect 61016 12223 61068 12232
rect 59544 12180 59596 12189
rect 61016 12189 61025 12223
rect 61025 12189 61059 12223
rect 61059 12189 61068 12223
rect 61016 12180 61068 12189
rect 47768 12044 47820 12053
rect 54576 12044 54628 12096
rect 55312 12044 55364 12096
rect 55496 12087 55548 12096
rect 55496 12053 55505 12087
rect 55505 12053 55539 12087
rect 55539 12053 55548 12087
rect 55496 12044 55548 12053
rect 62396 12180 62448 12232
rect 62488 12180 62540 12232
rect 61660 12112 61712 12164
rect 65800 12180 65852 12232
rect 72332 12316 72384 12368
rect 75368 12393 75377 12427
rect 75377 12393 75411 12427
rect 75411 12393 75420 12427
rect 75368 12384 75420 12393
rect 76196 12384 76248 12436
rect 77484 12384 77536 12436
rect 77760 12427 77812 12436
rect 77760 12393 77769 12427
rect 77769 12393 77803 12427
rect 77803 12393 77812 12427
rect 77760 12384 77812 12393
rect 84752 12384 84804 12436
rect 85212 12384 85264 12436
rect 85764 12384 85816 12436
rect 87328 12384 87380 12436
rect 87880 12384 87932 12436
rect 79692 12316 79744 12368
rect 80520 12316 80572 12368
rect 82176 12316 82228 12368
rect 88156 12316 88208 12368
rect 89168 12316 89220 12368
rect 89904 12316 89956 12368
rect 75920 12248 75972 12300
rect 76748 12248 76800 12300
rect 77392 12248 77444 12300
rect 77760 12248 77812 12300
rect 56784 12044 56836 12096
rect 68836 12112 68888 12164
rect 73160 12180 73212 12232
rect 66168 12044 66220 12096
rect 66812 12044 66864 12096
rect 68744 12044 68796 12096
rect 71136 12044 71188 12096
rect 71688 12087 71740 12096
rect 71688 12053 71697 12087
rect 71697 12053 71731 12087
rect 71731 12053 71740 12087
rect 71688 12044 71740 12053
rect 78588 12180 78640 12232
rect 77300 12155 77352 12164
rect 77300 12121 77309 12155
rect 77309 12121 77343 12155
rect 77343 12121 77352 12155
rect 77300 12112 77352 12121
rect 75276 12044 75328 12096
rect 75552 12044 75604 12096
rect 80520 12180 80572 12232
rect 81716 12180 81768 12232
rect 83096 12248 83148 12300
rect 84108 12248 84160 12300
rect 85396 12248 85448 12300
rect 82084 12223 82136 12232
rect 82084 12189 82093 12223
rect 82093 12189 82127 12223
rect 82127 12189 82136 12223
rect 82084 12180 82136 12189
rect 89536 12248 89588 12300
rect 90088 12248 90140 12300
rect 90180 12248 90232 12300
rect 86408 12223 86460 12232
rect 86408 12189 86417 12223
rect 86417 12189 86451 12223
rect 86451 12189 86460 12223
rect 86408 12180 86460 12189
rect 89168 12223 89220 12232
rect 89168 12189 89177 12223
rect 89177 12189 89211 12223
rect 89211 12189 89220 12223
rect 89168 12180 89220 12189
rect 89444 12180 89496 12232
rect 90364 12223 90416 12232
rect 77484 12044 77536 12096
rect 82452 12112 82504 12164
rect 79140 12044 79192 12096
rect 80704 12044 80756 12096
rect 81624 12087 81676 12096
rect 81624 12053 81633 12087
rect 81633 12053 81667 12087
rect 81667 12053 81676 12087
rect 81624 12044 81676 12053
rect 81716 12044 81768 12096
rect 82636 12087 82688 12096
rect 82636 12053 82645 12087
rect 82645 12053 82679 12087
rect 82679 12053 82688 12087
rect 82636 12044 82688 12053
rect 83280 12087 83332 12096
rect 83280 12053 83289 12087
rect 83289 12053 83323 12087
rect 83323 12053 83332 12087
rect 83280 12044 83332 12053
rect 84292 12044 84344 12096
rect 84476 12044 84528 12096
rect 84752 12112 84804 12164
rect 88064 12112 88116 12164
rect 88892 12155 88944 12164
rect 88892 12121 88910 12155
rect 88910 12121 88944 12155
rect 88892 12112 88944 12121
rect 90364 12189 90373 12223
rect 90373 12189 90407 12223
rect 90407 12189 90416 12223
rect 90364 12180 90416 12189
rect 93032 12248 93084 12300
rect 93308 12248 93360 12300
rect 96252 12384 96304 12436
rect 98736 12427 98788 12436
rect 98736 12393 98745 12427
rect 98745 12393 98779 12427
rect 98779 12393 98788 12427
rect 98736 12384 98788 12393
rect 99932 12384 99984 12436
rect 102048 12384 102100 12436
rect 104624 12384 104676 12436
rect 105084 12384 105136 12436
rect 105636 12384 105688 12436
rect 106740 12384 106792 12436
rect 107292 12384 107344 12436
rect 110236 12427 110288 12436
rect 98184 12316 98236 12368
rect 101404 12316 101456 12368
rect 101588 12248 101640 12300
rect 93676 12223 93728 12232
rect 93676 12189 93685 12223
rect 93685 12189 93719 12223
rect 93719 12189 93728 12223
rect 93676 12180 93728 12189
rect 96160 12223 96212 12232
rect 89904 12112 89956 12164
rect 90824 12112 90876 12164
rect 93124 12112 93176 12164
rect 93216 12112 93268 12164
rect 96160 12189 96169 12223
rect 96169 12189 96203 12223
rect 96203 12189 96212 12223
rect 96160 12180 96212 12189
rect 96988 12223 97040 12232
rect 96988 12189 96997 12223
rect 96997 12189 97031 12223
rect 97031 12189 97040 12223
rect 96988 12180 97040 12189
rect 99288 12180 99340 12232
rect 100300 12180 100352 12232
rect 102968 12223 103020 12232
rect 102968 12189 102977 12223
rect 102977 12189 103011 12223
rect 103011 12189 103020 12223
rect 102968 12180 103020 12189
rect 103060 12180 103112 12232
rect 104348 12223 104400 12232
rect 104348 12189 104357 12223
rect 104357 12189 104391 12223
rect 104391 12189 104400 12223
rect 104348 12180 104400 12189
rect 106372 12248 106424 12300
rect 108672 12316 108724 12368
rect 110236 12393 110245 12427
rect 110245 12393 110279 12427
rect 110279 12393 110288 12427
rect 110236 12384 110288 12393
rect 111708 12384 111760 12436
rect 112352 12384 112404 12436
rect 118516 12384 118568 12436
rect 121644 12384 121696 12436
rect 121828 12384 121880 12436
rect 126060 12384 126112 12436
rect 127164 12384 127216 12436
rect 128452 12427 128504 12436
rect 128452 12393 128461 12427
rect 128461 12393 128495 12427
rect 128495 12393 128504 12427
rect 128452 12384 128504 12393
rect 129096 12384 129148 12436
rect 130476 12384 130528 12436
rect 135076 12384 135128 12436
rect 135536 12427 135588 12436
rect 135536 12393 135545 12427
rect 135545 12393 135579 12427
rect 135579 12393 135588 12427
rect 135536 12384 135588 12393
rect 137192 12384 137244 12436
rect 141332 12427 141384 12436
rect 104624 12180 104676 12232
rect 106188 12223 106240 12232
rect 106188 12189 106197 12223
rect 106197 12189 106231 12223
rect 106231 12189 106240 12223
rect 106188 12180 106240 12189
rect 107292 12223 107344 12232
rect 107292 12189 107301 12223
rect 107301 12189 107335 12223
rect 107335 12189 107344 12223
rect 107292 12180 107344 12189
rect 107568 12180 107620 12232
rect 114284 12248 114336 12300
rect 110880 12223 110932 12232
rect 98184 12155 98236 12164
rect 98184 12121 98193 12155
rect 98193 12121 98227 12155
rect 98227 12121 98236 12155
rect 98184 12112 98236 12121
rect 101036 12112 101088 12164
rect 109408 12155 109460 12164
rect 91560 12087 91612 12096
rect 91560 12053 91569 12087
rect 91569 12053 91603 12087
rect 91603 12053 91612 12087
rect 91560 12044 91612 12053
rect 91836 12044 91888 12096
rect 94780 12087 94832 12096
rect 94780 12053 94789 12087
rect 94789 12053 94823 12087
rect 94823 12053 94832 12087
rect 94780 12044 94832 12053
rect 96528 12044 96580 12096
rect 100392 12087 100444 12096
rect 100392 12053 100401 12087
rect 100401 12053 100435 12087
rect 100435 12053 100444 12087
rect 100392 12044 100444 12053
rect 101312 12087 101364 12096
rect 101312 12053 101321 12087
rect 101321 12053 101355 12087
rect 101355 12053 101364 12087
rect 101312 12044 101364 12053
rect 101496 12044 101548 12096
rect 101956 12087 102008 12096
rect 101956 12053 101965 12087
rect 101965 12053 101999 12087
rect 101999 12053 102008 12087
rect 101956 12044 102008 12053
rect 102324 12044 102376 12096
rect 103612 12044 103664 12096
rect 105636 12044 105688 12096
rect 105820 12044 105872 12096
rect 107936 12044 107988 12096
rect 108028 12044 108080 12096
rect 109408 12121 109426 12155
rect 109426 12121 109460 12155
rect 109408 12112 109460 12121
rect 110880 12189 110889 12223
rect 110889 12189 110923 12223
rect 110923 12189 110932 12223
rect 110880 12180 110932 12189
rect 111248 12180 111300 12232
rect 114836 12180 114888 12232
rect 117964 12248 118016 12300
rect 116492 12223 116544 12232
rect 116492 12189 116501 12223
rect 116501 12189 116535 12223
rect 116535 12189 116544 12223
rect 116492 12180 116544 12189
rect 117228 12180 117280 12232
rect 118516 12180 118568 12232
rect 122748 12248 122800 12300
rect 125600 12316 125652 12368
rect 126796 12316 126848 12368
rect 127992 12316 128044 12368
rect 112536 12112 112588 12164
rect 115296 12112 115348 12164
rect 120448 12180 120500 12232
rect 121828 12180 121880 12232
rect 123852 12223 123904 12232
rect 123852 12189 123861 12223
rect 123861 12189 123895 12223
rect 123895 12189 123904 12223
rect 128452 12248 128504 12300
rect 128544 12248 128596 12300
rect 133880 12316 133932 12368
rect 123852 12180 123904 12189
rect 125508 12180 125560 12232
rect 126520 12180 126572 12232
rect 127440 12180 127492 12232
rect 127900 12180 127952 12232
rect 131764 12248 131816 12300
rect 130016 12223 130068 12232
rect 130016 12189 130025 12223
rect 130025 12189 130059 12223
rect 130059 12189 130068 12223
rect 130016 12180 130068 12189
rect 130108 12180 130160 12232
rect 132132 12180 132184 12232
rect 133144 12180 133196 12232
rect 135904 12180 135956 12232
rect 141332 12393 141341 12427
rect 141341 12393 141375 12427
rect 141375 12393 141384 12427
rect 141332 12384 141384 12393
rect 143172 12384 143224 12436
rect 141884 12359 141936 12368
rect 141884 12325 141893 12359
rect 141893 12325 141927 12359
rect 141927 12325 141936 12359
rect 141884 12316 141936 12325
rect 143264 12248 143316 12300
rect 138020 12223 138072 12232
rect 138020 12189 138029 12223
rect 138029 12189 138063 12223
rect 138063 12189 138072 12223
rect 140504 12223 140556 12232
rect 138020 12180 138072 12189
rect 140504 12189 140513 12223
rect 140513 12189 140547 12223
rect 140547 12189 140556 12223
rect 140504 12180 140556 12189
rect 140596 12180 140648 12232
rect 141240 12180 141292 12232
rect 111064 12044 111116 12096
rect 111616 12044 111668 12096
rect 113548 12087 113600 12096
rect 113548 12053 113557 12087
rect 113557 12053 113591 12087
rect 113591 12053 113600 12087
rect 113548 12044 113600 12053
rect 114284 12044 114336 12096
rect 114560 12087 114612 12096
rect 114560 12053 114569 12087
rect 114569 12053 114603 12087
rect 114603 12053 114612 12087
rect 114560 12044 114612 12053
rect 115204 12087 115256 12096
rect 115204 12053 115213 12087
rect 115213 12053 115247 12087
rect 115247 12053 115256 12087
rect 115204 12044 115256 12053
rect 116308 12087 116360 12096
rect 116308 12053 116317 12087
rect 116317 12053 116351 12087
rect 116351 12053 116360 12087
rect 116308 12044 116360 12053
rect 116400 12044 116452 12096
rect 118884 12087 118936 12096
rect 118884 12053 118893 12087
rect 118893 12053 118927 12087
rect 118927 12053 118936 12087
rect 118884 12044 118936 12053
rect 119896 12044 119948 12096
rect 120816 12087 120868 12096
rect 120816 12053 120825 12087
rect 120825 12053 120859 12087
rect 120859 12053 120868 12087
rect 120816 12044 120868 12053
rect 123760 12112 123812 12164
rect 124312 12044 124364 12096
rect 124864 12044 124916 12096
rect 126336 12044 126388 12096
rect 126704 12044 126756 12096
rect 126888 12044 126940 12096
rect 126980 12044 127032 12096
rect 130660 12087 130712 12096
rect 130660 12053 130669 12087
rect 130669 12053 130703 12087
rect 130703 12053 130712 12087
rect 130660 12044 130712 12053
rect 131212 12087 131264 12096
rect 131212 12053 131221 12087
rect 131221 12053 131255 12087
rect 131255 12053 131264 12087
rect 131212 12044 131264 12053
rect 131764 12087 131816 12096
rect 131764 12053 131773 12087
rect 131773 12053 131807 12087
rect 131807 12053 131816 12087
rect 131764 12044 131816 12053
rect 132408 12044 132460 12096
rect 133328 12087 133380 12096
rect 133328 12053 133337 12087
rect 133337 12053 133371 12087
rect 133371 12053 133380 12087
rect 133328 12044 133380 12053
rect 135352 12112 135404 12164
rect 141424 12112 141476 12164
rect 141884 12112 141936 12164
rect 144276 12155 144328 12164
rect 144276 12121 144294 12155
rect 144294 12121 144328 12155
rect 144276 12112 144328 12121
rect 144736 12180 144788 12232
rect 144828 12180 144880 12232
rect 146392 12223 146444 12232
rect 146116 12155 146168 12164
rect 138112 12044 138164 12096
rect 139124 12087 139176 12096
rect 139124 12053 139133 12087
rect 139133 12053 139167 12087
rect 139167 12053 139176 12087
rect 139124 12044 139176 12053
rect 140044 12044 140096 12096
rect 142344 12044 142396 12096
rect 143172 12087 143224 12096
rect 143172 12053 143181 12087
rect 143181 12053 143215 12087
rect 143215 12053 143224 12087
rect 143172 12044 143224 12053
rect 145012 12087 145064 12096
rect 145012 12053 145021 12087
rect 145021 12053 145055 12087
rect 145055 12053 145064 12087
rect 145012 12044 145064 12053
rect 146116 12121 146134 12155
rect 146134 12121 146168 12155
rect 146116 12112 146168 12121
rect 146392 12189 146401 12223
rect 146401 12189 146435 12223
rect 146435 12189 146444 12223
rect 146392 12180 146444 12189
rect 148140 12384 148192 12436
rect 153108 12384 153160 12436
rect 154764 12316 154816 12368
rect 148416 12248 148468 12300
rect 148048 12180 148100 12232
rect 148232 12180 148284 12232
rect 148600 12180 148652 12232
rect 150256 12180 150308 12232
rect 151360 12223 151412 12232
rect 151360 12189 151369 12223
rect 151369 12189 151403 12223
rect 151403 12189 151412 12223
rect 151360 12180 151412 12189
rect 152648 12223 152700 12232
rect 147680 12112 147732 12164
rect 150532 12112 150584 12164
rect 151084 12155 151136 12164
rect 151084 12121 151102 12155
rect 151102 12121 151136 12155
rect 152648 12189 152657 12223
rect 152657 12189 152691 12223
rect 152691 12189 152700 12223
rect 152648 12180 152700 12189
rect 153016 12180 153068 12232
rect 155868 12248 155920 12300
rect 151084 12112 151136 12121
rect 147588 12087 147640 12096
rect 147588 12053 147597 12087
rect 147597 12053 147631 12087
rect 147631 12053 147640 12087
rect 147588 12044 147640 12053
rect 148324 12087 148376 12096
rect 148324 12053 148333 12087
rect 148333 12053 148367 12087
rect 148367 12053 148376 12087
rect 148324 12044 148376 12053
rect 148416 12044 148468 12096
rect 149244 12044 149296 12096
rect 151912 12044 151964 12096
rect 153752 12112 153804 12164
rect 154672 12180 154724 12232
rect 155224 12180 155276 12232
rect 155500 12180 155552 12232
rect 159180 12180 159232 12232
rect 157064 12044 157116 12096
rect 40394 11942 40446 11994
rect 40458 11942 40510 11994
rect 40522 11942 40574 11994
rect 40586 11942 40638 11994
rect 40650 11942 40702 11994
rect 79839 11942 79891 11994
rect 79903 11942 79955 11994
rect 79967 11942 80019 11994
rect 80031 11942 80083 11994
rect 80095 11942 80147 11994
rect 119284 11942 119336 11994
rect 119348 11942 119400 11994
rect 119412 11942 119464 11994
rect 119476 11942 119528 11994
rect 119540 11942 119592 11994
rect 158729 11942 158781 11994
rect 158793 11942 158845 11994
rect 158857 11942 158909 11994
rect 158921 11942 158973 11994
rect 158985 11942 159037 11994
rect 13176 11840 13228 11892
rect 4068 11747 4120 11756
rect 4068 11713 4102 11747
rect 4102 11713 4120 11747
rect 8392 11747 8444 11756
rect 4068 11704 4120 11713
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 11244 11704 11296 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 12532 11704 12584 11756
rect 13360 11704 13412 11756
rect 14280 11840 14332 11892
rect 14924 11772 14976 11824
rect 15568 11772 15620 11824
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 14556 11704 14608 11756
rect 15200 11704 15252 11756
rect 15476 11704 15528 11756
rect 16120 11704 16172 11756
rect 17224 11704 17276 11756
rect 20168 11840 20220 11892
rect 20536 11840 20588 11892
rect 21640 11840 21692 11892
rect 27620 11840 27672 11892
rect 27988 11840 28040 11892
rect 31116 11840 31168 11892
rect 32312 11840 32364 11892
rect 32864 11883 32916 11892
rect 32864 11849 32873 11883
rect 32873 11849 32907 11883
rect 32907 11849 32916 11883
rect 32864 11840 32916 11849
rect 36360 11883 36412 11892
rect 36360 11849 36369 11883
rect 36369 11849 36403 11883
rect 36403 11849 36412 11883
rect 36360 11840 36412 11849
rect 37648 11840 37700 11892
rect 39304 11840 39356 11892
rect 39488 11840 39540 11892
rect 40224 11840 40276 11892
rect 41696 11840 41748 11892
rect 43260 11840 43312 11892
rect 19800 11772 19852 11824
rect 21916 11772 21968 11824
rect 6092 11568 6144 11620
rect 5540 11500 5592 11552
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 10324 11568 10376 11620
rect 12624 11636 12676 11688
rect 12900 11636 12952 11688
rect 17040 11636 17092 11688
rect 18144 11636 18196 11688
rect 19248 11636 19300 11688
rect 21088 11704 21140 11756
rect 29184 11772 29236 11824
rect 29552 11772 29604 11824
rect 30472 11772 30524 11824
rect 35900 11772 35952 11824
rect 40040 11772 40092 11824
rect 22192 11704 22244 11756
rect 24124 11747 24176 11756
rect 7748 11500 7800 11509
rect 10048 11500 10100 11552
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 18604 11568 18656 11620
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 15936 11500 15988 11552
rect 19340 11500 19392 11552
rect 20168 11543 20220 11552
rect 20168 11509 20177 11543
rect 20177 11509 20211 11543
rect 20211 11509 20220 11543
rect 20168 11500 20220 11509
rect 20260 11500 20312 11552
rect 22100 11500 22152 11552
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 24952 11704 25004 11756
rect 27712 11704 27764 11756
rect 28816 11704 28868 11756
rect 23756 11636 23808 11688
rect 26240 11636 26292 11688
rect 26608 11636 26660 11688
rect 25964 11568 26016 11620
rect 22284 11500 22336 11509
rect 27068 11500 27120 11552
rect 30196 11704 30248 11756
rect 31668 11704 31720 11756
rect 32036 11704 32088 11756
rect 34060 11704 34112 11756
rect 29000 11636 29052 11688
rect 29644 11679 29696 11688
rect 29644 11645 29653 11679
rect 29653 11645 29687 11679
rect 29687 11645 29696 11679
rect 29644 11636 29696 11645
rect 30840 11636 30892 11688
rect 39120 11704 39172 11756
rect 41512 11704 41564 11756
rect 41972 11704 42024 11756
rect 43628 11772 43680 11824
rect 43904 11772 43956 11824
rect 42156 11704 42208 11756
rect 42800 11704 42852 11756
rect 44180 11747 44232 11756
rect 44180 11713 44189 11747
rect 44189 11713 44223 11747
rect 44223 11713 44232 11747
rect 44180 11704 44232 11713
rect 45652 11747 45704 11756
rect 45652 11713 45661 11747
rect 45661 11713 45695 11747
rect 45695 11713 45704 11747
rect 45652 11704 45704 11713
rect 46388 11772 46440 11824
rect 46940 11840 46992 11892
rect 48136 11840 48188 11892
rect 50988 11840 51040 11892
rect 48228 11772 48280 11824
rect 49516 11772 49568 11824
rect 52368 11840 52420 11892
rect 52828 11840 52880 11892
rect 54300 11883 54352 11892
rect 54300 11849 54309 11883
rect 54309 11849 54343 11883
rect 54343 11849 54352 11883
rect 54300 11840 54352 11849
rect 54392 11840 54444 11892
rect 56048 11840 56100 11892
rect 47676 11704 47728 11756
rect 49148 11704 49200 11756
rect 49332 11747 49384 11756
rect 49332 11713 49341 11747
rect 49341 11713 49375 11747
rect 49375 11713 49384 11747
rect 49332 11704 49384 11713
rect 50068 11747 50120 11756
rect 50068 11713 50102 11747
rect 50102 11713 50120 11747
rect 51908 11747 51960 11756
rect 50068 11704 50120 11713
rect 51908 11713 51917 11747
rect 51917 11713 51951 11747
rect 51951 11713 51960 11747
rect 51908 11704 51960 11713
rect 52460 11704 52512 11756
rect 53564 11747 53616 11756
rect 53564 11713 53573 11747
rect 53573 11713 53607 11747
rect 53607 11713 53616 11747
rect 53564 11704 53616 11713
rect 55220 11772 55272 11824
rect 55312 11772 55364 11824
rect 57244 11840 57296 11892
rect 58624 11840 58676 11892
rect 59084 11840 59136 11892
rect 59452 11883 59504 11892
rect 59452 11849 59461 11883
rect 59461 11849 59495 11883
rect 59495 11849 59504 11883
rect 59452 11840 59504 11849
rect 56416 11815 56468 11824
rect 56416 11781 56439 11815
rect 56439 11781 56468 11815
rect 56416 11772 56468 11781
rect 57336 11704 57388 11756
rect 57888 11704 57940 11756
rect 37188 11636 37240 11688
rect 42616 11636 42668 11688
rect 30656 11568 30708 11620
rect 34796 11611 34848 11620
rect 30748 11500 30800 11552
rect 31760 11500 31812 11552
rect 33876 11500 33928 11552
rect 34244 11543 34296 11552
rect 34244 11509 34253 11543
rect 34253 11509 34287 11543
rect 34287 11509 34296 11543
rect 34244 11500 34296 11509
rect 34796 11577 34805 11611
rect 34805 11577 34839 11611
rect 34839 11577 34848 11611
rect 34796 11568 34848 11577
rect 36544 11500 36596 11552
rect 37832 11543 37884 11552
rect 37832 11509 37841 11543
rect 37841 11509 37875 11543
rect 37875 11509 37884 11543
rect 37832 11500 37884 11509
rect 39304 11568 39356 11620
rect 41328 11568 41380 11620
rect 39212 11500 39264 11552
rect 42432 11500 42484 11552
rect 44364 11636 44416 11688
rect 46664 11636 46716 11688
rect 49240 11636 49292 11688
rect 49792 11679 49844 11688
rect 49792 11645 49801 11679
rect 49801 11645 49835 11679
rect 49835 11645 49844 11679
rect 49792 11636 49844 11645
rect 51080 11636 51132 11688
rect 51540 11636 51592 11688
rect 52092 11636 52144 11688
rect 53012 11636 53064 11688
rect 54024 11636 54076 11688
rect 55772 11636 55824 11688
rect 56140 11679 56192 11688
rect 56140 11645 56149 11679
rect 56149 11645 56183 11679
rect 56183 11645 56192 11679
rect 56140 11636 56192 11645
rect 59544 11704 59596 11756
rect 60004 11840 60056 11892
rect 60924 11840 60976 11892
rect 61016 11840 61068 11892
rect 61292 11840 61344 11892
rect 62304 11840 62356 11892
rect 62580 11840 62632 11892
rect 60096 11772 60148 11824
rect 60648 11747 60700 11756
rect 60648 11713 60657 11747
rect 60657 11713 60691 11747
rect 60691 11713 60700 11747
rect 60648 11704 60700 11713
rect 61568 11747 61620 11756
rect 46756 11568 46808 11620
rect 46020 11500 46072 11552
rect 46388 11500 46440 11552
rect 47584 11500 47636 11552
rect 47676 11500 47728 11552
rect 48780 11568 48832 11620
rect 61568 11713 61602 11747
rect 61602 11713 61620 11747
rect 61568 11704 61620 11713
rect 61936 11704 61988 11756
rect 67180 11772 67232 11824
rect 61016 11636 61068 11688
rect 61292 11679 61344 11688
rect 61292 11645 61301 11679
rect 61301 11645 61335 11679
rect 61335 11645 61344 11679
rect 61292 11636 61344 11645
rect 62304 11636 62356 11688
rect 65708 11704 65760 11756
rect 70952 11840 71004 11892
rect 49056 11500 49108 11552
rect 52552 11500 52604 11552
rect 54392 11500 54444 11552
rect 60372 11568 60424 11620
rect 60096 11500 60148 11552
rect 60556 11500 60608 11552
rect 68560 11747 68612 11756
rect 68560 11713 68569 11747
rect 68569 11713 68603 11747
rect 68603 11713 68612 11747
rect 68560 11704 68612 11713
rect 72332 11815 72384 11824
rect 72332 11781 72341 11815
rect 72341 11781 72375 11815
rect 72375 11781 72384 11815
rect 72332 11772 72384 11781
rect 72608 11772 72660 11824
rect 74724 11772 74776 11824
rect 78772 11772 78824 11824
rect 78956 11840 79008 11892
rect 81348 11840 81400 11892
rect 82636 11840 82688 11892
rect 84200 11840 84252 11892
rect 86408 11840 86460 11892
rect 86868 11840 86920 11892
rect 88984 11883 89036 11892
rect 88984 11849 88993 11883
rect 88993 11849 89027 11883
rect 89027 11849 89036 11883
rect 88984 11840 89036 11849
rect 81440 11772 81492 11824
rect 68928 11636 68980 11688
rect 70952 11636 71004 11688
rect 72700 11636 72752 11688
rect 63592 11500 63644 11552
rect 65064 11543 65116 11552
rect 65064 11509 65073 11543
rect 65073 11509 65107 11543
rect 65107 11509 65116 11543
rect 65064 11500 65116 11509
rect 65616 11500 65668 11552
rect 65892 11500 65944 11552
rect 68376 11543 68428 11552
rect 68376 11509 68385 11543
rect 68385 11509 68419 11543
rect 68419 11509 68428 11543
rect 68376 11500 68428 11509
rect 68744 11500 68796 11552
rect 70216 11568 70268 11620
rect 72608 11568 72660 11620
rect 70308 11500 70360 11552
rect 70584 11543 70636 11552
rect 70584 11509 70593 11543
rect 70593 11509 70627 11543
rect 70627 11509 70636 11543
rect 70584 11500 70636 11509
rect 71872 11500 71924 11552
rect 75920 11704 75972 11756
rect 76196 11704 76248 11756
rect 77300 11704 77352 11756
rect 72976 11543 73028 11552
rect 72976 11509 72985 11543
rect 72985 11509 73019 11543
rect 73019 11509 73028 11543
rect 72976 11500 73028 11509
rect 74724 11500 74776 11552
rect 75920 11568 75972 11620
rect 75276 11500 75328 11552
rect 78680 11636 78732 11688
rect 80520 11747 80572 11756
rect 80520 11713 80529 11747
rect 80529 11713 80563 11747
rect 80563 11713 80572 11747
rect 80520 11704 80572 11713
rect 81624 11704 81676 11756
rect 86224 11704 86276 11756
rect 79140 11568 79192 11620
rect 83924 11636 83976 11688
rect 84108 11636 84160 11688
rect 86868 11704 86920 11756
rect 86960 11704 87012 11756
rect 87512 11772 87564 11824
rect 89260 11772 89312 11824
rect 89904 11772 89956 11824
rect 93676 11772 93728 11824
rect 94596 11840 94648 11892
rect 96160 11840 96212 11892
rect 98184 11840 98236 11892
rect 98460 11883 98512 11892
rect 98460 11849 98469 11883
rect 98469 11849 98503 11883
rect 98503 11849 98512 11883
rect 98460 11840 98512 11849
rect 99932 11883 99984 11892
rect 99932 11849 99941 11883
rect 99941 11849 99975 11883
rect 99975 11849 99984 11883
rect 99932 11840 99984 11849
rect 100208 11840 100260 11892
rect 103060 11840 103112 11892
rect 103520 11883 103572 11892
rect 103520 11849 103529 11883
rect 103529 11849 103563 11883
rect 103563 11849 103572 11883
rect 103520 11840 103572 11849
rect 104256 11840 104308 11892
rect 104716 11840 104768 11892
rect 106188 11840 106240 11892
rect 108672 11840 108724 11892
rect 109684 11883 109736 11892
rect 101588 11772 101640 11824
rect 109684 11849 109693 11883
rect 109693 11849 109727 11883
rect 109727 11849 109736 11883
rect 109684 11840 109736 11849
rect 112352 11840 112404 11892
rect 113272 11883 113324 11892
rect 113272 11849 113281 11883
rect 113281 11849 113315 11883
rect 113315 11849 113324 11883
rect 113272 11840 113324 11849
rect 114836 11883 114888 11892
rect 114836 11849 114845 11883
rect 114845 11849 114879 11883
rect 114879 11849 114888 11883
rect 114836 11840 114888 11849
rect 118700 11840 118752 11892
rect 119068 11883 119120 11892
rect 119068 11849 119077 11883
rect 119077 11849 119111 11883
rect 119111 11849 119120 11883
rect 119068 11840 119120 11849
rect 119436 11840 119488 11892
rect 125140 11840 125192 11892
rect 125600 11883 125652 11892
rect 125600 11849 125609 11883
rect 125609 11849 125643 11883
rect 125643 11849 125652 11883
rect 125600 11840 125652 11849
rect 130200 11883 130252 11892
rect 130200 11849 130209 11883
rect 130209 11849 130243 11883
rect 130243 11849 130252 11883
rect 130200 11840 130252 11849
rect 132316 11840 132368 11892
rect 134984 11840 135036 11892
rect 135260 11840 135312 11892
rect 87972 11679 88024 11688
rect 87972 11645 87981 11679
rect 87981 11645 88015 11679
rect 88015 11645 88024 11679
rect 87972 11636 88024 11645
rect 92756 11704 92808 11756
rect 92848 11704 92900 11756
rect 93400 11704 93452 11756
rect 94320 11704 94372 11756
rect 95056 11704 95108 11756
rect 90456 11636 90508 11688
rect 90640 11636 90692 11688
rect 77944 11500 77996 11552
rect 82820 11543 82872 11552
rect 82820 11509 82829 11543
rect 82829 11509 82863 11543
rect 82863 11509 82872 11543
rect 82820 11500 82872 11509
rect 83832 11543 83884 11552
rect 83832 11509 83841 11543
rect 83841 11509 83875 11543
rect 83875 11509 83884 11543
rect 83832 11500 83884 11509
rect 84844 11543 84896 11552
rect 84844 11509 84853 11543
rect 84853 11509 84887 11543
rect 84887 11509 84896 11543
rect 84844 11500 84896 11509
rect 86868 11568 86920 11620
rect 89260 11568 89312 11620
rect 94688 11636 94740 11688
rect 95240 11704 95292 11756
rect 96620 11704 96672 11756
rect 99012 11704 99064 11756
rect 101772 11747 101824 11756
rect 101772 11713 101790 11747
rect 101790 11713 101824 11747
rect 101772 11704 101824 11713
rect 101956 11704 102008 11756
rect 96436 11636 96488 11688
rect 96712 11636 96764 11688
rect 99380 11679 99432 11688
rect 99380 11645 99389 11679
rect 99389 11645 99423 11679
rect 99423 11645 99432 11679
rect 99380 11636 99432 11645
rect 87788 11500 87840 11552
rect 88064 11500 88116 11552
rect 89996 11500 90048 11552
rect 90088 11500 90140 11552
rect 93492 11568 93544 11620
rect 101036 11568 101088 11620
rect 94412 11500 94464 11552
rect 100668 11543 100720 11552
rect 100668 11509 100677 11543
rect 100677 11509 100711 11543
rect 100711 11509 100720 11543
rect 100668 11500 100720 11509
rect 103428 11500 103480 11552
rect 107476 11704 107528 11756
rect 108764 11704 108816 11756
rect 108856 11704 108908 11756
rect 112076 11704 112128 11756
rect 112168 11704 112220 11756
rect 113640 11704 113692 11756
rect 107568 11636 107620 11688
rect 108672 11636 108724 11688
rect 115480 11679 115532 11688
rect 115480 11645 115489 11679
rect 115489 11645 115523 11679
rect 115523 11645 115532 11679
rect 115480 11636 115532 11645
rect 115664 11747 115716 11756
rect 115664 11713 115673 11747
rect 115673 11713 115707 11747
rect 115707 11713 115716 11747
rect 115664 11704 115716 11713
rect 116400 11704 116452 11756
rect 106372 11611 106424 11620
rect 106372 11577 106381 11611
rect 106381 11577 106415 11611
rect 106415 11577 106424 11611
rect 106372 11568 106424 11577
rect 107200 11568 107252 11620
rect 107292 11568 107344 11620
rect 107016 11543 107068 11552
rect 107016 11509 107025 11543
rect 107025 11509 107059 11543
rect 107059 11509 107068 11543
rect 107016 11500 107068 11509
rect 107384 11500 107436 11552
rect 109040 11500 109092 11552
rect 109684 11500 109736 11552
rect 110420 11500 110472 11552
rect 112536 11568 112588 11620
rect 112720 11500 112772 11552
rect 115848 11543 115900 11552
rect 115848 11509 115857 11543
rect 115857 11509 115891 11543
rect 115891 11509 115900 11543
rect 115848 11500 115900 11509
rect 117320 11500 117372 11552
rect 117412 11500 117464 11552
rect 118240 11704 118292 11756
rect 121184 11747 121236 11756
rect 121184 11713 121193 11747
rect 121193 11713 121227 11747
rect 121227 11713 121236 11747
rect 121184 11704 121236 11713
rect 118516 11679 118568 11688
rect 118516 11645 118525 11679
rect 118525 11645 118559 11679
rect 118559 11645 118568 11679
rect 118516 11636 118568 11645
rect 118700 11636 118752 11688
rect 118884 11568 118936 11620
rect 119160 11636 119212 11688
rect 125048 11747 125100 11756
rect 125048 11713 125057 11747
rect 125057 11713 125091 11747
rect 125091 11713 125100 11747
rect 125048 11704 125100 11713
rect 121368 11679 121420 11688
rect 121368 11645 121377 11679
rect 121377 11645 121411 11679
rect 121411 11645 121420 11679
rect 121368 11636 121420 11645
rect 122012 11636 122064 11688
rect 123852 11636 123904 11688
rect 125140 11636 125192 11688
rect 125968 11704 126020 11756
rect 118148 11543 118200 11552
rect 118148 11509 118157 11543
rect 118157 11509 118191 11543
rect 118191 11509 118200 11543
rect 118148 11500 118200 11509
rect 118516 11500 118568 11552
rect 119620 11500 119672 11552
rect 124956 11568 125008 11620
rect 126980 11747 127032 11756
rect 126980 11713 126989 11747
rect 126989 11713 127023 11747
rect 127023 11713 127032 11747
rect 126980 11704 127032 11713
rect 127164 11747 127216 11756
rect 127164 11713 127173 11747
rect 127173 11713 127207 11747
rect 127207 11713 127216 11747
rect 127164 11704 127216 11713
rect 127348 11747 127400 11756
rect 127348 11713 127357 11747
rect 127357 11713 127391 11747
rect 127391 11713 127400 11747
rect 127348 11704 127400 11713
rect 129372 11772 129424 11824
rect 128636 11747 128688 11756
rect 128636 11713 128645 11747
rect 128645 11713 128679 11747
rect 128679 11713 128688 11747
rect 128636 11704 128688 11713
rect 127256 11636 127308 11688
rect 128360 11636 128412 11688
rect 132500 11679 132552 11688
rect 132500 11645 132509 11679
rect 132509 11645 132543 11679
rect 132543 11645 132552 11679
rect 132500 11636 132552 11645
rect 133420 11636 133472 11688
rect 134432 11679 134484 11688
rect 134432 11645 134441 11679
rect 134441 11645 134475 11679
rect 134475 11645 134484 11679
rect 134432 11636 134484 11645
rect 120448 11500 120500 11552
rect 120540 11500 120592 11552
rect 121920 11543 121972 11552
rect 121920 11509 121929 11543
rect 121929 11509 121963 11543
rect 121963 11509 121972 11543
rect 121920 11500 121972 11509
rect 122748 11500 122800 11552
rect 123208 11543 123260 11552
rect 123208 11509 123217 11543
rect 123217 11509 123251 11543
rect 123251 11509 123260 11543
rect 123208 11500 123260 11509
rect 123668 11543 123720 11552
rect 123668 11509 123677 11543
rect 123677 11509 123711 11543
rect 123711 11509 123720 11543
rect 123668 11500 123720 11509
rect 124220 11543 124272 11552
rect 124220 11509 124229 11543
rect 124229 11509 124263 11543
rect 124263 11509 124272 11543
rect 124220 11500 124272 11509
rect 125508 11500 125560 11552
rect 133236 11568 133288 11620
rect 134984 11636 135036 11688
rect 137192 11772 137244 11824
rect 138480 11840 138532 11892
rect 138664 11840 138716 11892
rect 136456 11747 136508 11756
rect 136456 11713 136474 11747
rect 136474 11713 136508 11747
rect 136456 11704 136508 11713
rect 136732 11679 136784 11688
rect 136732 11645 136741 11679
rect 136741 11645 136775 11679
rect 136775 11645 136784 11679
rect 136732 11636 136784 11645
rect 137008 11704 137060 11756
rect 138664 11704 138716 11756
rect 139124 11704 139176 11756
rect 135720 11568 135772 11620
rect 138204 11636 138256 11688
rect 140228 11636 140280 11688
rect 139952 11611 140004 11620
rect 127900 11500 127952 11552
rect 128452 11543 128504 11552
rect 128452 11509 128461 11543
rect 128461 11509 128495 11543
rect 128495 11509 128504 11543
rect 128452 11500 128504 11509
rect 128728 11500 128780 11552
rect 131856 11500 131908 11552
rect 132132 11500 132184 11552
rect 132408 11500 132460 11552
rect 133052 11543 133104 11552
rect 133052 11509 133061 11543
rect 133061 11509 133095 11543
rect 133095 11509 133104 11543
rect 133052 11500 133104 11509
rect 138204 11500 138256 11552
rect 139952 11577 139961 11611
rect 139961 11577 139995 11611
rect 139995 11577 140004 11611
rect 139952 11568 140004 11577
rect 141516 11636 141568 11688
rect 141148 11500 141200 11552
rect 141516 11543 141568 11552
rect 141516 11509 141525 11543
rect 141525 11509 141559 11543
rect 141559 11509 141568 11543
rect 141516 11500 141568 11509
rect 143816 11840 143868 11892
rect 143908 11840 143960 11892
rect 148324 11840 148376 11892
rect 148692 11840 148744 11892
rect 142988 11704 143040 11756
rect 144184 11704 144236 11756
rect 144460 11747 144512 11756
rect 146392 11772 146444 11824
rect 144460 11713 144478 11747
rect 144478 11713 144512 11747
rect 144460 11704 144512 11713
rect 144828 11704 144880 11756
rect 146944 11704 146996 11756
rect 147588 11772 147640 11824
rect 142896 11679 142948 11688
rect 142896 11645 142905 11679
rect 142905 11645 142939 11679
rect 142939 11645 142948 11679
rect 142896 11636 142948 11645
rect 147128 11636 147180 11688
rect 147496 11636 147548 11688
rect 148324 11704 148376 11756
rect 150440 11772 150492 11824
rect 152556 11840 152608 11892
rect 153292 11840 153344 11892
rect 157616 11883 157668 11892
rect 157616 11849 157625 11883
rect 157625 11849 157659 11883
rect 157659 11849 157668 11883
rect 157616 11840 157668 11849
rect 150164 11704 150216 11756
rect 153292 11704 153344 11756
rect 153936 11704 153988 11756
rect 154212 11772 154264 11824
rect 155316 11772 155368 11824
rect 155684 11772 155736 11824
rect 154580 11704 154632 11756
rect 154672 11747 154724 11756
rect 154672 11713 154681 11747
rect 154681 11713 154715 11747
rect 154715 11713 154724 11747
rect 154672 11704 154724 11713
rect 156144 11745 156196 11756
rect 156144 11711 156153 11745
rect 156153 11711 156187 11745
rect 156187 11711 156196 11745
rect 156144 11704 156196 11711
rect 150348 11636 150400 11688
rect 150808 11679 150860 11688
rect 150808 11645 150817 11679
rect 150817 11645 150851 11679
rect 150851 11645 150860 11679
rect 150808 11636 150860 11645
rect 154304 11636 154356 11688
rect 154396 11636 154448 11688
rect 155684 11636 155736 11688
rect 143264 11500 143316 11552
rect 144920 11500 144972 11552
rect 145656 11543 145708 11552
rect 145656 11509 145665 11543
rect 145665 11509 145699 11543
rect 145699 11509 145708 11543
rect 145656 11500 145708 11509
rect 147496 11543 147548 11552
rect 147496 11509 147505 11543
rect 147505 11509 147539 11543
rect 147539 11509 147548 11543
rect 147496 11500 147548 11509
rect 147588 11500 147640 11552
rect 148140 11500 148192 11552
rect 148508 11500 148560 11552
rect 150164 11568 150216 11620
rect 149612 11500 149664 11552
rect 149980 11500 150032 11552
rect 152372 11568 152424 11620
rect 155500 11568 155552 11620
rect 155316 11543 155368 11552
rect 155316 11509 155325 11543
rect 155325 11509 155359 11543
rect 155359 11509 155368 11543
rect 155316 11500 155368 11509
rect 155408 11500 155460 11552
rect 155684 11500 155736 11552
rect 156144 11568 156196 11620
rect 155868 11500 155920 11552
rect 156512 11500 156564 11552
rect 158260 11543 158312 11552
rect 158260 11509 158269 11543
rect 158269 11509 158303 11543
rect 158303 11509 158312 11543
rect 158260 11500 158312 11509
rect 20672 11398 20724 11450
rect 20736 11398 20788 11450
rect 20800 11398 20852 11450
rect 20864 11398 20916 11450
rect 20928 11398 20980 11450
rect 60117 11398 60169 11450
rect 60181 11398 60233 11450
rect 60245 11398 60297 11450
rect 60309 11398 60361 11450
rect 60373 11398 60425 11450
rect 99562 11398 99614 11450
rect 99626 11398 99678 11450
rect 99690 11398 99742 11450
rect 99754 11398 99806 11450
rect 99818 11398 99870 11450
rect 139007 11398 139059 11450
rect 139071 11398 139123 11450
rect 139135 11398 139187 11450
rect 139199 11398 139251 11450
rect 139263 11398 139315 11450
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 11244 11296 11296 11348
rect 8392 11228 8444 11280
rect 13636 11296 13688 11348
rect 25596 11296 25648 11348
rect 28172 11296 28224 11348
rect 17592 11271 17644 11280
rect 4896 11160 4948 11212
rect 10508 11160 10560 11212
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 17592 11237 17601 11271
rect 17601 11237 17635 11271
rect 17635 11237 17644 11271
rect 17592 11228 17644 11237
rect 30932 11296 30984 11348
rect 31392 11296 31444 11348
rect 30748 11228 30800 11280
rect 36176 11296 36228 11348
rect 36728 11296 36780 11348
rect 37832 11296 37884 11348
rect 40040 11296 40092 11348
rect 40776 11296 40828 11348
rect 34888 11228 34940 11280
rect 38568 11228 38620 11280
rect 16212 11203 16264 11212
rect 7748 11092 7800 11144
rect 8208 11092 8260 11144
rect 9588 11092 9640 11144
rect 10876 11092 10928 11144
rect 11888 11092 11940 11144
rect 11060 11024 11112 11076
rect 11152 11024 11204 11076
rect 12256 11092 12308 11144
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 17316 11160 17368 11212
rect 19432 11203 19484 11212
rect 11428 10956 11480 11008
rect 15200 11092 15252 11144
rect 18420 11092 18472 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 20536 11160 20588 11212
rect 21088 11092 21140 11144
rect 24400 11160 24452 11212
rect 29552 11160 29604 11212
rect 13636 10956 13688 11008
rect 18328 11024 18380 11076
rect 18512 11024 18564 11076
rect 20260 11024 20312 11076
rect 21364 11024 21416 11076
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 18604 10956 18656 11008
rect 24584 11092 24636 11144
rect 26608 11135 26660 11144
rect 21916 11067 21968 11076
rect 21916 11033 21950 11067
rect 21950 11033 21968 11067
rect 21916 11024 21968 11033
rect 22100 11024 22152 11076
rect 25136 11067 25188 11076
rect 25136 11033 25145 11067
rect 25145 11033 25179 11067
rect 25179 11033 25188 11067
rect 25136 11024 25188 11033
rect 26240 11024 26292 11076
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 27712 11092 27764 11144
rect 29644 11092 29696 11144
rect 33600 11160 33652 11212
rect 34336 11160 34388 11212
rect 42248 11228 42300 11280
rect 43260 11296 43312 11348
rect 51632 11296 51684 11348
rect 53472 11296 53524 11348
rect 42708 11228 42760 11280
rect 45376 11271 45428 11280
rect 45376 11237 45385 11271
rect 45385 11237 45419 11271
rect 45419 11237 45428 11271
rect 45376 11228 45428 11237
rect 45652 11228 45704 11280
rect 31668 11135 31720 11144
rect 26884 11024 26936 11076
rect 27160 11024 27212 11076
rect 27344 11024 27396 11076
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 31760 11092 31812 11144
rect 22008 10956 22060 11008
rect 27252 10956 27304 11008
rect 29092 10999 29144 11008
rect 29092 10965 29101 10999
rect 29101 10965 29135 10999
rect 29135 10965 29144 10999
rect 29092 10956 29144 10965
rect 29920 11024 29972 11076
rect 31116 11024 31168 11076
rect 34060 11092 34112 11144
rect 34980 11092 35032 11144
rect 35900 11024 35952 11076
rect 35992 11024 36044 11076
rect 37740 11092 37792 11144
rect 37556 11024 37608 11076
rect 31208 10956 31260 11008
rect 31484 10956 31536 11008
rect 33324 10956 33376 11008
rect 33508 10999 33560 11008
rect 33508 10965 33517 10999
rect 33517 10965 33551 10999
rect 33551 10965 33560 10999
rect 33508 10956 33560 10965
rect 33784 10956 33836 11008
rect 39120 11024 39172 11076
rect 41236 11160 41288 11212
rect 41328 11160 41380 11212
rect 42524 11160 42576 11212
rect 40224 11092 40276 11144
rect 41420 11092 41472 11144
rect 41788 11135 41840 11144
rect 41788 11101 41797 11135
rect 41797 11101 41831 11135
rect 41831 11101 41840 11135
rect 41788 11092 41840 11101
rect 40132 11067 40184 11076
rect 37832 10956 37884 11008
rect 40132 11033 40141 11067
rect 40141 11033 40175 11067
rect 40175 11033 40184 11067
rect 40132 11024 40184 11033
rect 40776 10956 40828 11008
rect 41512 10956 41564 11008
rect 42616 10956 42668 11008
rect 48320 11228 48372 11280
rect 48504 11228 48556 11280
rect 48596 11228 48648 11280
rect 47308 11160 47360 11212
rect 49516 11160 49568 11212
rect 49792 11160 49844 11212
rect 51724 11203 51776 11212
rect 51724 11169 51733 11203
rect 51733 11169 51767 11203
rect 51767 11169 51776 11203
rect 51724 11160 51776 11169
rect 55404 11228 55456 11280
rect 59268 11296 59320 11348
rect 60004 11339 60056 11348
rect 60004 11305 60013 11339
rect 60013 11305 60047 11339
rect 60047 11305 60056 11339
rect 60004 11296 60056 11305
rect 62028 11296 62080 11348
rect 58808 11228 58860 11280
rect 45652 11092 45704 11144
rect 45744 11135 45796 11144
rect 45744 11101 45753 11135
rect 45753 11101 45787 11135
rect 45787 11101 45796 11135
rect 46204 11135 46256 11144
rect 45744 11092 45796 11101
rect 46204 11101 46213 11135
rect 46213 11101 46247 11135
rect 46247 11101 46256 11135
rect 46204 11092 46256 11101
rect 46296 11092 46348 11144
rect 48596 11092 48648 11144
rect 48688 11135 48740 11144
rect 48688 11101 48697 11135
rect 48697 11101 48731 11135
rect 48731 11101 48740 11135
rect 48688 11092 48740 11101
rect 49148 11092 49200 11144
rect 43352 11024 43404 11076
rect 45468 11024 45520 11076
rect 46848 11024 46900 11076
rect 48412 10956 48464 11008
rect 48780 11024 48832 11076
rect 49240 11024 49292 11076
rect 50896 11092 50948 11144
rect 48596 10956 48648 11008
rect 50436 10956 50488 11008
rect 51080 11024 51132 11076
rect 55312 11092 55364 11144
rect 55588 11092 55640 11144
rect 57704 11135 57756 11144
rect 52552 11024 52604 11076
rect 55220 11024 55272 11076
rect 55680 11024 55732 11076
rect 57704 11101 57713 11135
rect 57713 11101 57747 11135
rect 57747 11101 57756 11135
rect 57704 11092 57756 11101
rect 58164 11092 58216 11144
rect 58624 11135 58676 11144
rect 58624 11101 58633 11135
rect 58633 11101 58667 11135
rect 58667 11101 58676 11135
rect 58624 11092 58676 11101
rect 58992 11092 59044 11144
rect 62028 11160 62080 11212
rect 56140 11024 56192 11076
rect 62120 11092 62172 11144
rect 62764 11135 62816 11144
rect 62764 11101 62773 11135
rect 62773 11101 62807 11135
rect 62807 11101 62816 11135
rect 62764 11092 62816 11101
rect 63224 11024 63276 11076
rect 65248 11203 65300 11212
rect 65248 11169 65257 11203
rect 65257 11169 65291 11203
rect 65291 11169 65300 11203
rect 70216 11296 70268 11348
rect 70584 11296 70636 11348
rect 81440 11296 81492 11348
rect 81532 11296 81584 11348
rect 65248 11160 65300 11169
rect 64512 11092 64564 11144
rect 66720 11228 66772 11280
rect 66996 11160 67048 11212
rect 68376 11092 68428 11144
rect 68560 11092 68612 11144
rect 75644 11228 75696 11280
rect 83556 11296 83608 11348
rect 87512 11296 87564 11348
rect 70308 11160 70360 11212
rect 71872 11203 71924 11212
rect 71872 11169 71881 11203
rect 71881 11169 71915 11203
rect 71915 11169 71924 11203
rect 71872 11160 71924 11169
rect 73620 11160 73672 11212
rect 84200 11228 84252 11280
rect 86868 11228 86920 11280
rect 88708 11228 88760 11280
rect 90364 11228 90416 11280
rect 90824 11271 90876 11280
rect 90824 11237 90833 11271
rect 90833 11237 90867 11271
rect 90867 11237 90876 11271
rect 90824 11228 90876 11237
rect 92480 11271 92532 11280
rect 92480 11237 92489 11271
rect 92489 11237 92523 11271
rect 92523 11237 92532 11271
rect 92480 11228 92532 11237
rect 94228 11228 94280 11280
rect 95608 11228 95660 11280
rect 96436 11228 96488 11280
rect 96804 11271 96856 11280
rect 96804 11237 96813 11271
rect 96813 11237 96847 11271
rect 96847 11237 96856 11271
rect 96804 11228 96856 11237
rect 101680 11228 101732 11280
rect 107476 11296 107528 11348
rect 107568 11296 107620 11348
rect 108764 11339 108816 11348
rect 108764 11305 108773 11339
rect 108773 11305 108807 11339
rect 108807 11305 108816 11339
rect 108764 11296 108816 11305
rect 109592 11339 109644 11348
rect 109592 11305 109601 11339
rect 109601 11305 109635 11339
rect 109635 11305 109644 11339
rect 109592 11296 109644 11305
rect 112076 11296 112128 11348
rect 113824 11339 113876 11348
rect 113824 11305 113833 11339
rect 113833 11305 113867 11339
rect 113867 11305 113876 11339
rect 113824 11296 113876 11305
rect 114560 11296 114612 11348
rect 115204 11296 115256 11348
rect 77944 11203 77996 11212
rect 77944 11169 77953 11203
rect 77953 11169 77987 11203
rect 77987 11169 77996 11203
rect 77944 11160 77996 11169
rect 55956 10956 56008 11008
rect 56692 10956 56744 11008
rect 61016 10956 61068 11008
rect 62028 10999 62080 11008
rect 62028 10965 62037 10999
rect 62037 10965 62071 10999
rect 62071 10965 62080 10999
rect 62028 10956 62080 10965
rect 63408 10999 63460 11008
rect 63408 10965 63417 10999
rect 63417 10965 63451 10999
rect 63451 10965 63460 10999
rect 63408 10956 63460 10965
rect 63868 10999 63920 11008
rect 63868 10965 63877 10999
rect 63877 10965 63911 10999
rect 63911 10965 63920 10999
rect 63868 10956 63920 10965
rect 64788 11024 64840 11076
rect 66720 11024 66772 11076
rect 69296 11067 69348 11076
rect 69296 11033 69305 11067
rect 69305 11033 69339 11067
rect 69339 11033 69348 11067
rect 69296 11024 69348 11033
rect 70032 11135 70084 11144
rect 70032 11101 70041 11135
rect 70041 11101 70075 11135
rect 70075 11101 70084 11135
rect 70032 11092 70084 11101
rect 72976 11092 73028 11144
rect 75276 11135 75328 11144
rect 75276 11101 75285 11135
rect 75285 11101 75319 11135
rect 75319 11101 75328 11135
rect 75276 11092 75328 11101
rect 76748 11092 76800 11144
rect 78864 11135 78916 11144
rect 78864 11101 78873 11135
rect 78873 11101 78907 11135
rect 78907 11101 78916 11135
rect 78864 11092 78916 11101
rect 83924 11092 83976 11144
rect 86684 11160 86736 11212
rect 98184 11203 98236 11212
rect 90272 11092 90324 11144
rect 90640 11092 90692 11144
rect 98184 11169 98193 11203
rect 98193 11169 98227 11203
rect 98227 11169 98236 11203
rect 98184 11160 98236 11169
rect 102232 11160 102284 11212
rect 103796 11203 103848 11212
rect 72332 11024 72384 11076
rect 74632 11067 74684 11076
rect 74632 11033 74641 11067
rect 74641 11033 74675 11067
rect 74675 11033 74684 11067
rect 74632 11024 74684 11033
rect 77300 11024 77352 11076
rect 82820 11024 82872 11076
rect 83556 11067 83608 11076
rect 83556 11033 83596 11067
rect 83596 11033 83608 11067
rect 83556 11024 83608 11033
rect 85028 11024 85080 11076
rect 88524 11024 88576 11076
rect 93032 11024 93084 11076
rect 93216 11092 93268 11144
rect 98736 11092 98788 11144
rect 101404 11092 101456 11144
rect 103428 11092 103480 11144
rect 103796 11169 103805 11203
rect 103805 11169 103839 11203
rect 103839 11169 103848 11203
rect 103796 11160 103848 11169
rect 106464 11160 106516 11212
rect 106648 11160 106700 11212
rect 109224 11228 109276 11280
rect 105820 11092 105872 11144
rect 68928 10956 68980 11008
rect 70032 10956 70084 11008
rect 74356 10956 74408 11008
rect 75460 10999 75512 11008
rect 75460 10965 75469 10999
rect 75469 10965 75503 10999
rect 75503 10965 75512 10999
rect 75460 10956 75512 10965
rect 77116 10956 77168 11008
rect 81256 10956 81308 11008
rect 81348 10956 81400 11008
rect 84568 10956 84620 11008
rect 84752 10956 84804 11008
rect 84936 10956 84988 11008
rect 89720 10956 89772 11008
rect 90640 10956 90692 11008
rect 92020 10956 92072 11008
rect 94412 11067 94464 11076
rect 94412 11033 94421 11067
rect 94421 11033 94455 11067
rect 94455 11033 94464 11067
rect 94412 11024 94464 11033
rect 98276 11024 98328 11076
rect 94780 10956 94832 11008
rect 98644 10999 98696 11008
rect 98644 10965 98653 10999
rect 98653 10965 98687 10999
rect 98687 10965 98696 10999
rect 98644 10956 98696 10965
rect 98828 10956 98880 11008
rect 99472 10956 99524 11008
rect 101128 10956 101180 11008
rect 103520 11024 103572 11076
rect 105728 11067 105780 11076
rect 103336 10956 103388 11008
rect 105176 10999 105228 11008
rect 105176 10965 105185 10999
rect 105185 10965 105219 10999
rect 105219 10965 105228 10999
rect 105176 10956 105228 10965
rect 105728 11033 105737 11067
rect 105737 11033 105771 11067
rect 105771 11033 105780 11067
rect 105728 11024 105780 11033
rect 106740 11092 106792 11144
rect 108304 11135 108356 11144
rect 108304 11101 108313 11135
rect 108313 11101 108347 11135
rect 108347 11101 108356 11135
rect 108304 11092 108356 11101
rect 108580 11092 108632 11144
rect 109132 11135 109184 11144
rect 106372 11024 106424 11076
rect 107384 11024 107436 11076
rect 109132 11101 109141 11135
rect 109141 11101 109175 11135
rect 109175 11101 109184 11135
rect 109132 11092 109184 11101
rect 109040 11024 109092 11076
rect 111156 11228 111208 11280
rect 111064 11160 111116 11212
rect 109592 11092 109644 11144
rect 111616 11135 111668 11144
rect 111616 11101 111625 11135
rect 111625 11101 111659 11135
rect 111659 11101 111668 11135
rect 111616 11092 111668 11101
rect 113180 11160 113232 11212
rect 113364 11203 113416 11212
rect 113364 11169 113373 11203
rect 113373 11169 113407 11203
rect 113407 11169 113416 11203
rect 113364 11160 113416 11169
rect 115296 11160 115348 11212
rect 118424 11296 118476 11348
rect 115480 11228 115532 11280
rect 115940 11228 115992 11280
rect 116584 11228 116636 11280
rect 117504 11228 117556 11280
rect 119436 11296 119488 11348
rect 119620 11339 119672 11348
rect 119620 11305 119629 11339
rect 119629 11305 119663 11339
rect 119663 11305 119672 11339
rect 119620 11296 119672 11305
rect 121000 11296 121052 11348
rect 129096 11339 129148 11348
rect 118608 11228 118660 11280
rect 115756 11203 115808 11212
rect 115756 11169 115765 11203
rect 115765 11169 115799 11203
rect 115799 11169 115808 11203
rect 115756 11160 115808 11169
rect 115848 11160 115900 11212
rect 118424 11160 118476 11212
rect 110420 11024 110472 11076
rect 111708 11024 111760 11076
rect 112168 11067 112220 11076
rect 112168 11033 112177 11067
rect 112177 11033 112211 11067
rect 112211 11033 112220 11067
rect 112168 11024 112220 11033
rect 105912 10956 105964 11008
rect 111064 10956 111116 11008
rect 111248 10956 111300 11008
rect 115388 11024 115440 11076
rect 117412 11092 117464 11144
rect 117504 11135 117556 11144
rect 117504 11101 117513 11135
rect 117513 11101 117547 11135
rect 117547 11101 117556 11135
rect 117504 11092 117556 11101
rect 117780 11092 117832 11144
rect 120172 11135 120224 11144
rect 120172 11101 120181 11135
rect 120181 11101 120215 11135
rect 120215 11101 120224 11135
rect 120172 11092 120224 11101
rect 123024 11160 123076 11212
rect 125692 11228 125744 11280
rect 129096 11305 129105 11339
rect 129105 11305 129139 11339
rect 129139 11305 129148 11339
rect 129096 11296 129148 11305
rect 129280 11296 129332 11348
rect 132776 11296 132828 11348
rect 133052 11296 133104 11348
rect 134524 11339 134576 11348
rect 134524 11305 134533 11339
rect 134533 11305 134567 11339
rect 134567 11305 134576 11339
rect 134524 11296 134576 11305
rect 134708 11296 134760 11348
rect 137008 11296 137060 11348
rect 138480 11339 138532 11348
rect 138480 11305 138489 11339
rect 138489 11305 138523 11339
rect 138523 11305 138532 11339
rect 138480 11296 138532 11305
rect 139768 11296 139820 11348
rect 121000 11135 121052 11144
rect 121000 11101 121009 11135
rect 121009 11101 121043 11135
rect 121043 11101 121052 11135
rect 121000 11092 121052 11101
rect 121920 11092 121972 11144
rect 122564 11092 122616 11144
rect 122656 11092 122708 11144
rect 124772 11092 124824 11144
rect 115940 10956 115992 11008
rect 117228 11024 117280 11076
rect 117320 11024 117372 11076
rect 119160 11024 119212 11076
rect 119620 11024 119672 11076
rect 116308 10956 116360 11008
rect 121828 10956 121880 11008
rect 122104 11024 122156 11076
rect 125407 11135 125459 11144
rect 125407 11101 125418 11135
rect 125418 11101 125452 11135
rect 125452 11101 125459 11135
rect 125407 11092 125459 11101
rect 125600 11092 125652 11144
rect 126244 11135 126296 11144
rect 126244 11101 126253 11135
rect 126253 11101 126287 11135
rect 126287 11101 126296 11135
rect 127808 11135 127860 11144
rect 126244 11092 126296 11101
rect 127808 11101 127817 11135
rect 127817 11101 127851 11135
rect 127851 11101 127860 11135
rect 127808 11092 127860 11101
rect 128084 11135 128136 11144
rect 128084 11101 128093 11135
rect 128093 11101 128127 11135
rect 128127 11101 128136 11135
rect 128084 11092 128136 11101
rect 128268 11092 128320 11144
rect 129372 11092 129424 11144
rect 132500 11160 132552 11212
rect 130200 11135 130252 11144
rect 130200 11101 130218 11135
rect 130218 11101 130252 11135
rect 130200 11092 130252 11101
rect 130936 11092 130988 11144
rect 122932 10956 122984 11008
rect 125232 11024 125284 11076
rect 125692 11024 125744 11076
rect 125784 11024 125836 11076
rect 126888 11024 126940 11076
rect 130384 11024 130436 11076
rect 130752 11024 130804 11076
rect 133144 11203 133196 11212
rect 133144 11169 133153 11203
rect 133153 11169 133187 11203
rect 133187 11169 133196 11203
rect 133144 11160 133196 11169
rect 137284 11160 137336 11212
rect 138664 11228 138716 11280
rect 141516 11296 141568 11348
rect 147128 11296 147180 11348
rect 147312 11339 147364 11348
rect 147312 11305 147321 11339
rect 147321 11305 147355 11339
rect 147355 11305 147364 11339
rect 147312 11296 147364 11305
rect 147496 11296 147548 11348
rect 147772 11296 147824 11348
rect 149336 11296 149388 11348
rect 143816 11228 143868 11280
rect 133236 11092 133288 11144
rect 138296 11092 138348 11144
rect 139492 11092 139544 11144
rect 123668 10956 123720 11008
rect 125048 10956 125100 11008
rect 129372 10956 129424 11008
rect 130568 10956 130620 11008
rect 133696 11024 133748 11076
rect 134708 11024 134760 11076
rect 135536 11067 135588 11076
rect 135536 11033 135545 11067
rect 135545 11033 135579 11067
rect 135579 11033 135588 11067
rect 135536 11024 135588 11033
rect 135812 11024 135864 11076
rect 136088 11067 136140 11076
rect 136088 11033 136097 11067
rect 136097 11033 136131 11067
rect 136131 11033 136140 11067
rect 136088 11024 136140 11033
rect 140596 11092 140648 11144
rect 141332 11092 141384 11144
rect 141608 11160 141660 11212
rect 144828 11203 144880 11212
rect 140688 11024 140740 11076
rect 141056 11067 141108 11076
rect 141056 11033 141065 11067
rect 141065 11033 141099 11067
rect 141099 11033 141108 11067
rect 141056 11024 141108 11033
rect 141608 11024 141660 11076
rect 142988 11092 143040 11144
rect 144828 11169 144837 11203
rect 144837 11169 144871 11203
rect 144871 11169 144880 11203
rect 144828 11160 144880 11169
rect 144920 11160 144972 11212
rect 146576 11092 146628 11144
rect 146852 11092 146904 11144
rect 144000 11024 144052 11076
rect 144552 11067 144604 11076
rect 144552 11033 144570 11067
rect 144570 11033 144604 11067
rect 144552 11024 144604 11033
rect 148232 11067 148284 11076
rect 148232 11033 148241 11067
rect 148241 11033 148275 11067
rect 148275 11033 148284 11067
rect 148232 11024 148284 11033
rect 148416 11135 148468 11144
rect 148416 11101 148425 11135
rect 148425 11101 148459 11135
rect 148459 11101 148468 11135
rect 148416 11092 148468 11101
rect 149980 11296 150032 11348
rect 150440 11296 150492 11348
rect 150808 11296 150860 11348
rect 150992 11296 151044 11348
rect 153200 11296 153252 11348
rect 153476 11296 153528 11348
rect 149612 11092 149664 11144
rect 151360 11160 151412 11212
rect 152464 11203 152516 11212
rect 152464 11169 152473 11203
rect 152473 11169 152507 11203
rect 152507 11169 152516 11203
rect 152464 11160 152516 11169
rect 151268 11092 151320 11144
rect 155224 11160 155276 11212
rect 155684 11296 155736 11348
rect 156052 11296 156104 11348
rect 159456 11296 159508 11348
rect 158352 11228 158404 11280
rect 155500 11160 155552 11212
rect 149520 11024 149572 11076
rect 134432 10956 134484 11008
rect 134984 10999 135036 11008
rect 134984 10965 134993 10999
rect 134993 10965 135027 10999
rect 135027 10965 135036 10999
rect 134984 10956 135036 10965
rect 135076 10956 135128 11008
rect 141332 10956 141384 11008
rect 143172 10956 143224 11008
rect 143448 10999 143500 11008
rect 143448 10965 143457 10999
rect 143457 10965 143491 10999
rect 143491 10965 143500 10999
rect 143448 10956 143500 10965
rect 145288 10999 145340 11008
rect 145288 10965 145297 10999
rect 145297 10965 145331 10999
rect 145331 10965 145340 10999
rect 145288 10956 145340 10965
rect 145380 10956 145432 11008
rect 149336 10956 149388 11008
rect 151544 10956 151596 11008
rect 154028 11024 154080 11076
rect 154396 11024 154448 11076
rect 155960 11092 156012 11144
rect 156236 11135 156288 11144
rect 156236 11101 156245 11135
rect 156245 11101 156279 11135
rect 156279 11101 156288 11135
rect 156236 11092 156288 11101
rect 158628 11092 158680 11144
rect 154856 11024 154908 11076
rect 156144 11024 156196 11076
rect 156420 11067 156472 11076
rect 156420 11033 156429 11067
rect 156429 11033 156463 11067
rect 156463 11033 156472 11067
rect 156420 11024 156472 11033
rect 155408 10956 155460 11008
rect 157432 10956 157484 11008
rect 40394 10854 40446 10906
rect 40458 10854 40510 10906
rect 40522 10854 40574 10906
rect 40586 10854 40638 10906
rect 40650 10854 40702 10906
rect 79839 10854 79891 10906
rect 79903 10854 79955 10906
rect 79967 10854 80019 10906
rect 80031 10854 80083 10906
rect 80095 10854 80147 10906
rect 119284 10854 119336 10906
rect 119348 10854 119400 10906
rect 119412 10854 119464 10906
rect 119476 10854 119528 10906
rect 119540 10854 119592 10906
rect 158729 10854 158781 10906
rect 158793 10854 158845 10906
rect 158857 10854 158909 10906
rect 158921 10854 158973 10906
rect 158985 10854 159037 10906
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 12256 10752 12308 10804
rect 15292 10795 15344 10804
rect 4160 10684 4212 10736
rect 8392 10616 8444 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 12072 10727 12124 10736
rect 12072 10693 12106 10727
rect 12106 10693 12124 10727
rect 12072 10684 12124 10693
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 18604 10752 18656 10804
rect 16948 10684 17000 10736
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 15384 10616 15436 10668
rect 16580 10616 16632 10668
rect 17040 10616 17092 10668
rect 19432 10752 19484 10804
rect 20536 10752 20588 10804
rect 22008 10752 22060 10804
rect 25136 10752 25188 10804
rect 26608 10795 26660 10804
rect 26608 10761 26617 10795
rect 26617 10761 26651 10795
rect 26651 10761 26660 10795
rect 26608 10752 26660 10761
rect 27620 10752 27672 10804
rect 27712 10752 27764 10804
rect 29092 10752 29144 10804
rect 30104 10752 30156 10804
rect 30196 10752 30248 10804
rect 33232 10752 33284 10804
rect 33324 10752 33376 10804
rect 37648 10752 37700 10804
rect 40040 10795 40092 10804
rect 40040 10761 40049 10795
rect 40049 10761 40083 10795
rect 40083 10761 40092 10795
rect 40040 10752 40092 10761
rect 40408 10752 40460 10804
rect 41512 10752 41564 10804
rect 42616 10752 42668 10804
rect 44824 10752 44876 10804
rect 44916 10752 44968 10804
rect 46112 10752 46164 10804
rect 48504 10752 48556 10804
rect 49424 10752 49476 10804
rect 27252 10684 27304 10736
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 28356 10616 28408 10668
rect 22192 10548 22244 10600
rect 23020 10591 23072 10600
rect 23020 10557 23029 10591
rect 23029 10557 23063 10591
rect 23063 10557 23072 10591
rect 23020 10548 23072 10557
rect 27344 10548 27396 10600
rect 29552 10616 29604 10668
rect 33508 10684 33560 10736
rect 30104 10616 30156 10668
rect 30012 10591 30064 10600
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 15660 10480 15712 10532
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 8208 10412 8260 10464
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 13636 10412 13688 10464
rect 16672 10412 16724 10464
rect 18512 10480 18564 10532
rect 19984 10412 20036 10464
rect 21364 10455 21416 10464
rect 21364 10421 21373 10455
rect 21373 10421 21407 10455
rect 21407 10421 21416 10455
rect 21364 10412 21416 10421
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 25596 10412 25648 10464
rect 26976 10412 27028 10464
rect 27252 10455 27304 10464
rect 27252 10421 27261 10455
rect 27261 10421 27295 10455
rect 27295 10421 27304 10455
rect 27252 10412 27304 10421
rect 31208 10548 31260 10600
rect 33876 10659 33928 10668
rect 33876 10625 33885 10659
rect 33885 10625 33919 10659
rect 33919 10625 33928 10659
rect 33876 10616 33928 10625
rect 33600 10548 33652 10600
rect 34428 10548 34480 10600
rect 40224 10616 40276 10668
rect 41144 10616 41196 10668
rect 41328 10659 41380 10668
rect 41328 10625 41337 10659
rect 41337 10625 41371 10659
rect 41371 10625 41380 10659
rect 41328 10616 41380 10625
rect 45928 10684 45980 10736
rect 46020 10684 46072 10736
rect 48596 10684 48648 10736
rect 52644 10752 52696 10804
rect 55680 10795 55732 10804
rect 55680 10761 55689 10795
rect 55689 10761 55723 10795
rect 55723 10761 55732 10795
rect 55680 10752 55732 10761
rect 56324 10752 56376 10804
rect 57704 10752 57756 10804
rect 58256 10752 58308 10804
rect 59176 10752 59228 10804
rect 81072 10795 81124 10804
rect 53564 10684 53616 10736
rect 35256 10548 35308 10600
rect 41788 10548 41840 10600
rect 44916 10548 44968 10600
rect 31300 10412 31352 10464
rect 40040 10480 40092 10532
rect 41236 10480 41288 10532
rect 33784 10412 33836 10464
rect 36452 10412 36504 10464
rect 39396 10455 39448 10464
rect 39396 10421 39405 10455
rect 39405 10421 39439 10455
rect 39439 10421 39448 10455
rect 39396 10412 39448 10421
rect 40132 10412 40184 10464
rect 40960 10412 41012 10464
rect 41696 10412 41748 10464
rect 42616 10455 42668 10464
rect 42616 10421 42625 10455
rect 42625 10421 42659 10455
rect 42659 10421 42668 10455
rect 42616 10412 42668 10421
rect 45192 10412 45244 10464
rect 45376 10616 45428 10668
rect 47216 10659 47268 10668
rect 47216 10625 47225 10659
rect 47225 10625 47259 10659
rect 47259 10625 47268 10659
rect 47216 10616 47268 10625
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 48412 10659 48464 10668
rect 48412 10625 48421 10659
rect 48421 10625 48455 10659
rect 48455 10625 48464 10659
rect 48412 10616 48464 10625
rect 49884 10616 49936 10668
rect 50436 10659 50488 10668
rect 50436 10625 50445 10659
rect 50445 10625 50479 10659
rect 50479 10625 50488 10659
rect 50436 10616 50488 10625
rect 50896 10659 50948 10668
rect 50896 10625 50905 10659
rect 50905 10625 50939 10659
rect 50939 10625 50948 10659
rect 50896 10616 50948 10625
rect 49424 10548 49476 10600
rect 51908 10659 51960 10668
rect 51908 10625 51917 10659
rect 51917 10625 51951 10659
rect 51951 10625 51960 10659
rect 51908 10616 51960 10625
rect 52644 10616 52696 10668
rect 55220 10684 55272 10736
rect 56048 10616 56100 10668
rect 56508 10684 56560 10736
rect 58072 10684 58124 10736
rect 58348 10616 58400 10668
rect 51172 10548 51224 10600
rect 49516 10480 49568 10532
rect 50436 10480 50488 10532
rect 53012 10548 53064 10600
rect 47860 10412 47912 10464
rect 48044 10412 48096 10464
rect 55312 10548 55364 10600
rect 55772 10548 55824 10600
rect 59084 10616 59136 10668
rect 60004 10616 60056 10668
rect 60740 10684 60792 10736
rect 64236 10684 64288 10736
rect 69296 10684 69348 10736
rect 60648 10616 60700 10668
rect 63868 10659 63920 10668
rect 63868 10625 63877 10659
rect 63877 10625 63911 10659
rect 63911 10625 63920 10659
rect 63868 10616 63920 10625
rect 64144 10616 64196 10668
rect 68928 10616 68980 10668
rect 70492 10616 70544 10668
rect 74448 10684 74500 10736
rect 72608 10616 72660 10668
rect 78956 10684 79008 10736
rect 79140 10727 79192 10736
rect 79140 10693 79149 10727
rect 79149 10693 79183 10727
rect 79183 10693 79192 10727
rect 79140 10684 79192 10693
rect 79876 10684 79928 10736
rect 81072 10761 81081 10795
rect 81081 10761 81115 10795
rect 81115 10761 81124 10795
rect 81072 10752 81124 10761
rect 84936 10752 84988 10804
rect 86684 10752 86736 10804
rect 74632 10616 74684 10668
rect 76196 10659 76248 10668
rect 76196 10625 76205 10659
rect 76205 10625 76239 10659
rect 76239 10625 76248 10659
rect 76196 10616 76248 10625
rect 76472 10616 76524 10668
rect 76748 10659 76800 10668
rect 76748 10625 76757 10659
rect 76757 10625 76791 10659
rect 76791 10625 76800 10659
rect 76748 10616 76800 10625
rect 77852 10616 77904 10668
rect 83832 10684 83884 10736
rect 87236 10684 87288 10736
rect 59176 10548 59228 10600
rect 62212 10548 62264 10600
rect 63408 10548 63460 10600
rect 67180 10591 67232 10600
rect 57428 10480 57480 10532
rect 55312 10412 55364 10464
rect 58072 10412 58124 10464
rect 58624 10480 58676 10532
rect 62488 10523 62540 10532
rect 62488 10489 62497 10523
rect 62497 10489 62531 10523
rect 62531 10489 62540 10523
rect 62488 10480 62540 10489
rect 62028 10412 62080 10464
rect 64604 10412 64656 10464
rect 64696 10455 64748 10464
rect 64696 10421 64705 10455
rect 64705 10421 64739 10455
rect 64739 10421 64748 10455
rect 67180 10557 67189 10591
rect 67189 10557 67223 10591
rect 67223 10557 67232 10591
rect 67180 10548 67232 10557
rect 65800 10523 65852 10532
rect 65800 10489 65809 10523
rect 65809 10489 65843 10523
rect 65843 10489 65852 10523
rect 65800 10480 65852 10489
rect 64696 10412 64748 10421
rect 66260 10412 66312 10464
rect 67824 10455 67876 10464
rect 67824 10421 67833 10455
rect 67833 10421 67867 10455
rect 67867 10421 67876 10455
rect 67824 10412 67876 10421
rect 68376 10412 68428 10464
rect 68744 10412 68796 10464
rect 71780 10548 71832 10600
rect 74356 10548 74408 10600
rect 74724 10480 74776 10532
rect 71780 10455 71832 10464
rect 71780 10421 71789 10455
rect 71789 10421 71823 10455
rect 71823 10421 71832 10455
rect 71780 10412 71832 10421
rect 74816 10455 74868 10464
rect 74816 10421 74825 10455
rect 74825 10421 74859 10455
rect 74859 10421 74868 10455
rect 74816 10412 74868 10421
rect 78864 10548 78916 10600
rect 79692 10591 79744 10600
rect 79692 10557 79701 10591
rect 79701 10557 79735 10591
rect 79735 10557 79744 10591
rect 79692 10548 79744 10557
rect 82544 10591 82596 10600
rect 82544 10557 82553 10591
rect 82553 10557 82587 10591
rect 82587 10557 82596 10591
rect 82544 10548 82596 10557
rect 93216 10795 93268 10804
rect 93216 10761 93225 10795
rect 93225 10761 93259 10795
rect 93259 10761 93268 10795
rect 93216 10752 93268 10761
rect 94412 10752 94464 10804
rect 88340 10684 88392 10736
rect 98828 10684 98880 10736
rect 87696 10616 87748 10668
rect 83004 10548 83056 10600
rect 83372 10548 83424 10600
rect 84844 10548 84896 10600
rect 86868 10548 86920 10600
rect 88432 10616 88484 10668
rect 89168 10616 89220 10668
rect 90456 10616 90508 10668
rect 94320 10616 94372 10668
rect 94780 10616 94832 10668
rect 87236 10523 87288 10532
rect 76380 10412 76432 10464
rect 81900 10455 81952 10464
rect 81900 10421 81909 10455
rect 81909 10421 81943 10455
rect 81943 10421 81952 10455
rect 81900 10412 81952 10421
rect 83832 10412 83884 10464
rect 84568 10412 84620 10464
rect 85304 10455 85356 10464
rect 85304 10421 85313 10455
rect 85313 10421 85347 10455
rect 85347 10421 85356 10455
rect 85304 10412 85356 10421
rect 87236 10489 87245 10523
rect 87245 10489 87279 10523
rect 87279 10489 87288 10523
rect 87236 10480 87288 10489
rect 88892 10548 88944 10600
rect 92020 10591 92072 10600
rect 92020 10557 92029 10591
rect 92029 10557 92063 10591
rect 92063 10557 92072 10591
rect 92020 10548 92072 10557
rect 92296 10548 92348 10600
rect 93032 10548 93084 10600
rect 98828 10548 98880 10600
rect 100852 10795 100904 10804
rect 100852 10761 100861 10795
rect 100861 10761 100895 10795
rect 100895 10761 100904 10795
rect 100852 10752 100904 10761
rect 102140 10752 102192 10804
rect 102232 10752 102284 10804
rect 102324 10684 102376 10736
rect 103796 10752 103848 10804
rect 107752 10752 107804 10804
rect 103428 10684 103480 10736
rect 104348 10684 104400 10736
rect 103336 10659 103388 10668
rect 103336 10625 103345 10659
rect 103345 10625 103379 10659
rect 103379 10625 103388 10659
rect 107568 10684 107620 10736
rect 108948 10752 109000 10804
rect 109040 10752 109092 10804
rect 110604 10752 110656 10804
rect 110880 10752 110932 10804
rect 111524 10752 111576 10804
rect 112720 10752 112772 10804
rect 112904 10752 112956 10804
rect 115296 10752 115348 10804
rect 115664 10752 115716 10804
rect 116216 10752 116268 10804
rect 103336 10616 103388 10625
rect 107476 10616 107528 10668
rect 88340 10412 88392 10464
rect 88524 10412 88576 10464
rect 90272 10412 90324 10464
rect 101128 10480 101180 10532
rect 92756 10455 92808 10464
rect 92756 10421 92765 10455
rect 92765 10421 92799 10455
rect 92799 10421 92808 10455
rect 92756 10412 92808 10421
rect 93952 10412 94004 10464
rect 94872 10455 94924 10464
rect 94872 10421 94881 10455
rect 94881 10421 94915 10455
rect 94915 10421 94924 10455
rect 94872 10412 94924 10421
rect 95332 10412 95384 10464
rect 95516 10412 95568 10464
rect 97080 10412 97132 10464
rect 98276 10455 98328 10464
rect 98276 10421 98285 10455
rect 98285 10421 98319 10455
rect 98319 10421 98328 10455
rect 98276 10412 98328 10421
rect 98368 10412 98420 10464
rect 100852 10412 100904 10464
rect 104072 10548 104124 10600
rect 104532 10548 104584 10600
rect 107844 10548 107896 10600
rect 108212 10616 108264 10668
rect 116952 10684 117004 10736
rect 117688 10752 117740 10804
rect 110604 10659 110656 10668
rect 110604 10625 110613 10659
rect 110613 10625 110647 10659
rect 110647 10625 110656 10659
rect 110604 10616 110656 10625
rect 110880 10616 110932 10668
rect 110972 10616 111024 10668
rect 111432 10659 111484 10668
rect 111432 10625 111441 10659
rect 111441 10625 111475 10659
rect 111475 10625 111484 10659
rect 111432 10616 111484 10625
rect 111524 10659 111576 10668
rect 111524 10625 111533 10659
rect 111533 10625 111567 10659
rect 111567 10625 111576 10659
rect 111524 10616 111576 10625
rect 111800 10616 111852 10668
rect 113732 10616 113784 10668
rect 114560 10616 114612 10668
rect 109132 10548 109184 10600
rect 110420 10591 110472 10600
rect 110420 10557 110429 10591
rect 110429 10557 110463 10591
rect 110463 10557 110472 10591
rect 110420 10548 110472 10557
rect 110696 10548 110748 10600
rect 117872 10616 117924 10668
rect 115664 10548 115716 10600
rect 116216 10548 116268 10600
rect 117320 10591 117372 10600
rect 117320 10557 117329 10591
rect 117329 10557 117363 10591
rect 117363 10557 117372 10591
rect 117320 10548 117372 10557
rect 107476 10480 107528 10532
rect 107844 10412 107896 10464
rect 108488 10412 108540 10464
rect 111616 10480 111668 10532
rect 122656 10752 122708 10804
rect 122932 10752 122984 10804
rect 125692 10752 125744 10804
rect 130200 10795 130252 10804
rect 120172 10684 120224 10736
rect 130200 10761 130209 10795
rect 130209 10761 130243 10795
rect 130243 10761 130252 10795
rect 130200 10752 130252 10761
rect 126796 10684 126848 10736
rect 136180 10752 136232 10804
rect 136916 10752 136968 10804
rect 137652 10752 137704 10804
rect 138664 10752 138716 10804
rect 138756 10752 138808 10804
rect 139860 10752 139912 10804
rect 140780 10752 140832 10804
rect 141332 10752 141384 10804
rect 147312 10752 147364 10804
rect 141240 10684 141292 10736
rect 144920 10684 144972 10736
rect 148784 10752 148836 10804
rect 150256 10752 150308 10804
rect 150716 10752 150768 10804
rect 150900 10752 150952 10804
rect 152556 10752 152608 10804
rect 153936 10752 153988 10804
rect 154580 10752 154632 10804
rect 155316 10795 155368 10804
rect 155316 10761 155325 10795
rect 155325 10761 155359 10795
rect 155359 10761 155368 10795
rect 155316 10752 155368 10761
rect 155684 10752 155736 10804
rect 158260 10795 158312 10804
rect 158260 10761 158269 10795
rect 158269 10761 158303 10795
rect 158303 10761 158312 10795
rect 158260 10752 158312 10761
rect 118608 10616 118660 10668
rect 120540 10659 120592 10668
rect 119160 10591 119212 10600
rect 119160 10557 119169 10591
rect 119169 10557 119203 10591
rect 119203 10557 119212 10591
rect 119160 10548 119212 10557
rect 120540 10625 120549 10659
rect 120549 10625 120583 10659
rect 120583 10625 120592 10659
rect 120540 10616 120592 10625
rect 122104 10659 122156 10668
rect 122104 10625 122122 10659
rect 122122 10625 122156 10659
rect 122104 10616 122156 10625
rect 122288 10616 122340 10668
rect 123760 10616 123812 10668
rect 125232 10616 125284 10668
rect 125692 10616 125744 10668
rect 126152 10616 126204 10668
rect 126888 10659 126940 10668
rect 126888 10625 126897 10659
rect 126897 10625 126931 10659
rect 126931 10625 126940 10659
rect 126888 10616 126940 10625
rect 126980 10616 127032 10668
rect 128084 10616 128136 10668
rect 128360 10616 128412 10668
rect 128452 10616 128504 10668
rect 128912 10616 128964 10668
rect 130568 10616 130620 10668
rect 122380 10591 122432 10600
rect 110604 10412 110656 10464
rect 110788 10455 110840 10464
rect 110788 10421 110797 10455
rect 110797 10421 110831 10455
rect 110831 10421 110840 10455
rect 110788 10412 110840 10421
rect 111340 10412 111392 10464
rect 111432 10412 111484 10464
rect 113456 10412 113508 10464
rect 113824 10412 113876 10464
rect 115848 10412 115900 10464
rect 117872 10412 117924 10464
rect 120172 10412 120224 10464
rect 120356 10455 120408 10464
rect 120356 10421 120365 10455
rect 120365 10421 120399 10455
rect 120399 10421 120408 10455
rect 120356 10412 120408 10421
rect 121000 10455 121052 10464
rect 121000 10421 121009 10455
rect 121009 10421 121043 10455
rect 121043 10421 121052 10455
rect 121000 10412 121052 10421
rect 122380 10557 122389 10591
rect 122389 10557 122423 10591
rect 122423 10557 122432 10591
rect 122380 10548 122432 10557
rect 125600 10548 125652 10600
rect 132408 10616 132460 10668
rect 122564 10480 122616 10532
rect 122840 10412 122892 10464
rect 123668 10455 123720 10464
rect 123668 10421 123677 10455
rect 123677 10421 123711 10455
rect 123711 10421 123720 10455
rect 123668 10412 123720 10421
rect 123760 10412 123812 10464
rect 125600 10412 125652 10464
rect 127072 10480 127124 10532
rect 126152 10412 126204 10464
rect 127532 10412 127584 10464
rect 128176 10412 128228 10464
rect 130200 10412 130252 10464
rect 130292 10412 130344 10464
rect 136732 10548 136784 10600
rect 138020 10616 138072 10668
rect 137652 10548 137704 10600
rect 140320 10616 140372 10668
rect 141148 10659 141200 10668
rect 139492 10548 139544 10600
rect 140504 10548 140556 10600
rect 141148 10625 141157 10659
rect 141157 10625 141191 10659
rect 141191 10625 141200 10659
rect 141148 10616 141200 10625
rect 141332 10616 141384 10668
rect 144184 10659 144236 10668
rect 144184 10625 144193 10659
rect 144193 10625 144227 10659
rect 144227 10625 144236 10659
rect 144184 10616 144236 10625
rect 144736 10616 144788 10668
rect 145196 10616 145248 10668
rect 146944 10616 146996 10668
rect 133052 10412 133104 10464
rect 133696 10455 133748 10464
rect 133696 10421 133705 10455
rect 133705 10421 133739 10455
rect 133739 10421 133748 10455
rect 133696 10412 133748 10421
rect 134984 10412 135036 10464
rect 135536 10412 135588 10464
rect 136548 10412 136600 10464
rect 136640 10412 136692 10464
rect 138664 10480 138716 10532
rect 139860 10412 139912 10464
rect 139952 10412 140004 10464
rect 141332 10412 141384 10464
rect 142896 10412 142948 10464
rect 143540 10480 143592 10532
rect 146668 10548 146720 10600
rect 149428 10659 149480 10668
rect 149428 10625 149437 10659
rect 149437 10625 149471 10659
rect 149471 10625 149480 10659
rect 149428 10616 149480 10625
rect 150164 10616 150216 10668
rect 155408 10684 155460 10736
rect 150440 10548 150492 10600
rect 151636 10616 151688 10668
rect 152096 10616 152148 10668
rect 152464 10616 152516 10668
rect 154396 10616 154448 10668
rect 154672 10659 154724 10668
rect 154672 10625 154681 10659
rect 154681 10625 154715 10659
rect 154715 10625 154724 10659
rect 154672 10616 154724 10625
rect 156144 10659 156196 10668
rect 154028 10591 154080 10600
rect 146852 10412 146904 10464
rect 147036 10455 147088 10464
rect 147036 10421 147045 10455
rect 147045 10421 147079 10455
rect 147079 10421 147088 10455
rect 147036 10412 147088 10421
rect 149980 10480 150032 10532
rect 150900 10480 150952 10532
rect 149060 10412 149112 10464
rect 150256 10412 150308 10464
rect 154028 10557 154037 10591
rect 154037 10557 154071 10591
rect 154071 10557 154080 10591
rect 154028 10548 154080 10557
rect 154212 10548 154264 10600
rect 156144 10625 156153 10659
rect 156153 10625 156187 10659
rect 156187 10625 156196 10659
rect 156144 10616 156196 10625
rect 156972 10659 157024 10668
rect 156972 10625 156981 10659
rect 156981 10625 157015 10659
rect 157015 10625 157024 10659
rect 156972 10616 157024 10625
rect 159088 10616 159140 10668
rect 152648 10523 152700 10532
rect 152648 10489 152657 10523
rect 152657 10489 152691 10523
rect 152691 10489 152700 10523
rect 152648 10480 152700 10489
rect 154304 10480 154356 10532
rect 158444 10480 158496 10532
rect 152280 10412 152332 10464
rect 155224 10412 155276 10464
rect 155408 10412 155460 10464
rect 155868 10412 155920 10464
rect 157156 10455 157208 10464
rect 157156 10421 157165 10455
rect 157165 10421 157199 10455
rect 157199 10421 157208 10455
rect 157156 10412 157208 10421
rect 20672 10310 20724 10362
rect 20736 10310 20788 10362
rect 20800 10310 20852 10362
rect 20864 10310 20916 10362
rect 20928 10310 20980 10362
rect 60117 10310 60169 10362
rect 60181 10310 60233 10362
rect 60245 10310 60297 10362
rect 60309 10310 60361 10362
rect 60373 10310 60425 10362
rect 99562 10310 99614 10362
rect 99626 10310 99678 10362
rect 99690 10310 99742 10362
rect 99754 10310 99806 10362
rect 99818 10310 99870 10362
rect 139007 10310 139059 10362
rect 139071 10310 139123 10362
rect 139135 10310 139187 10362
rect 139199 10310 139251 10362
rect 139263 10310 139315 10362
rect 5724 10208 5776 10260
rect 9496 10208 9548 10260
rect 13636 10140 13688 10192
rect 16764 10140 16816 10192
rect 17316 10140 17368 10192
rect 3792 10004 3844 10056
rect 5724 10004 5776 10056
rect 1584 9936 1636 9988
rect 4988 9936 5040 9988
rect 8208 9936 8260 9988
rect 14188 10072 14240 10124
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 15108 10004 15160 10056
rect 16948 10072 17000 10124
rect 17040 10072 17092 10124
rect 18144 10072 18196 10124
rect 16672 10004 16724 10056
rect 19340 10004 19392 10056
rect 20076 10208 20128 10260
rect 23756 10208 23808 10260
rect 24584 10208 24636 10260
rect 27252 10208 27304 10260
rect 27344 10208 27396 10260
rect 30840 10208 30892 10260
rect 30196 10140 30248 10192
rect 25136 10004 25188 10056
rect 29460 10004 29512 10056
rect 29552 10004 29604 10056
rect 39396 10208 39448 10260
rect 40408 10208 40460 10260
rect 40776 10208 40828 10260
rect 41052 10208 41104 10260
rect 41420 10251 41472 10260
rect 41420 10217 41429 10251
rect 41429 10217 41463 10251
rect 41463 10217 41472 10251
rect 41420 10208 41472 10217
rect 33232 10140 33284 10192
rect 36268 10140 36320 10192
rect 41236 10140 41288 10192
rect 44456 10208 44508 10260
rect 46020 10208 46072 10260
rect 46572 10208 46624 10260
rect 47492 10208 47544 10260
rect 48688 10208 48740 10260
rect 50344 10208 50396 10260
rect 51264 10251 51316 10260
rect 51264 10217 51273 10251
rect 51273 10217 51307 10251
rect 51307 10217 51316 10251
rect 51264 10208 51316 10217
rect 52460 10208 52512 10260
rect 38568 10072 38620 10124
rect 31300 10004 31352 10056
rect 32772 10047 32824 10056
rect 32772 10013 32781 10047
rect 32781 10013 32815 10047
rect 32815 10013 32824 10047
rect 32772 10004 32824 10013
rect 12532 9936 12584 9988
rect 5448 9868 5500 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 13544 9868 13596 9920
rect 16856 9936 16908 9988
rect 18512 9936 18564 9988
rect 17132 9911 17184 9920
rect 17132 9877 17141 9911
rect 17141 9877 17175 9911
rect 17175 9877 17184 9911
rect 17132 9868 17184 9877
rect 19340 9868 19392 9920
rect 20076 9911 20128 9920
rect 20076 9877 20085 9911
rect 20085 9877 20119 9911
rect 20119 9877 20128 9911
rect 20076 9868 20128 9877
rect 25688 9868 25740 9920
rect 29000 9868 29052 9920
rect 29276 9868 29328 9920
rect 30104 9868 30156 9920
rect 31576 9936 31628 9988
rect 32036 9911 32088 9920
rect 32036 9877 32045 9911
rect 32045 9877 32079 9911
rect 32079 9877 32088 9911
rect 32036 9868 32088 9877
rect 35348 10004 35400 10056
rect 35900 10004 35952 10056
rect 33600 9868 33652 9920
rect 34520 9936 34572 9988
rect 36636 9936 36688 9988
rect 41052 10004 41104 10056
rect 42708 10004 42760 10056
rect 43168 10004 43220 10056
rect 43536 10047 43588 10056
rect 43536 10013 43570 10047
rect 43570 10013 43588 10047
rect 43536 10004 43588 10013
rect 44640 10004 44692 10056
rect 44916 10004 44968 10056
rect 46112 10004 46164 10056
rect 48780 10140 48832 10192
rect 46940 10047 46992 10056
rect 46940 10013 46949 10047
rect 46949 10013 46983 10047
rect 46983 10013 46992 10047
rect 46940 10004 46992 10013
rect 47308 10004 47360 10056
rect 47492 10004 47544 10056
rect 48228 10072 48280 10124
rect 34980 9911 35032 9920
rect 34980 9877 34989 9911
rect 34989 9877 35023 9911
rect 35023 9877 35032 9911
rect 34980 9868 35032 9877
rect 35900 9868 35952 9920
rect 39396 9911 39448 9920
rect 39396 9877 39405 9911
rect 39405 9877 39439 9911
rect 39439 9877 39448 9911
rect 39396 9868 39448 9877
rect 41788 9868 41840 9920
rect 47860 9936 47912 9988
rect 49148 9936 49200 9988
rect 49516 9979 49568 9988
rect 49516 9945 49534 9979
rect 49534 9945 49568 9979
rect 49516 9936 49568 9945
rect 49700 10004 49752 10056
rect 52460 10072 52512 10124
rect 49976 10004 50028 10056
rect 51172 10004 51224 10056
rect 51448 10004 51500 10056
rect 52000 10047 52052 10056
rect 52000 10013 52009 10047
rect 52009 10013 52043 10047
rect 52043 10013 52052 10047
rect 52000 10004 52052 10013
rect 64236 10208 64288 10260
rect 54024 10183 54076 10192
rect 54024 10149 54033 10183
rect 54033 10149 54067 10183
rect 54067 10149 54076 10183
rect 54024 10140 54076 10149
rect 55956 10140 56008 10192
rect 56232 10183 56284 10192
rect 56232 10149 56241 10183
rect 56241 10149 56275 10183
rect 56275 10149 56284 10183
rect 56232 10140 56284 10149
rect 52644 10115 52696 10124
rect 52644 10081 52653 10115
rect 52653 10081 52687 10115
rect 52687 10081 52696 10115
rect 52644 10072 52696 10081
rect 54392 10072 54444 10124
rect 57060 10140 57112 10192
rect 57612 10140 57664 10192
rect 57888 10183 57940 10192
rect 57888 10149 57897 10183
rect 57897 10149 57931 10183
rect 57931 10149 57940 10183
rect 57888 10140 57940 10149
rect 58716 10140 58768 10192
rect 59820 10140 59872 10192
rect 62028 10183 62080 10192
rect 62028 10149 62037 10183
rect 62037 10149 62071 10183
rect 62071 10149 62080 10183
rect 62028 10140 62080 10149
rect 74816 10208 74868 10260
rect 60648 10115 60700 10124
rect 53196 9936 53248 9988
rect 53288 9936 53340 9988
rect 55036 10004 55088 10056
rect 54576 9936 54628 9988
rect 56692 10004 56744 10056
rect 56876 10004 56928 10056
rect 58808 10047 58860 10056
rect 45560 9868 45612 9920
rect 48412 9911 48464 9920
rect 48412 9877 48421 9911
rect 48421 9877 48455 9911
rect 48455 9877 48464 9911
rect 48412 9868 48464 9877
rect 50620 9868 50672 9920
rect 54392 9868 54444 9920
rect 54852 9911 54904 9920
rect 54852 9877 54861 9911
rect 54861 9877 54895 9911
rect 54895 9877 54904 9911
rect 54852 9868 54904 9877
rect 54944 9868 54996 9920
rect 58808 10013 58817 10047
rect 58817 10013 58851 10047
rect 58851 10013 58860 10047
rect 58808 10004 58860 10013
rect 60648 10081 60657 10115
rect 60657 10081 60691 10115
rect 60691 10081 60700 10115
rect 60648 10072 60700 10081
rect 68836 10140 68888 10192
rect 73712 10140 73764 10192
rect 74724 10140 74776 10192
rect 75828 10140 75880 10192
rect 62396 10072 62448 10124
rect 65248 10115 65300 10124
rect 63040 10047 63092 10056
rect 57704 9979 57756 9988
rect 57704 9945 57713 9979
rect 57713 9945 57747 9979
rect 57747 9945 57756 9979
rect 57704 9936 57756 9945
rect 57796 9936 57848 9988
rect 57060 9868 57112 9920
rect 57520 9868 57572 9920
rect 57612 9868 57664 9920
rect 60464 9868 60516 9920
rect 60648 9868 60700 9920
rect 61016 9868 61068 9920
rect 63040 10013 63049 10047
rect 63049 10013 63083 10047
rect 63083 10013 63092 10047
rect 63040 10004 63092 10013
rect 65248 10081 65257 10115
rect 65257 10081 65291 10115
rect 65291 10081 65300 10115
rect 65248 10072 65300 10081
rect 67180 10115 67232 10124
rect 67180 10081 67189 10115
rect 67189 10081 67223 10115
rect 67223 10081 67232 10115
rect 67180 10072 67232 10081
rect 64696 10004 64748 10056
rect 62580 9868 62632 9920
rect 63408 9911 63460 9920
rect 63408 9877 63417 9911
rect 63417 9877 63451 9911
rect 63451 9877 63460 9911
rect 63408 9868 63460 9877
rect 63960 9936 64012 9988
rect 66720 9936 66772 9988
rect 69020 10072 69072 10124
rect 69480 10072 69532 10124
rect 71228 10047 71280 10056
rect 71228 10013 71237 10047
rect 71237 10013 71271 10047
rect 71271 10013 71280 10047
rect 71228 10004 71280 10013
rect 73436 9936 73488 9988
rect 64420 9868 64472 9920
rect 66076 9868 66128 9920
rect 67732 9868 67784 9920
rect 67824 9868 67876 9920
rect 70032 9868 70084 9920
rect 71780 9868 71832 9920
rect 72608 9911 72660 9920
rect 72608 9877 72617 9911
rect 72617 9877 72651 9911
rect 72651 9877 72660 9911
rect 72608 9868 72660 9877
rect 73160 9911 73212 9920
rect 73160 9877 73169 9911
rect 73169 9877 73203 9911
rect 73203 9877 73212 9911
rect 76380 10047 76432 10056
rect 76380 10013 76389 10047
rect 76389 10013 76423 10047
rect 76423 10013 76432 10047
rect 76380 10004 76432 10013
rect 76656 10004 76708 10056
rect 74724 9936 74776 9988
rect 73160 9868 73212 9877
rect 75184 9868 75236 9920
rect 76564 9868 76616 9920
rect 84108 10208 84160 10260
rect 84568 10208 84620 10260
rect 100760 10251 100812 10260
rect 82728 10140 82780 10192
rect 83096 10140 83148 10192
rect 84752 10140 84804 10192
rect 86408 10140 86460 10192
rect 86776 10140 86828 10192
rect 89720 10183 89772 10192
rect 89720 10149 89729 10183
rect 89729 10149 89763 10183
rect 89763 10149 89772 10183
rect 89720 10140 89772 10149
rect 90548 10140 90600 10192
rect 92848 10183 92900 10192
rect 92848 10149 92857 10183
rect 92857 10149 92891 10183
rect 92891 10149 92900 10183
rect 92848 10140 92900 10149
rect 86960 10072 87012 10124
rect 89536 10072 89588 10124
rect 93216 10072 93268 10124
rect 81256 10047 81308 10056
rect 81256 10013 81265 10047
rect 81265 10013 81299 10047
rect 81299 10013 81308 10047
rect 81256 10004 81308 10013
rect 84568 10004 84620 10056
rect 84752 10004 84804 10056
rect 85488 10004 85540 10056
rect 91652 10047 91704 10056
rect 91652 10013 91661 10047
rect 91661 10013 91695 10047
rect 91695 10013 91704 10047
rect 91652 10004 91704 10013
rect 93584 10004 93636 10056
rect 94872 10004 94924 10056
rect 98828 10183 98880 10192
rect 98828 10149 98837 10183
rect 98837 10149 98871 10183
rect 98871 10149 98880 10183
rect 98828 10140 98880 10149
rect 100760 10217 100769 10251
rect 100769 10217 100803 10251
rect 100803 10217 100812 10251
rect 100760 10208 100812 10217
rect 101128 10140 101180 10192
rect 98368 10072 98420 10124
rect 102232 10208 102284 10260
rect 102876 10208 102928 10260
rect 104348 10251 104400 10260
rect 101864 10183 101916 10192
rect 101864 10149 101873 10183
rect 101873 10149 101907 10183
rect 101907 10149 101916 10183
rect 101864 10140 101916 10149
rect 104348 10217 104357 10251
rect 104357 10217 104391 10251
rect 104391 10217 104400 10251
rect 104348 10208 104400 10217
rect 104532 10208 104584 10260
rect 106832 10208 106884 10260
rect 107568 10208 107620 10260
rect 107752 10208 107804 10260
rect 112536 10251 112588 10260
rect 105912 10140 105964 10192
rect 103428 10072 103480 10124
rect 104072 10072 104124 10124
rect 107476 10072 107528 10124
rect 110696 10140 110748 10192
rect 111248 10140 111300 10192
rect 112536 10217 112545 10251
rect 112545 10217 112579 10251
rect 112579 10217 112588 10251
rect 112536 10208 112588 10217
rect 112996 10140 113048 10192
rect 97080 10047 97132 10056
rect 97080 10013 97089 10047
rect 97089 10013 97123 10047
rect 97123 10013 97132 10047
rect 97080 10004 97132 10013
rect 79600 9936 79652 9988
rect 81900 9936 81952 9988
rect 77852 9911 77904 9920
rect 77852 9877 77861 9911
rect 77861 9877 77895 9911
rect 77895 9877 77904 9911
rect 77852 9868 77904 9877
rect 83096 9911 83148 9920
rect 83096 9877 83105 9911
rect 83105 9877 83139 9911
rect 83139 9877 83148 9911
rect 83096 9868 83148 9877
rect 83464 9868 83516 9920
rect 84844 9936 84896 9988
rect 88340 9936 88392 9988
rect 87696 9868 87748 9920
rect 87880 9911 87932 9920
rect 87880 9877 87889 9911
rect 87889 9877 87923 9911
rect 87923 9877 87932 9911
rect 87880 9868 87932 9877
rect 87972 9868 88024 9920
rect 90824 9936 90876 9988
rect 93860 9936 93912 9988
rect 93952 9979 94004 9988
rect 93952 9945 93970 9979
rect 93970 9945 94004 9979
rect 98276 10004 98328 10056
rect 115572 10072 115624 10124
rect 108396 10047 108448 10056
rect 108396 10013 108405 10047
rect 108405 10013 108439 10047
rect 108439 10013 108448 10047
rect 108396 10004 108448 10013
rect 110420 10004 110472 10056
rect 110604 10004 110656 10056
rect 111524 10004 111576 10056
rect 111616 10004 111668 10056
rect 112904 10004 112956 10056
rect 113548 10004 113600 10056
rect 114744 10004 114796 10056
rect 115848 10072 115900 10124
rect 118516 10208 118568 10260
rect 122564 10208 122616 10260
rect 122932 10208 122984 10260
rect 118792 10140 118844 10192
rect 118976 10140 119028 10192
rect 115940 10004 115992 10056
rect 120724 10072 120776 10124
rect 117228 10004 117280 10056
rect 93952 9936 94004 9945
rect 91100 9868 91152 9920
rect 92388 9868 92440 9920
rect 94872 9868 94924 9920
rect 95700 9868 95752 9920
rect 96160 9911 96212 9920
rect 96160 9877 96169 9911
rect 96169 9877 96203 9911
rect 96203 9877 96212 9911
rect 96160 9868 96212 9877
rect 99472 9936 99524 9988
rect 100760 9936 100812 9988
rect 101128 9936 101180 9988
rect 102876 9936 102928 9988
rect 103428 9936 103480 9988
rect 98092 9868 98144 9920
rect 104532 9868 104584 9920
rect 104808 9911 104860 9920
rect 104808 9877 104817 9911
rect 104817 9877 104851 9911
rect 104851 9877 104860 9911
rect 104808 9868 104860 9877
rect 104992 9936 105044 9988
rect 107752 9936 107804 9988
rect 108672 9979 108724 9988
rect 108672 9945 108706 9979
rect 108706 9945 108724 9979
rect 108672 9936 108724 9945
rect 110328 9936 110380 9988
rect 113916 9936 113968 9988
rect 115848 9936 115900 9988
rect 116032 9936 116084 9988
rect 118608 10004 118660 10056
rect 119160 10047 119212 10056
rect 119160 10013 119169 10047
rect 119169 10013 119203 10047
rect 119203 10013 119212 10047
rect 119160 10004 119212 10013
rect 121092 10047 121144 10056
rect 121092 10013 121101 10047
rect 121101 10013 121135 10047
rect 121135 10013 121144 10047
rect 121092 10004 121144 10013
rect 122288 10140 122340 10192
rect 123392 10140 123444 10192
rect 123760 10140 123812 10192
rect 126152 10208 126204 10260
rect 133696 10208 133748 10260
rect 133788 10208 133840 10260
rect 128176 10140 128228 10192
rect 128360 10183 128412 10192
rect 128360 10149 128369 10183
rect 128369 10149 128403 10183
rect 128403 10149 128412 10183
rect 137744 10208 137796 10260
rect 140320 10208 140372 10260
rect 140504 10208 140556 10260
rect 128360 10140 128412 10149
rect 121920 10072 121972 10124
rect 122380 10072 122432 10124
rect 122748 10072 122800 10124
rect 122564 10004 122616 10056
rect 122840 10004 122892 10056
rect 128084 10072 128136 10124
rect 130200 10072 130252 10124
rect 137560 10072 137612 10124
rect 140872 10140 140924 10192
rect 142160 10208 142212 10260
rect 108212 9868 108264 9920
rect 108764 9868 108816 9920
rect 110696 9868 110748 9920
rect 110880 9911 110932 9920
rect 110880 9877 110889 9911
rect 110889 9877 110923 9911
rect 110923 9877 110932 9911
rect 110880 9868 110932 9877
rect 113088 9911 113140 9920
rect 113088 9877 113097 9911
rect 113097 9877 113131 9911
rect 113131 9877 113140 9911
rect 113088 9868 113140 9877
rect 113548 9868 113600 9920
rect 114100 9868 114152 9920
rect 115480 9911 115532 9920
rect 115480 9877 115489 9911
rect 115489 9877 115523 9911
rect 115523 9877 115532 9911
rect 115480 9868 115532 9877
rect 115572 9868 115624 9920
rect 118332 9936 118384 9988
rect 117412 9868 117464 9920
rect 117964 9868 118016 9920
rect 120448 9936 120500 9988
rect 123576 9936 123628 9988
rect 119988 9868 120040 9920
rect 121552 9868 121604 9920
rect 124404 9911 124456 9920
rect 124404 9877 124413 9911
rect 124413 9877 124447 9911
rect 124447 9877 124456 9911
rect 124404 9868 124456 9877
rect 129740 10047 129792 10056
rect 129740 10013 129749 10047
rect 129749 10013 129783 10047
rect 129783 10013 129792 10047
rect 130016 10047 130068 10056
rect 129740 10004 129792 10013
rect 130016 10013 130025 10047
rect 130025 10013 130059 10047
rect 130059 10013 130068 10047
rect 130016 10004 130068 10013
rect 130568 10004 130620 10056
rect 130936 10004 130988 10056
rect 132684 10004 132736 10056
rect 134156 10004 134208 10056
rect 135444 10004 135496 10056
rect 135536 10047 135588 10056
rect 135536 10013 135545 10047
rect 135545 10013 135579 10047
rect 135579 10013 135588 10047
rect 135536 10004 135588 10013
rect 126428 9868 126480 9920
rect 126796 9868 126848 9920
rect 132776 9936 132828 9988
rect 134064 9936 134116 9988
rect 135628 9936 135680 9988
rect 133512 9911 133564 9920
rect 133512 9877 133521 9911
rect 133521 9877 133555 9911
rect 133555 9877 133564 9911
rect 133512 9868 133564 9877
rect 133972 9868 134024 9920
rect 134708 9868 134760 9920
rect 136272 9979 136324 9988
rect 136272 9945 136306 9979
rect 136306 9945 136324 9979
rect 140044 10004 140096 10056
rect 144368 10140 144420 10192
rect 144920 10140 144972 10192
rect 146668 10208 146720 10260
rect 147036 10251 147088 10260
rect 147036 10217 147045 10251
rect 147045 10217 147079 10251
rect 147079 10217 147088 10251
rect 147036 10208 147088 10217
rect 147772 10208 147824 10260
rect 147864 10208 147916 10260
rect 147312 10140 147364 10192
rect 145196 10115 145248 10124
rect 145196 10081 145205 10115
rect 145205 10081 145239 10115
rect 145239 10081 145248 10115
rect 145196 10072 145248 10081
rect 146208 10072 146260 10124
rect 148600 10072 148652 10124
rect 149612 10115 149664 10124
rect 149612 10081 149621 10115
rect 149621 10081 149655 10115
rect 149655 10081 149664 10115
rect 149612 10072 149664 10081
rect 136272 9936 136324 9945
rect 136732 9936 136784 9988
rect 139768 9936 139820 9988
rect 136456 9868 136508 9920
rect 138204 9911 138256 9920
rect 138204 9877 138213 9911
rect 138213 9877 138247 9911
rect 138247 9877 138256 9911
rect 138204 9868 138256 9877
rect 138664 9868 138716 9920
rect 139860 9868 139912 9920
rect 140320 9868 140372 9920
rect 140780 9936 140832 9988
rect 142896 10004 142948 10056
rect 143448 10004 143500 10056
rect 141148 9911 141200 9920
rect 141148 9877 141157 9911
rect 141157 9877 141191 9911
rect 141191 9877 141200 9911
rect 141148 9868 141200 9877
rect 142160 9936 142212 9988
rect 144920 10004 144972 10056
rect 146024 10004 146076 10056
rect 147036 10004 147088 10056
rect 147220 10004 147272 10056
rect 144644 9936 144696 9988
rect 146116 9936 146168 9988
rect 148048 10004 148100 10056
rect 149336 10047 149388 10056
rect 149336 10013 149354 10047
rect 149354 10013 149388 10047
rect 149336 10004 149388 10013
rect 150256 10140 150308 10192
rect 150072 10072 150124 10124
rect 150440 10072 150492 10124
rect 153660 10140 153712 10192
rect 153844 10183 153896 10192
rect 153844 10149 153853 10183
rect 153853 10149 153887 10183
rect 153887 10149 153896 10183
rect 153844 10140 153896 10149
rect 144092 9868 144144 9920
rect 144276 9868 144328 9920
rect 144736 9911 144788 9920
rect 144736 9877 144745 9911
rect 144745 9877 144779 9911
rect 144779 9877 144788 9911
rect 144736 9868 144788 9877
rect 144828 9868 144880 9920
rect 145472 9868 145524 9920
rect 147864 9868 147916 9920
rect 153936 10072 153988 10124
rect 156236 10140 156288 10192
rect 150256 9936 150308 9988
rect 151360 9936 151412 9988
rect 152004 9936 152056 9988
rect 150072 9911 150124 9920
rect 150072 9877 150081 9911
rect 150081 9877 150115 9911
rect 150115 9877 150124 9911
rect 150072 9868 150124 9877
rect 150716 9868 150768 9920
rect 150900 9868 150952 9920
rect 151452 9868 151504 9920
rect 154672 10004 154724 10056
rect 155408 10072 155460 10124
rect 157708 10072 157760 10124
rect 152188 9868 152240 9920
rect 152280 9868 152332 9920
rect 154028 9868 154080 9920
rect 155776 10004 155828 10056
rect 155960 10004 156012 10056
rect 156604 10047 156656 10056
rect 156604 10013 156613 10047
rect 156613 10013 156647 10047
rect 156647 10013 156656 10047
rect 156604 10004 156656 10013
rect 157524 10047 157576 10056
rect 155408 9868 155460 9920
rect 157524 10013 157533 10047
rect 157533 10013 157567 10047
rect 157567 10013 157576 10047
rect 157524 10004 157576 10013
rect 157892 9868 157944 9920
rect 40394 9766 40446 9818
rect 40458 9766 40510 9818
rect 40522 9766 40574 9818
rect 40586 9766 40638 9818
rect 40650 9766 40702 9818
rect 79839 9766 79891 9818
rect 79903 9766 79955 9818
rect 79967 9766 80019 9818
rect 80031 9766 80083 9818
rect 80095 9766 80147 9818
rect 119284 9766 119336 9818
rect 119348 9766 119400 9818
rect 119412 9766 119464 9818
rect 119476 9766 119528 9818
rect 119540 9766 119592 9818
rect 158729 9766 158781 9818
rect 158793 9766 158845 9818
rect 158857 9766 158909 9818
rect 158921 9766 158973 9818
rect 158985 9766 159037 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 5172 9596 5224 9648
rect 29092 9664 29144 9716
rect 29460 9664 29512 9716
rect 10048 9596 10100 9648
rect 13452 9596 13504 9648
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 5724 9528 5776 9580
rect 12348 9528 12400 9580
rect 14280 9596 14332 9648
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 17776 9596 17828 9648
rect 14096 9528 14148 9580
rect 14188 9528 14240 9580
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16672 9528 16724 9580
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 19340 9596 19392 9648
rect 20536 9596 20588 9648
rect 23388 9596 23440 9648
rect 28632 9596 28684 9648
rect 30656 9596 30708 9648
rect 31300 9664 31352 9716
rect 31668 9707 31720 9716
rect 31668 9673 31677 9707
rect 31677 9673 31711 9707
rect 31711 9673 31720 9707
rect 31668 9664 31720 9673
rect 15016 9460 15068 9512
rect 19432 9528 19484 9580
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 26884 9528 26936 9580
rect 30748 9528 30800 9580
rect 32036 9596 32088 9648
rect 34244 9596 34296 9648
rect 35900 9664 35952 9716
rect 36728 9664 36780 9716
rect 38660 9664 38712 9716
rect 38568 9596 38620 9648
rect 19524 9460 19576 9512
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 26332 9503 26384 9512
rect 26332 9469 26341 9503
rect 26341 9469 26375 9503
rect 26375 9469 26384 9503
rect 26332 9460 26384 9469
rect 29092 9503 29144 9512
rect 8024 9324 8076 9376
rect 14464 9324 14516 9376
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 17500 9324 17552 9376
rect 19800 9392 19852 9444
rect 27068 9392 27120 9444
rect 19892 9324 19944 9376
rect 26516 9324 26568 9376
rect 27712 9324 27764 9376
rect 29092 9469 29101 9503
rect 29101 9469 29135 9503
rect 29135 9469 29144 9503
rect 29092 9460 29144 9469
rect 31024 9460 31076 9512
rect 33324 9528 33376 9580
rect 34520 9571 34572 9580
rect 34520 9537 34529 9571
rect 34529 9537 34563 9571
rect 34563 9537 34572 9571
rect 34520 9528 34572 9537
rect 39396 9596 39448 9648
rect 40224 9639 40276 9648
rect 33876 9460 33928 9512
rect 40224 9605 40233 9639
rect 40233 9605 40267 9639
rect 40267 9605 40276 9639
rect 40224 9596 40276 9605
rect 40960 9639 41012 9648
rect 40960 9605 40994 9639
rect 40994 9605 41012 9639
rect 40960 9596 41012 9605
rect 42892 9596 42944 9648
rect 45192 9664 45244 9716
rect 47124 9664 47176 9716
rect 47768 9664 47820 9716
rect 48228 9664 48280 9716
rect 49884 9664 49936 9716
rect 54208 9664 54260 9716
rect 48136 9596 48188 9648
rect 49700 9596 49752 9648
rect 40040 9460 40092 9512
rect 41512 9528 41564 9580
rect 41788 9528 41840 9580
rect 43076 9528 43128 9580
rect 46756 9528 46808 9580
rect 47032 9571 47084 9580
rect 47032 9537 47041 9571
rect 47041 9537 47075 9571
rect 47075 9537 47084 9571
rect 47032 9528 47084 9537
rect 47676 9528 47728 9580
rect 48596 9528 48648 9580
rect 48872 9528 48924 9580
rect 49792 9528 49844 9580
rect 43168 9503 43220 9512
rect 37556 9435 37608 9444
rect 30012 9324 30064 9376
rect 37556 9401 37565 9435
rect 37565 9401 37599 9435
rect 37599 9401 37608 9435
rect 37556 9392 37608 9401
rect 33048 9324 33100 9376
rect 33876 9324 33928 9376
rect 38568 9324 38620 9376
rect 38752 9324 38804 9376
rect 43168 9469 43177 9503
rect 43177 9469 43211 9503
rect 43211 9469 43220 9503
rect 43168 9460 43220 9469
rect 50620 9596 50672 9648
rect 50804 9596 50856 9648
rect 51448 9596 51500 9648
rect 53012 9528 53064 9580
rect 53472 9528 53524 9580
rect 53840 9596 53892 9648
rect 54484 9596 54536 9648
rect 56600 9664 56652 9716
rect 57060 9664 57112 9716
rect 61200 9664 61252 9716
rect 63040 9664 63092 9716
rect 64972 9664 65024 9716
rect 65248 9664 65300 9716
rect 54300 9528 54352 9580
rect 55496 9528 55548 9580
rect 56232 9528 56284 9580
rect 57152 9596 57204 9648
rect 58072 9596 58124 9648
rect 57520 9571 57572 9580
rect 57520 9537 57529 9571
rect 57529 9537 57563 9571
rect 57563 9537 57572 9571
rect 57520 9528 57572 9537
rect 57704 9528 57756 9580
rect 41880 9392 41932 9444
rect 40224 9324 40276 9376
rect 41972 9324 42024 9376
rect 43076 9324 43128 9376
rect 43904 9324 43956 9376
rect 44732 9392 44784 9444
rect 45192 9367 45244 9376
rect 45192 9333 45201 9367
rect 45201 9333 45235 9367
rect 45235 9333 45244 9367
rect 45192 9324 45244 9333
rect 45744 9367 45796 9376
rect 45744 9333 45753 9367
rect 45753 9333 45787 9367
rect 45787 9333 45796 9367
rect 45744 9324 45796 9333
rect 46296 9367 46348 9376
rect 46296 9333 46305 9367
rect 46305 9333 46339 9367
rect 46339 9333 46348 9367
rect 46296 9324 46348 9333
rect 46756 9324 46808 9376
rect 47308 9324 47360 9376
rect 48688 9324 48740 9376
rect 49240 9392 49292 9444
rect 49516 9392 49568 9444
rect 52828 9392 52880 9444
rect 51172 9324 51224 9376
rect 52184 9324 52236 9376
rect 56692 9460 56744 9512
rect 56876 9460 56928 9512
rect 60004 9528 60056 9580
rect 60740 9571 60792 9580
rect 60740 9537 60749 9571
rect 60749 9537 60783 9571
rect 60783 9537 60792 9571
rect 62120 9596 62172 9648
rect 60740 9528 60792 9537
rect 63500 9528 63552 9580
rect 64880 9571 64932 9580
rect 64880 9537 64889 9571
rect 64889 9537 64923 9571
rect 64923 9537 64932 9571
rect 64880 9528 64932 9537
rect 64972 9571 65024 9580
rect 64972 9537 64981 9571
rect 64981 9537 65015 9571
rect 65015 9537 65024 9571
rect 64972 9528 65024 9537
rect 63684 9460 63736 9512
rect 72608 9664 72660 9716
rect 73712 9664 73764 9716
rect 82728 9664 82780 9716
rect 88340 9707 88392 9716
rect 66904 9596 66956 9648
rect 71780 9596 71832 9648
rect 67456 9528 67508 9580
rect 73436 9596 73488 9648
rect 74724 9639 74776 9648
rect 73712 9571 73764 9580
rect 73712 9537 73721 9571
rect 73721 9537 73755 9571
rect 73755 9537 73764 9571
rect 73712 9528 73764 9537
rect 74724 9605 74733 9639
rect 74733 9605 74767 9639
rect 74767 9605 74776 9639
rect 74724 9596 74776 9605
rect 75920 9596 75972 9648
rect 76656 9596 76708 9648
rect 74448 9460 74500 9512
rect 76564 9503 76616 9512
rect 54208 9324 54260 9376
rect 56600 9392 56652 9444
rect 58440 9435 58492 9444
rect 58440 9401 58449 9435
rect 58449 9401 58483 9435
rect 58483 9401 58492 9435
rect 58440 9392 58492 9401
rect 66260 9392 66312 9444
rect 56416 9324 56468 9376
rect 58072 9324 58124 9376
rect 61660 9367 61712 9376
rect 61660 9333 61669 9367
rect 61669 9333 61703 9367
rect 61703 9333 61712 9367
rect 61660 9324 61712 9333
rect 63776 9367 63828 9376
rect 63776 9333 63785 9367
rect 63785 9333 63819 9367
rect 63819 9333 63828 9367
rect 63776 9324 63828 9333
rect 65800 9324 65852 9376
rect 66720 9324 66772 9376
rect 73528 9367 73580 9376
rect 73528 9333 73537 9367
rect 73537 9333 73571 9367
rect 73571 9333 73580 9367
rect 73528 9324 73580 9333
rect 76564 9469 76573 9503
rect 76573 9469 76607 9503
rect 76607 9469 76616 9503
rect 76564 9460 76616 9469
rect 79876 9596 79928 9648
rect 84844 9596 84896 9648
rect 85120 9596 85172 9648
rect 88340 9673 88349 9707
rect 88349 9673 88383 9707
rect 88383 9673 88392 9707
rect 88340 9664 88392 9673
rect 89076 9664 89128 9716
rect 79692 9528 79744 9580
rect 82544 9460 82596 9512
rect 83004 9460 83056 9512
rect 85396 9528 85448 9580
rect 88248 9528 88300 9580
rect 88340 9528 88392 9580
rect 90456 9596 90508 9648
rect 93860 9596 93912 9648
rect 95424 9664 95476 9716
rect 98092 9664 98144 9716
rect 95700 9596 95752 9648
rect 98736 9639 98788 9648
rect 77300 9392 77352 9444
rect 78680 9392 78732 9444
rect 79968 9392 80020 9444
rect 82268 9392 82320 9444
rect 90088 9460 90140 9512
rect 92296 9503 92348 9512
rect 85212 9392 85264 9444
rect 89076 9392 89128 9444
rect 79600 9324 79652 9376
rect 81440 9324 81492 9376
rect 82636 9324 82688 9376
rect 84200 9324 84252 9376
rect 84292 9324 84344 9376
rect 84476 9324 84528 9376
rect 90456 9367 90508 9376
rect 90456 9333 90465 9367
rect 90465 9333 90499 9367
rect 90499 9333 90508 9367
rect 90456 9324 90508 9333
rect 92296 9469 92305 9503
rect 92305 9469 92339 9503
rect 92339 9469 92348 9503
rect 92296 9460 92348 9469
rect 92940 9460 92992 9512
rect 98736 9605 98745 9639
rect 98745 9605 98779 9639
rect 98779 9605 98788 9639
rect 98736 9596 98788 9605
rect 98920 9664 98972 9716
rect 113548 9664 113600 9716
rect 113732 9664 113784 9716
rect 108028 9596 108080 9648
rect 92848 9324 92900 9376
rect 93860 9324 93912 9376
rect 94504 9324 94556 9376
rect 99380 9528 99432 9580
rect 104256 9528 104308 9580
rect 104440 9571 104492 9580
rect 104440 9537 104449 9571
rect 104449 9537 104483 9571
rect 104483 9537 104492 9571
rect 104440 9528 104492 9537
rect 104624 9571 104676 9580
rect 104624 9537 104633 9571
rect 104633 9537 104667 9571
rect 104667 9537 104676 9571
rect 104624 9528 104676 9537
rect 105636 9571 105688 9580
rect 105636 9537 105645 9571
rect 105645 9537 105679 9571
rect 105679 9537 105688 9571
rect 105636 9528 105688 9537
rect 105820 9528 105872 9580
rect 107844 9528 107896 9580
rect 110788 9528 110840 9580
rect 97356 9392 97408 9444
rect 107660 9460 107712 9512
rect 113824 9596 113876 9648
rect 116308 9596 116360 9648
rect 116584 9639 116636 9648
rect 116584 9605 116602 9639
rect 116602 9605 116636 9639
rect 117320 9664 117372 9716
rect 121000 9664 121052 9716
rect 130292 9639 130344 9648
rect 116584 9596 116636 9605
rect 113272 9503 113324 9512
rect 113272 9469 113281 9503
rect 113281 9469 113315 9503
rect 113315 9469 113324 9503
rect 113272 9460 113324 9469
rect 101220 9435 101272 9444
rect 101220 9401 101229 9435
rect 101229 9401 101263 9435
rect 101263 9401 101272 9435
rect 101220 9392 101272 9401
rect 108396 9392 108448 9444
rect 108672 9392 108724 9444
rect 113824 9460 113876 9512
rect 114744 9503 114796 9512
rect 114744 9469 114753 9503
rect 114753 9469 114787 9503
rect 114787 9469 114796 9503
rect 114744 9460 114796 9469
rect 115388 9460 115440 9512
rect 115848 9460 115900 9512
rect 117136 9460 117188 9512
rect 103244 9324 103296 9376
rect 103428 9367 103480 9376
rect 103428 9333 103437 9367
rect 103437 9333 103471 9367
rect 103471 9333 103480 9367
rect 103428 9324 103480 9333
rect 105360 9324 105412 9376
rect 105452 9367 105504 9376
rect 105452 9333 105461 9367
rect 105461 9333 105495 9367
rect 105495 9333 105504 9367
rect 107200 9367 107252 9376
rect 105452 9324 105504 9333
rect 107200 9333 107209 9367
rect 107209 9333 107243 9367
rect 107243 9333 107252 9367
rect 107200 9324 107252 9333
rect 107292 9324 107344 9376
rect 117964 9528 118016 9580
rect 121092 9528 121144 9580
rect 121920 9528 121972 9580
rect 124404 9571 124456 9580
rect 121736 9460 121788 9512
rect 124404 9537 124413 9571
rect 124413 9537 124447 9571
rect 124447 9537 124456 9571
rect 124404 9528 124456 9537
rect 127900 9528 127952 9580
rect 130292 9605 130301 9639
rect 130301 9605 130335 9639
rect 130335 9605 130344 9639
rect 130292 9596 130344 9605
rect 130936 9596 130988 9648
rect 133788 9664 133840 9716
rect 136916 9664 136968 9716
rect 125692 9503 125744 9512
rect 110052 9367 110104 9376
rect 110052 9333 110061 9367
rect 110061 9333 110095 9367
rect 110095 9333 110104 9367
rect 110052 9324 110104 9333
rect 110788 9324 110840 9376
rect 110972 9324 111024 9376
rect 111248 9324 111300 9376
rect 114008 9324 114060 9376
rect 114192 9324 114244 9376
rect 115388 9324 115440 9376
rect 117504 9324 117556 9376
rect 118332 9324 118384 9376
rect 119804 9324 119856 9376
rect 119988 9324 120040 9376
rect 121368 9324 121420 9376
rect 123300 9392 123352 9444
rect 125692 9469 125701 9503
rect 125701 9469 125735 9503
rect 125735 9469 125744 9503
rect 125692 9460 125744 9469
rect 125968 9460 126020 9512
rect 127532 9460 127584 9512
rect 130200 9460 130252 9512
rect 130292 9460 130344 9512
rect 137560 9596 137612 9648
rect 132592 9528 132644 9580
rect 133512 9528 133564 9580
rect 134064 9528 134116 9580
rect 134984 9528 135036 9580
rect 137468 9528 137520 9580
rect 133144 9460 133196 9512
rect 123852 9324 123904 9376
rect 125600 9324 125652 9376
rect 126152 9367 126204 9376
rect 126152 9333 126161 9367
rect 126161 9333 126195 9367
rect 126195 9333 126204 9367
rect 126152 9324 126204 9333
rect 126244 9324 126296 9376
rect 127072 9324 127124 9376
rect 128268 9367 128320 9376
rect 128268 9333 128277 9367
rect 128277 9333 128311 9367
rect 128311 9333 128320 9367
rect 128268 9324 128320 9333
rect 129648 9392 129700 9444
rect 131120 9392 131172 9444
rect 132224 9392 132276 9444
rect 132500 9324 132552 9376
rect 135536 9392 135588 9444
rect 136916 9392 136968 9444
rect 134800 9367 134852 9376
rect 134800 9333 134809 9367
rect 134809 9333 134843 9367
rect 134843 9333 134852 9367
rect 134800 9324 134852 9333
rect 137376 9367 137428 9376
rect 137376 9333 137385 9367
rect 137385 9333 137419 9367
rect 137419 9333 137428 9367
rect 139492 9596 139544 9648
rect 140596 9596 140648 9648
rect 143540 9664 143592 9716
rect 143908 9664 143960 9716
rect 147404 9664 147456 9716
rect 147956 9664 148008 9716
rect 149520 9664 149572 9716
rect 150992 9664 151044 9716
rect 151268 9707 151320 9716
rect 151268 9673 151277 9707
rect 151277 9673 151311 9707
rect 151311 9673 151320 9707
rect 151268 9664 151320 9673
rect 151728 9664 151780 9716
rect 158076 9664 158128 9716
rect 158260 9707 158312 9716
rect 158260 9673 158269 9707
rect 158269 9673 158303 9707
rect 158303 9673 158312 9707
rect 158260 9664 158312 9673
rect 140044 9528 140096 9580
rect 137376 9324 137428 9333
rect 137836 9324 137888 9376
rect 138940 9460 138992 9512
rect 139308 9435 139360 9444
rect 139308 9401 139317 9435
rect 139317 9401 139351 9435
rect 139351 9401 139360 9435
rect 139308 9392 139360 9401
rect 139492 9460 139544 9512
rect 141700 9460 141752 9512
rect 143448 9528 143500 9580
rect 143540 9528 143592 9580
rect 144368 9528 144420 9580
rect 145012 9528 145064 9580
rect 145472 9596 145524 9648
rect 149152 9596 149204 9648
rect 153936 9639 153988 9648
rect 153936 9605 153945 9639
rect 153945 9605 153979 9639
rect 153979 9605 153988 9639
rect 153936 9596 153988 9605
rect 147312 9528 147364 9580
rect 139860 9367 139912 9376
rect 139860 9333 139869 9367
rect 139869 9333 139903 9367
rect 139903 9333 139912 9367
rect 139860 9324 139912 9333
rect 140780 9367 140832 9376
rect 140780 9333 140789 9367
rect 140789 9333 140823 9367
rect 140823 9333 140832 9367
rect 140780 9324 140832 9333
rect 142160 9324 142212 9376
rect 143724 9367 143776 9376
rect 143724 9333 143733 9367
rect 143733 9333 143767 9367
rect 143767 9333 143776 9367
rect 143724 9324 143776 9333
rect 145196 9460 145248 9512
rect 145656 9460 145708 9512
rect 147128 9503 147180 9512
rect 147128 9469 147137 9503
rect 147137 9469 147171 9503
rect 147171 9469 147180 9503
rect 147128 9460 147180 9469
rect 149336 9528 149388 9580
rect 149520 9528 149572 9580
rect 150992 9528 151044 9580
rect 152096 9528 152148 9580
rect 152556 9528 152608 9580
rect 153292 9571 153344 9580
rect 153292 9537 153301 9571
rect 153301 9537 153335 9571
rect 153335 9537 153344 9571
rect 153292 9528 153344 9537
rect 153660 9528 153712 9580
rect 155316 9596 155368 9648
rect 151452 9460 151504 9512
rect 152648 9503 152700 9512
rect 152648 9469 152657 9503
rect 152657 9469 152691 9503
rect 152691 9469 152700 9503
rect 152648 9460 152700 9469
rect 153016 9460 153068 9512
rect 153476 9503 153528 9512
rect 153476 9469 153485 9503
rect 153485 9469 153519 9503
rect 153519 9469 153528 9503
rect 153476 9460 153528 9469
rect 149152 9392 149204 9444
rect 145564 9324 145616 9376
rect 145748 9367 145800 9376
rect 145748 9333 145757 9367
rect 145757 9333 145791 9367
rect 145791 9333 145800 9367
rect 145748 9324 145800 9333
rect 148876 9324 148928 9376
rect 149520 9324 149572 9376
rect 150532 9392 150584 9444
rect 151636 9392 151688 9444
rect 154672 9528 154724 9580
rect 155040 9571 155092 9580
rect 155040 9537 155049 9571
rect 155049 9537 155083 9571
rect 155083 9537 155092 9571
rect 155040 9528 155092 9537
rect 156144 9571 156196 9580
rect 156144 9537 156153 9571
rect 156153 9537 156187 9571
rect 156187 9537 156196 9571
rect 156144 9528 156196 9537
rect 156328 9528 156380 9580
rect 157800 9571 157852 9580
rect 157800 9537 157809 9571
rect 157809 9537 157843 9571
rect 157843 9537 157852 9571
rect 157800 9528 157852 9537
rect 154304 9503 154356 9512
rect 154304 9469 154313 9503
rect 154313 9469 154347 9503
rect 154347 9469 154356 9503
rect 154304 9460 154356 9469
rect 154764 9460 154816 9512
rect 155500 9460 155552 9512
rect 155868 9460 155920 9512
rect 154028 9392 154080 9444
rect 154120 9392 154172 9444
rect 152280 9324 152332 9376
rect 153108 9367 153160 9376
rect 153108 9333 153117 9367
rect 153117 9333 153151 9367
rect 153151 9333 153160 9367
rect 153108 9324 153160 9333
rect 153844 9324 153896 9376
rect 156972 9392 157024 9444
rect 156236 9324 156288 9376
rect 157064 9324 157116 9376
rect 157984 9392 158036 9444
rect 157524 9324 157576 9376
rect 20672 9222 20724 9274
rect 20736 9222 20788 9274
rect 20800 9222 20852 9274
rect 20864 9222 20916 9274
rect 20928 9222 20980 9274
rect 60117 9222 60169 9274
rect 60181 9222 60233 9274
rect 60245 9222 60297 9274
rect 60309 9222 60361 9274
rect 60373 9222 60425 9274
rect 99562 9222 99614 9274
rect 99626 9222 99678 9274
rect 99690 9222 99742 9274
rect 99754 9222 99806 9274
rect 99818 9222 99870 9274
rect 139007 9222 139059 9274
rect 139071 9222 139123 9274
rect 139135 9222 139187 9274
rect 139199 9222 139251 9274
rect 139263 9222 139315 9274
rect 11060 9120 11112 9172
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 12440 8916 12492 8968
rect 5264 8848 5316 8900
rect 17684 9120 17736 9172
rect 17776 9052 17828 9104
rect 18604 9095 18656 9104
rect 18604 9061 18613 9095
rect 18613 9061 18647 9095
rect 18647 9061 18656 9095
rect 18604 9052 18656 9061
rect 26332 9120 26384 9172
rect 26516 9120 26568 9172
rect 29736 9052 29788 9104
rect 38660 9120 38712 9172
rect 39396 9163 39448 9172
rect 39396 9129 39405 9163
rect 39405 9129 39439 9163
rect 39439 9129 39448 9163
rect 39396 9120 39448 9129
rect 13452 8984 13504 9036
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 15108 9027 15160 9036
rect 15108 8993 15117 9027
rect 15117 8993 15151 9027
rect 15151 8993 15160 9027
rect 15108 8984 15160 8993
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 17684 8984 17736 9036
rect 19432 9027 19484 9036
rect 16764 8916 16816 8968
rect 17776 8959 17828 8968
rect 12164 8780 12216 8832
rect 12348 8780 12400 8832
rect 14372 8780 14424 8832
rect 15660 8848 15712 8900
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 19432 8993 19441 9027
rect 19441 8993 19475 9027
rect 19475 8993 19484 9027
rect 19432 8984 19484 8993
rect 21180 8916 21232 8968
rect 17592 8848 17644 8900
rect 19340 8848 19392 8900
rect 27620 8984 27672 9036
rect 27712 8984 27764 9036
rect 31668 8984 31720 9036
rect 33232 8984 33284 9036
rect 33600 8984 33652 9036
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 16120 8780 16172 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 18052 8780 18104 8832
rect 18696 8780 18748 8832
rect 20996 8780 21048 8832
rect 26056 8780 26108 8832
rect 29092 8916 29144 8968
rect 30472 8916 30524 8968
rect 32864 8916 32916 8968
rect 32956 8916 33008 8968
rect 40224 9052 40276 9104
rect 36728 9027 36780 9036
rect 36728 8993 36737 9027
rect 36737 8993 36771 9027
rect 36771 8993 36780 9027
rect 44732 9120 44784 9172
rect 45468 9120 45520 9172
rect 47032 9052 47084 9104
rect 48320 9052 48372 9104
rect 49608 9120 49660 9172
rect 49700 9120 49752 9172
rect 53380 9163 53432 9172
rect 49424 9052 49476 9104
rect 49516 9052 49568 9104
rect 49884 9052 49936 9104
rect 53380 9129 53389 9163
rect 53389 9129 53423 9163
rect 53423 9129 53432 9163
rect 53380 9120 53432 9129
rect 36728 8984 36780 8993
rect 41052 8916 41104 8968
rect 41696 8916 41748 8968
rect 43168 8916 43220 8968
rect 43996 8916 44048 8968
rect 45560 8984 45612 9036
rect 47676 8984 47728 9036
rect 50344 8984 50396 9036
rect 54208 9052 54260 9104
rect 55864 9120 55916 9172
rect 56876 9120 56928 9172
rect 56968 9120 57020 9172
rect 59820 9120 59872 9172
rect 64880 9120 64932 9172
rect 64972 9120 65024 9172
rect 54024 8984 54076 9036
rect 57704 9052 57756 9104
rect 60648 9052 60700 9104
rect 63500 9052 63552 9104
rect 62120 9027 62172 9036
rect 45376 8916 45428 8968
rect 46664 8916 46716 8968
rect 48412 8916 48464 8968
rect 53380 8916 53432 8968
rect 53840 8916 53892 8968
rect 54116 8916 54168 8968
rect 54300 8959 54352 8968
rect 54300 8925 54309 8959
rect 54309 8925 54343 8959
rect 54343 8925 54352 8959
rect 54300 8916 54352 8925
rect 62120 8993 62129 9027
rect 62129 8993 62163 9027
rect 62163 8993 62172 9027
rect 62120 8984 62172 8993
rect 55404 8916 55456 8968
rect 57704 8959 57756 8968
rect 32404 8848 32456 8900
rect 33692 8848 33744 8900
rect 37280 8848 37332 8900
rect 40960 8848 41012 8900
rect 41512 8891 41564 8900
rect 41512 8857 41530 8891
rect 41530 8857 41564 8891
rect 41512 8848 41564 8857
rect 41880 8848 41932 8900
rect 33600 8823 33652 8832
rect 33600 8789 33609 8823
rect 33609 8789 33643 8823
rect 33643 8789 33652 8823
rect 33600 8780 33652 8789
rect 34152 8780 34204 8832
rect 38016 8780 38068 8832
rect 39764 8780 39816 8832
rect 40040 8780 40092 8832
rect 41052 8780 41104 8832
rect 44180 8780 44232 8832
rect 45468 8848 45520 8900
rect 45560 8848 45612 8900
rect 46388 8780 46440 8832
rect 47216 8780 47268 8832
rect 57704 8925 57713 8959
rect 57713 8925 57747 8959
rect 57747 8925 57756 8959
rect 57704 8916 57756 8925
rect 57796 8916 57848 8968
rect 57980 8959 58032 8968
rect 57980 8925 58014 8959
rect 58014 8925 58032 8959
rect 57980 8916 58032 8925
rect 61660 8916 61712 8968
rect 49240 8823 49292 8832
rect 49240 8789 49249 8823
rect 49249 8789 49283 8823
rect 49283 8789 49292 8823
rect 49240 8780 49292 8789
rect 49976 8780 50028 8832
rect 50068 8780 50120 8832
rect 50804 8780 50856 8832
rect 52736 8780 52788 8832
rect 53472 8780 53524 8832
rect 54576 8780 54628 8832
rect 54944 8780 54996 8832
rect 56416 8823 56468 8832
rect 56416 8789 56425 8823
rect 56425 8789 56459 8823
rect 56459 8789 56468 8823
rect 56416 8780 56468 8789
rect 58164 8848 58216 8900
rect 60832 8891 60884 8900
rect 60832 8857 60841 8891
rect 60841 8857 60875 8891
rect 60875 8857 60884 8891
rect 60832 8848 60884 8857
rect 61752 8848 61804 8900
rect 62672 8848 62724 8900
rect 65248 8916 65300 8968
rect 65800 8959 65852 8968
rect 65800 8925 65809 8959
rect 65809 8925 65843 8959
rect 65843 8925 65852 8959
rect 65800 8916 65852 8925
rect 65892 8916 65944 8968
rect 69020 9120 69072 9172
rect 75920 9120 75972 9172
rect 69756 9052 69808 9104
rect 82636 9120 82688 9172
rect 82728 9120 82780 9172
rect 83924 9052 83976 9104
rect 85396 9052 85448 9104
rect 88156 9120 88208 9172
rect 88340 9120 88392 9172
rect 90824 9120 90876 9172
rect 90916 9120 90968 9172
rect 101036 9120 101088 9172
rect 101220 9163 101272 9172
rect 101220 9129 101229 9163
rect 101229 9129 101263 9163
rect 101263 9129 101272 9163
rect 101220 9120 101272 9129
rect 103244 9120 103296 9172
rect 114468 9120 114520 9172
rect 114928 9163 114980 9172
rect 114928 9129 114937 9163
rect 114937 9129 114971 9163
rect 114971 9129 114980 9163
rect 114928 9120 114980 9129
rect 115572 9120 115624 9172
rect 115848 9120 115900 9172
rect 118332 9120 118384 9172
rect 128268 9120 128320 9172
rect 89628 9052 89680 9104
rect 71136 8984 71188 9036
rect 75184 8916 75236 8968
rect 69848 8848 69900 8900
rect 71688 8848 71740 8900
rect 75460 8984 75512 9036
rect 79692 8984 79744 9036
rect 75368 8916 75420 8968
rect 76656 8916 76708 8968
rect 84476 8984 84528 9036
rect 80336 8916 80388 8968
rect 86408 8959 86460 8968
rect 86408 8925 86417 8959
rect 86417 8925 86451 8959
rect 86451 8925 86460 8959
rect 86408 8916 86460 8925
rect 92940 9027 92992 9036
rect 92940 8993 92949 9027
rect 92949 8993 92983 9027
rect 92983 8993 92992 9027
rect 92940 8984 92992 8993
rect 89720 8916 89772 8968
rect 90916 8916 90968 8968
rect 95240 9052 95292 9104
rect 98092 9052 98144 9104
rect 99380 9052 99432 9104
rect 99748 9052 99800 9104
rect 95516 8984 95568 9036
rect 104440 9052 104492 9104
rect 107476 9052 107528 9104
rect 120724 9052 120776 9104
rect 121920 9052 121972 9104
rect 124220 9052 124272 9104
rect 126980 9095 127032 9104
rect 57336 8780 57388 8832
rect 57520 8780 57572 8832
rect 58256 8780 58308 8832
rect 59728 8780 59780 8832
rect 61292 8780 61344 8832
rect 61660 8823 61712 8832
rect 61660 8789 61669 8823
rect 61669 8789 61703 8823
rect 61703 8789 61712 8823
rect 61660 8780 61712 8789
rect 63592 8780 63644 8832
rect 65064 8780 65116 8832
rect 68376 8780 68428 8832
rect 73252 8780 73304 8832
rect 79968 8848 80020 8900
rect 86500 8848 86552 8900
rect 90456 8848 90508 8900
rect 90732 8848 90784 8900
rect 76012 8780 76064 8832
rect 76288 8780 76340 8832
rect 76380 8780 76432 8832
rect 84016 8780 84068 8832
rect 84292 8780 84344 8832
rect 87788 8780 87840 8832
rect 88340 8823 88392 8832
rect 88340 8789 88349 8823
rect 88349 8789 88383 8823
rect 88383 8789 88392 8823
rect 88340 8780 88392 8789
rect 89444 8823 89496 8832
rect 89444 8789 89453 8823
rect 89453 8789 89487 8823
rect 89487 8789 89496 8823
rect 89444 8780 89496 8789
rect 89628 8780 89680 8832
rect 92572 8848 92624 8900
rect 93676 8891 93728 8900
rect 93676 8857 93710 8891
rect 93710 8857 93728 8891
rect 93676 8848 93728 8857
rect 95424 8848 95476 8900
rect 104624 8984 104676 9036
rect 96160 8916 96212 8968
rect 97724 8848 97776 8900
rect 98000 8916 98052 8968
rect 99472 8916 99524 8968
rect 107200 8916 107252 8968
rect 107568 8959 107620 8968
rect 95056 8780 95108 8832
rect 97632 8780 97684 8832
rect 104624 8848 104676 8900
rect 107568 8925 107577 8959
rect 107577 8925 107611 8959
rect 107611 8925 107620 8959
rect 107568 8916 107620 8925
rect 111340 8916 111392 8968
rect 112352 8959 112404 8968
rect 112352 8925 112361 8959
rect 112361 8925 112395 8959
rect 112395 8925 112404 8959
rect 112352 8916 112404 8925
rect 118148 8959 118200 8968
rect 118148 8925 118157 8959
rect 118157 8925 118191 8959
rect 118191 8925 118200 8959
rect 118148 8916 118200 8925
rect 119620 8959 119672 8968
rect 119620 8925 119629 8959
rect 119629 8925 119663 8959
rect 119663 8925 119672 8959
rect 119620 8916 119672 8925
rect 107936 8848 107988 8900
rect 108948 8848 109000 8900
rect 109224 8848 109276 8900
rect 98184 8780 98236 8832
rect 99380 8823 99432 8832
rect 99380 8789 99389 8823
rect 99389 8789 99423 8823
rect 99423 8789 99432 8823
rect 108212 8823 108264 8832
rect 99380 8780 99432 8789
rect 108212 8789 108221 8823
rect 108221 8789 108255 8823
rect 108255 8789 108264 8823
rect 108212 8780 108264 8789
rect 110788 8780 110840 8832
rect 113272 8780 113324 8832
rect 115848 8780 115900 8832
rect 117228 8848 117280 8900
rect 118424 8848 118476 8900
rect 116952 8780 117004 8832
rect 117136 8780 117188 8832
rect 118976 8780 119028 8832
rect 119160 8780 119212 8832
rect 120908 8916 120960 8968
rect 121828 8959 121880 8968
rect 121828 8925 121837 8959
rect 121837 8925 121871 8959
rect 121871 8925 121880 8959
rect 121828 8916 121880 8925
rect 120448 8848 120500 8900
rect 120264 8780 120316 8832
rect 121368 8823 121420 8832
rect 121368 8789 121377 8823
rect 121377 8789 121411 8823
rect 121411 8789 121420 8823
rect 121368 8780 121420 8789
rect 122380 8780 122432 8832
rect 122472 8823 122524 8832
rect 122472 8789 122481 8823
rect 122481 8789 122515 8823
rect 122515 8789 122524 8823
rect 126612 9027 126664 9036
rect 126612 8993 126621 9027
rect 126621 8993 126655 9027
rect 126655 8993 126664 9027
rect 126980 9061 126989 9095
rect 126989 9061 127023 9095
rect 127023 9061 127032 9095
rect 126980 9052 127032 9061
rect 129096 9052 129148 9104
rect 126612 8984 126664 8993
rect 127532 8984 127584 9036
rect 130936 9120 130988 9172
rect 131028 9120 131080 9172
rect 130844 9052 130896 9104
rect 131120 9095 131172 9104
rect 131120 9061 131129 9095
rect 131129 9061 131163 9095
rect 131163 9061 131172 9095
rect 131120 9052 131172 9061
rect 131948 9120 132000 9172
rect 134800 9120 134852 9172
rect 135076 9120 135128 9172
rect 136456 9120 136508 9172
rect 136548 9120 136600 9172
rect 137836 9120 137888 9172
rect 132500 9052 132552 9104
rect 137928 9052 137980 9104
rect 138204 9120 138256 9172
rect 145748 9120 145800 9172
rect 146024 9120 146076 9172
rect 138664 9095 138716 9104
rect 138664 9061 138673 9095
rect 138673 9061 138707 9095
rect 138707 9061 138716 9095
rect 138664 9052 138716 9061
rect 139492 9052 139544 9104
rect 139768 9052 139820 9104
rect 140596 9052 140648 9104
rect 140688 9052 140740 9104
rect 143448 9052 143500 9104
rect 144644 9052 144696 9104
rect 145104 9052 145156 9104
rect 145472 9052 145524 9104
rect 147220 9052 147272 9104
rect 148600 9052 148652 9104
rect 123760 8916 123812 8968
rect 128820 8916 128872 8968
rect 131672 8916 131724 8968
rect 122472 8780 122524 8789
rect 123852 8780 123904 8832
rect 124404 8780 124456 8832
rect 125416 8780 125468 8832
rect 125692 8780 125744 8832
rect 126244 8780 126296 8832
rect 127716 8780 127768 8832
rect 128544 8780 128596 8832
rect 129556 8848 129608 8900
rect 130292 8848 130344 8900
rect 137376 8984 137428 9036
rect 137560 8984 137612 9036
rect 139584 8984 139636 9036
rect 133512 8916 133564 8968
rect 133696 8916 133748 8968
rect 135076 8916 135128 8968
rect 135260 8916 135312 8968
rect 135996 8916 136048 8968
rect 136456 8916 136508 8968
rect 138664 8916 138716 8968
rect 140964 8959 141016 8968
rect 140964 8925 140973 8959
rect 140973 8925 141007 8959
rect 141007 8925 141016 8959
rect 140964 8916 141016 8925
rect 141516 8916 141568 8968
rect 141976 8959 142028 8968
rect 141976 8925 141985 8959
rect 141985 8925 142019 8959
rect 142019 8925 142028 8959
rect 141976 8916 142028 8925
rect 143632 8916 143684 8968
rect 145840 8984 145892 9036
rect 147128 8984 147180 9036
rect 147496 8984 147548 9036
rect 144644 8916 144696 8968
rect 144828 8916 144880 8968
rect 145012 8916 145064 8968
rect 147404 8916 147456 8968
rect 148232 8984 148284 9036
rect 132132 8891 132184 8900
rect 132132 8857 132141 8891
rect 132141 8857 132175 8891
rect 132175 8857 132184 8891
rect 132132 8848 132184 8857
rect 130844 8780 130896 8832
rect 137376 8848 137428 8900
rect 132868 8780 132920 8832
rect 133512 8780 133564 8832
rect 133788 8780 133840 8832
rect 135260 8780 135312 8832
rect 135536 8780 135588 8832
rect 135996 8780 136048 8832
rect 136456 8823 136508 8832
rect 136456 8789 136465 8823
rect 136465 8789 136499 8823
rect 136499 8789 136508 8823
rect 136456 8780 136508 8789
rect 136916 8780 136968 8832
rect 137468 8780 137520 8832
rect 139676 8780 139728 8832
rect 140596 8780 140648 8832
rect 141332 8848 141384 8900
rect 142896 8780 142948 8832
rect 143080 8823 143132 8832
rect 143080 8789 143089 8823
rect 143089 8789 143123 8823
rect 143123 8789 143132 8823
rect 143080 8780 143132 8789
rect 144552 8780 144604 8832
rect 145932 8780 145984 8832
rect 147128 8848 147180 8900
rect 147496 8823 147548 8832
rect 147496 8789 147505 8823
rect 147505 8789 147539 8823
rect 147539 8789 147548 8823
rect 148324 8823 148376 8832
rect 147496 8780 147548 8789
rect 148324 8789 148333 8823
rect 148333 8789 148367 8823
rect 148367 8789 148376 8823
rect 148324 8780 148376 8789
rect 148784 9163 148836 9172
rect 148784 9129 148793 9163
rect 148793 9129 148827 9163
rect 148827 9129 148836 9163
rect 148784 9120 148836 9129
rect 148876 9052 148928 9104
rect 150440 9052 150492 9104
rect 151820 9052 151872 9104
rect 152832 9052 152884 9104
rect 153568 9120 153620 9172
rect 154672 9120 154724 9172
rect 157800 9120 157852 9172
rect 153660 9052 153712 9104
rect 154764 9052 154816 9104
rect 156880 9052 156932 9104
rect 149612 8916 149664 8968
rect 150256 8916 150308 8968
rect 152004 8984 152056 9036
rect 150900 8848 150952 8900
rect 150532 8780 150584 8832
rect 150992 8823 151044 8832
rect 150992 8789 151001 8823
rect 151001 8789 151035 8823
rect 151035 8789 151044 8823
rect 150992 8780 151044 8789
rect 151636 8959 151688 8968
rect 151636 8925 151645 8959
rect 151645 8925 151679 8959
rect 151679 8925 151688 8959
rect 151636 8916 151688 8925
rect 152096 8916 152148 8968
rect 152464 8959 152516 8968
rect 152464 8925 152473 8959
rect 152473 8925 152507 8959
rect 152507 8925 152516 8959
rect 152464 8916 152516 8925
rect 152556 8959 152608 8968
rect 152556 8925 152565 8959
rect 152565 8925 152599 8959
rect 152599 8925 152608 8959
rect 153476 8959 153528 8968
rect 152556 8916 152608 8925
rect 153476 8925 153485 8959
rect 153485 8925 153519 8959
rect 153519 8925 153528 8959
rect 153476 8916 153528 8925
rect 155040 8984 155092 9036
rect 153936 8916 153988 8968
rect 154212 8959 154264 8968
rect 154212 8925 154221 8959
rect 154221 8925 154255 8959
rect 154255 8925 154264 8959
rect 154212 8916 154264 8925
rect 155960 8984 156012 9036
rect 151728 8848 151780 8900
rect 153660 8848 153712 8900
rect 152832 8780 152884 8832
rect 155224 8959 155276 8968
rect 155224 8925 155233 8959
rect 155233 8925 155267 8959
rect 155267 8925 155276 8959
rect 156052 8959 156104 8968
rect 155224 8916 155276 8925
rect 156052 8925 156061 8959
rect 156061 8925 156095 8959
rect 156095 8925 156104 8959
rect 156052 8916 156104 8925
rect 156144 8959 156196 8968
rect 156144 8925 156153 8959
rect 156153 8925 156187 8959
rect 156187 8925 156196 8959
rect 156144 8916 156196 8925
rect 156328 8916 156380 8968
rect 156788 8916 156840 8968
rect 157708 8959 157760 8968
rect 157708 8925 157717 8959
rect 157717 8925 157751 8959
rect 157751 8925 157760 8959
rect 157708 8916 157760 8925
rect 158536 8848 158588 8900
rect 155040 8780 155092 8832
rect 156880 8780 156932 8832
rect 40394 8678 40446 8730
rect 40458 8678 40510 8730
rect 40522 8678 40574 8730
rect 40586 8678 40638 8730
rect 40650 8678 40702 8730
rect 79839 8678 79891 8730
rect 79903 8678 79955 8730
rect 79967 8678 80019 8730
rect 80031 8678 80083 8730
rect 80095 8678 80147 8730
rect 119284 8678 119336 8730
rect 119348 8678 119400 8730
rect 119412 8678 119464 8730
rect 119476 8678 119528 8730
rect 119540 8678 119592 8730
rect 158729 8678 158781 8730
rect 158793 8678 158845 8730
rect 158857 8678 158909 8730
rect 158921 8678 158973 8730
rect 158985 8678 159037 8730
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5816 8576 5868 8628
rect 12440 8576 12492 8628
rect 12900 8576 12952 8628
rect 13268 8508 13320 8560
rect 5540 8440 5592 8492
rect 18236 8576 18288 8628
rect 18696 8576 18748 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 28540 8619 28592 8628
rect 28540 8585 28549 8619
rect 28549 8585 28583 8619
rect 28583 8585 28592 8619
rect 28540 8576 28592 8585
rect 29552 8619 29604 8628
rect 29552 8585 29561 8619
rect 29561 8585 29595 8619
rect 29595 8585 29604 8619
rect 29552 8576 29604 8585
rect 29644 8576 29696 8628
rect 33324 8619 33376 8628
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 14924 8483 14976 8492
rect 14924 8449 14958 8483
rect 14958 8449 14976 8483
rect 14924 8440 14976 8449
rect 16488 8440 16540 8492
rect 17684 8440 17736 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18236 8440 18288 8492
rect 5632 8372 5684 8424
rect 5356 8304 5408 8356
rect 6736 8304 6788 8356
rect 5080 8236 5132 8288
rect 8208 8304 8260 8356
rect 11980 8304 12032 8356
rect 16764 8372 16816 8424
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 19800 8372 19852 8424
rect 19984 8372 20036 8424
rect 26332 8440 26384 8492
rect 29092 8508 29144 8560
rect 31024 8508 31076 8560
rect 33324 8585 33333 8619
rect 33333 8585 33367 8619
rect 33367 8585 33376 8619
rect 33324 8576 33376 8585
rect 34244 8576 34296 8628
rect 35256 8576 35308 8628
rect 35900 8619 35952 8628
rect 35900 8585 35909 8619
rect 35909 8585 35943 8619
rect 35943 8585 35952 8619
rect 35900 8576 35952 8585
rect 41052 8576 41104 8628
rect 41788 8576 41840 8628
rect 45468 8576 45520 8628
rect 45652 8576 45704 8628
rect 45928 8576 45980 8628
rect 27252 8440 27304 8492
rect 27712 8440 27764 8492
rect 30472 8440 30524 8492
rect 30840 8473 30892 8476
rect 30840 8439 30852 8473
rect 30852 8439 30886 8473
rect 30886 8439 30892 8473
rect 30840 8424 30892 8439
rect 33140 8440 33192 8492
rect 16488 8304 16540 8356
rect 17776 8304 17828 8356
rect 21916 8304 21968 8356
rect 27068 8304 27120 8356
rect 8668 8236 8720 8288
rect 10692 8236 10744 8288
rect 14280 8236 14332 8288
rect 15752 8236 15804 8288
rect 16948 8236 17000 8288
rect 17316 8236 17368 8288
rect 18972 8236 19024 8288
rect 24216 8236 24268 8288
rect 28172 8372 28224 8424
rect 29644 8372 29696 8424
rect 30564 8372 30616 8424
rect 31116 8372 31168 8424
rect 35256 8440 35308 8492
rect 36544 8483 36596 8492
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 37648 8508 37700 8560
rect 38476 8508 38528 8560
rect 38936 8551 38988 8560
rect 38936 8517 38970 8551
rect 38970 8517 38988 8551
rect 38936 8508 38988 8517
rect 39396 8508 39448 8560
rect 49424 8619 49476 8628
rect 49424 8585 49433 8619
rect 49433 8585 49467 8619
rect 49467 8585 49476 8619
rect 49424 8576 49476 8585
rect 51448 8619 51500 8628
rect 51448 8585 51457 8619
rect 51457 8585 51491 8619
rect 51491 8585 51500 8619
rect 51448 8576 51500 8585
rect 56140 8576 56192 8628
rect 60004 8619 60056 8628
rect 60004 8585 60013 8619
rect 60013 8585 60047 8619
rect 60047 8585 60056 8619
rect 60004 8576 60056 8585
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 38660 8483 38712 8492
rect 38660 8449 38669 8483
rect 38669 8449 38703 8483
rect 38703 8449 38712 8483
rect 38660 8440 38712 8449
rect 37004 8372 37056 8424
rect 31392 8236 31444 8288
rect 36544 8304 36596 8356
rect 32956 8236 33008 8288
rect 39304 8236 39356 8288
rect 41144 8440 41196 8492
rect 46388 8551 46440 8560
rect 46388 8517 46406 8551
rect 46406 8517 46440 8551
rect 46388 8508 46440 8517
rect 40776 8304 40828 8356
rect 41236 8304 41288 8356
rect 44180 8440 44232 8492
rect 44732 8440 44784 8492
rect 48872 8440 48924 8492
rect 50436 8508 50488 8560
rect 53380 8508 53432 8560
rect 55220 8508 55272 8560
rect 58072 8508 58124 8560
rect 60832 8508 60884 8560
rect 49148 8440 49200 8492
rect 52184 8483 52236 8492
rect 52184 8449 52193 8483
rect 52193 8449 52227 8483
rect 52227 8449 52236 8483
rect 52184 8440 52236 8449
rect 52276 8483 52328 8492
rect 52276 8449 52285 8483
rect 52285 8449 52319 8483
rect 52319 8449 52328 8483
rect 52276 8440 52328 8449
rect 52552 8440 52604 8492
rect 55680 8440 55732 8492
rect 57336 8483 57388 8492
rect 57336 8449 57345 8483
rect 57345 8449 57379 8483
rect 57379 8449 57388 8483
rect 57336 8440 57388 8449
rect 43996 8415 44048 8424
rect 43996 8381 44005 8415
rect 44005 8381 44039 8415
rect 44039 8381 44048 8415
rect 43996 8372 44048 8381
rect 45376 8372 45428 8424
rect 46664 8415 46716 8424
rect 46664 8381 46673 8415
rect 46673 8381 46707 8415
rect 46707 8381 46716 8415
rect 46664 8372 46716 8381
rect 49792 8372 49844 8424
rect 51080 8372 51132 8424
rect 51356 8372 51408 8424
rect 52092 8372 52144 8424
rect 52736 8372 52788 8424
rect 54116 8372 54168 8424
rect 59820 8440 59872 8492
rect 60648 8483 60700 8492
rect 60648 8449 60657 8483
rect 60657 8449 60691 8483
rect 60691 8449 60700 8483
rect 60648 8440 60700 8449
rect 62212 8576 62264 8628
rect 62672 8619 62724 8628
rect 62672 8585 62681 8619
rect 62681 8585 62715 8619
rect 62715 8585 62724 8619
rect 62672 8576 62724 8585
rect 65156 8576 65208 8628
rect 67456 8619 67508 8628
rect 67456 8585 67465 8619
rect 67465 8585 67499 8619
rect 67499 8585 67508 8619
rect 67456 8576 67508 8585
rect 69756 8619 69808 8628
rect 69756 8585 69765 8619
rect 69765 8585 69799 8619
rect 69799 8585 69808 8619
rect 69756 8576 69808 8585
rect 69848 8576 69900 8628
rect 83924 8576 83976 8628
rect 84016 8576 84068 8628
rect 64236 8551 64288 8560
rect 64236 8517 64245 8551
rect 64245 8517 64279 8551
rect 64279 8517 64288 8551
rect 64236 8508 64288 8517
rect 42064 8304 42116 8356
rect 44088 8304 44140 8356
rect 50988 8304 51040 8356
rect 53932 8347 53984 8356
rect 53932 8313 53941 8347
rect 53941 8313 53975 8347
rect 53975 8313 53984 8347
rect 53932 8304 53984 8313
rect 41788 8236 41840 8288
rect 42340 8236 42392 8288
rect 46020 8236 46072 8288
rect 46756 8236 46808 8288
rect 47032 8236 47084 8288
rect 51908 8236 51960 8288
rect 54208 8236 54260 8288
rect 54576 8236 54628 8288
rect 57520 8415 57572 8424
rect 57520 8381 57529 8415
rect 57529 8381 57563 8415
rect 57563 8381 57572 8415
rect 57520 8372 57572 8381
rect 56048 8304 56100 8356
rect 59728 8372 59780 8424
rect 85212 8508 85264 8560
rect 87880 8551 87932 8560
rect 87880 8517 87898 8551
rect 87898 8517 87932 8551
rect 89352 8576 89404 8628
rect 89444 8576 89496 8628
rect 117320 8576 117372 8628
rect 117504 8576 117556 8628
rect 121920 8576 121972 8628
rect 87880 8508 87932 8517
rect 90916 8508 90968 8560
rect 92480 8508 92532 8560
rect 108672 8508 108724 8560
rect 67640 8483 67692 8492
rect 67640 8449 67649 8483
rect 67649 8449 67683 8483
rect 67683 8449 67692 8483
rect 67640 8440 67692 8449
rect 70216 8483 70268 8492
rect 70216 8449 70225 8483
rect 70225 8449 70259 8483
rect 70259 8449 70268 8483
rect 70216 8440 70268 8449
rect 72332 8440 72384 8492
rect 76472 8440 76524 8492
rect 76564 8440 76616 8492
rect 83648 8440 83700 8492
rect 83832 8483 83884 8492
rect 83832 8449 83841 8483
rect 83841 8449 83875 8483
rect 83875 8449 83884 8483
rect 83832 8440 83884 8449
rect 67824 8415 67876 8424
rect 67824 8381 67833 8415
rect 67833 8381 67867 8415
rect 67867 8381 67876 8415
rect 67824 8372 67876 8381
rect 68376 8415 68428 8424
rect 68376 8381 68385 8415
rect 68385 8381 68419 8415
rect 68419 8381 68428 8415
rect 68376 8372 68428 8381
rect 73344 8372 73396 8424
rect 65892 8304 65944 8356
rect 73160 8304 73212 8356
rect 78864 8304 78916 8356
rect 80336 8304 80388 8356
rect 88432 8440 88484 8492
rect 90088 8483 90140 8492
rect 90088 8449 90106 8483
rect 90106 8449 90140 8483
rect 90088 8440 90140 8449
rect 90456 8440 90508 8492
rect 91008 8440 91060 8492
rect 91928 8483 91980 8492
rect 91928 8449 91946 8483
rect 91946 8449 91980 8483
rect 91928 8440 91980 8449
rect 92204 8483 92256 8492
rect 92204 8449 92206 8483
rect 92206 8449 92240 8483
rect 92240 8449 92256 8483
rect 92204 8440 92256 8449
rect 92388 8440 92440 8492
rect 88892 8372 88944 8424
rect 90364 8415 90416 8424
rect 90364 8381 90373 8415
rect 90373 8381 90407 8415
rect 90407 8381 90416 8415
rect 90364 8372 90416 8381
rect 90916 8372 90968 8424
rect 92296 8372 92348 8424
rect 94044 8372 94096 8424
rect 94320 8483 94372 8492
rect 94320 8449 94329 8483
rect 94329 8449 94363 8483
rect 94363 8449 94372 8483
rect 98184 8483 98236 8492
rect 94320 8440 94372 8449
rect 98184 8449 98193 8483
rect 98193 8449 98227 8483
rect 98227 8449 98236 8483
rect 98184 8440 98236 8449
rect 100392 8372 100444 8424
rect 101036 8440 101088 8492
rect 107568 8440 107620 8492
rect 107936 8440 107988 8492
rect 108488 8440 108540 8492
rect 109132 8440 109184 8492
rect 109592 8483 109644 8492
rect 109592 8449 109601 8483
rect 109601 8449 109635 8483
rect 109635 8449 109644 8483
rect 109592 8440 109644 8449
rect 107292 8372 107344 8424
rect 107384 8372 107436 8424
rect 112352 8508 112404 8560
rect 115296 8551 115348 8560
rect 115296 8517 115305 8551
rect 115305 8517 115339 8551
rect 115339 8517 115348 8551
rect 115296 8508 115348 8517
rect 112720 8440 112772 8492
rect 115572 8440 115624 8492
rect 114192 8372 114244 8424
rect 116676 8372 116728 8424
rect 117320 8440 117372 8492
rect 118976 8483 119028 8492
rect 118976 8449 118985 8483
rect 118985 8449 119019 8483
rect 119019 8449 119028 8483
rect 118976 8440 119028 8449
rect 122840 8440 122892 8492
rect 117504 8372 117556 8424
rect 117596 8372 117648 8424
rect 118332 8415 118384 8424
rect 118332 8381 118341 8415
rect 118341 8381 118375 8415
rect 118375 8381 118384 8415
rect 118332 8372 118384 8381
rect 118516 8372 118568 8424
rect 119160 8415 119212 8424
rect 119160 8381 119169 8415
rect 119169 8381 119203 8415
rect 119203 8381 119212 8415
rect 119160 8372 119212 8381
rect 119988 8372 120040 8424
rect 130292 8508 130344 8560
rect 123300 8483 123352 8492
rect 123300 8449 123334 8483
rect 123334 8449 123352 8483
rect 123300 8440 123352 8449
rect 123576 8440 123628 8492
rect 126612 8440 126664 8492
rect 127256 8483 127308 8492
rect 127256 8449 127265 8483
rect 127265 8449 127299 8483
rect 127299 8449 127308 8483
rect 127256 8440 127308 8449
rect 127348 8440 127400 8492
rect 86500 8304 86552 8356
rect 92204 8304 92256 8356
rect 93308 8347 93360 8356
rect 59084 8236 59136 8288
rect 60004 8236 60056 8288
rect 65248 8236 65300 8288
rect 74356 8279 74408 8288
rect 74356 8245 74365 8279
rect 74365 8245 74399 8279
rect 74399 8245 74408 8279
rect 74356 8236 74408 8245
rect 75092 8236 75144 8288
rect 83924 8236 83976 8288
rect 84108 8236 84160 8288
rect 90732 8236 90784 8288
rect 90824 8279 90876 8288
rect 90824 8245 90833 8279
rect 90833 8245 90867 8279
rect 90867 8245 90876 8279
rect 90824 8236 90876 8245
rect 92388 8236 92440 8288
rect 93308 8313 93317 8347
rect 93317 8313 93351 8347
rect 93351 8313 93360 8347
rect 93308 8304 93360 8313
rect 95332 8304 95384 8356
rect 95424 8304 95476 8356
rect 101680 8304 101732 8356
rect 104256 8304 104308 8356
rect 112812 8304 112864 8356
rect 97540 8236 97592 8288
rect 98276 8236 98328 8288
rect 101864 8236 101916 8288
rect 108672 8236 108724 8288
rect 112076 8236 112128 8288
rect 115940 8236 115992 8288
rect 116032 8236 116084 8288
rect 117504 8236 117556 8288
rect 119436 8304 119488 8356
rect 123024 8415 123076 8424
rect 123024 8381 123033 8415
rect 123033 8381 123067 8415
rect 123067 8381 123076 8415
rect 125140 8415 125192 8424
rect 123024 8372 123076 8381
rect 120172 8236 120224 8288
rect 122012 8304 122064 8356
rect 125140 8381 125149 8415
rect 125149 8381 125183 8415
rect 125183 8381 125192 8415
rect 125140 8372 125192 8381
rect 126152 8372 126204 8424
rect 126796 8415 126848 8424
rect 126796 8381 126805 8415
rect 126805 8381 126839 8415
rect 126839 8381 126848 8415
rect 126796 8372 126848 8381
rect 127624 8372 127676 8424
rect 131304 8576 131356 8628
rect 131672 8576 131724 8628
rect 132316 8576 132368 8628
rect 132776 8576 132828 8628
rect 143356 8576 143408 8628
rect 144920 8576 144972 8628
rect 146024 8576 146076 8628
rect 147772 8576 147824 8628
rect 132408 8440 132460 8492
rect 135352 8440 135404 8492
rect 135720 8440 135772 8492
rect 137836 8440 137888 8492
rect 138204 8440 138256 8492
rect 121460 8236 121512 8288
rect 123300 8236 123352 8288
rect 127716 8304 127768 8356
rect 128360 8304 128412 8356
rect 128452 8304 128504 8356
rect 133144 8372 133196 8424
rect 130292 8304 130344 8356
rect 131948 8304 132000 8356
rect 124128 8236 124180 8288
rect 129648 8236 129700 8288
rect 130660 8236 130712 8288
rect 131304 8236 131356 8288
rect 134708 8372 134760 8424
rect 136916 8415 136968 8424
rect 133788 8236 133840 8288
rect 134064 8236 134116 8288
rect 136916 8381 136925 8415
rect 136925 8381 136959 8415
rect 136959 8381 136968 8415
rect 136916 8372 136968 8381
rect 137192 8372 137244 8424
rect 135720 8304 135772 8356
rect 138572 8347 138624 8356
rect 138572 8313 138581 8347
rect 138581 8313 138615 8347
rect 138615 8313 138624 8347
rect 138572 8304 138624 8313
rect 139860 8372 139912 8424
rect 140964 8372 141016 8424
rect 140688 8347 140740 8356
rect 137468 8236 137520 8288
rect 138664 8236 138716 8288
rect 139768 8236 139820 8288
rect 140688 8313 140697 8347
rect 140697 8313 140731 8347
rect 140731 8313 140740 8347
rect 140688 8304 140740 8313
rect 140596 8236 140648 8288
rect 141332 8483 141384 8492
rect 141332 8449 141341 8483
rect 141341 8449 141375 8483
rect 141375 8449 141384 8483
rect 141332 8440 141384 8449
rect 141516 8440 141568 8492
rect 143080 8440 143132 8492
rect 143264 8440 143316 8492
rect 143908 8483 143960 8492
rect 143908 8449 143942 8483
rect 143942 8449 143960 8483
rect 143908 8440 143960 8449
rect 145656 8483 145708 8492
rect 145656 8449 145665 8483
rect 145665 8449 145699 8483
rect 145699 8449 145708 8483
rect 145656 8440 145708 8449
rect 147404 8440 147456 8492
rect 148232 8508 148284 8560
rect 148324 8508 148376 8560
rect 148692 8508 148744 8560
rect 149888 8576 149940 8628
rect 150808 8619 150860 8628
rect 150808 8585 150817 8619
rect 150817 8585 150851 8619
rect 150851 8585 150860 8619
rect 150808 8576 150860 8585
rect 150900 8576 150952 8628
rect 151084 8576 151136 8628
rect 155316 8619 155368 8628
rect 151636 8508 151688 8560
rect 141608 8372 141660 8424
rect 141976 8372 142028 8424
rect 144920 8372 144972 8424
rect 145564 8372 145616 8424
rect 147128 8372 147180 8424
rect 148968 8372 149020 8424
rect 149520 8483 149572 8492
rect 149520 8449 149529 8483
rect 149529 8449 149563 8483
rect 149563 8449 149572 8483
rect 149520 8440 149572 8449
rect 149888 8440 149940 8492
rect 151176 8440 151228 8492
rect 153752 8508 153804 8560
rect 151820 8440 151872 8492
rect 152832 8483 152884 8492
rect 152832 8449 152841 8483
rect 152841 8449 152875 8483
rect 152875 8449 152884 8483
rect 152832 8440 152884 8449
rect 141792 8347 141844 8356
rect 141792 8313 141801 8347
rect 141801 8313 141835 8347
rect 141835 8313 141844 8347
rect 141792 8304 141844 8313
rect 147220 8304 147272 8356
rect 147404 8304 147456 8356
rect 149060 8304 149112 8356
rect 150164 8372 150216 8424
rect 150900 8372 150952 8424
rect 152004 8415 152056 8424
rect 152004 8381 152013 8415
rect 152013 8381 152047 8415
rect 152047 8381 152056 8415
rect 152004 8372 152056 8381
rect 152280 8415 152332 8424
rect 152280 8381 152289 8415
rect 152289 8381 152323 8415
rect 152323 8381 152332 8415
rect 152280 8372 152332 8381
rect 142068 8236 142120 8288
rect 144920 8236 144972 8288
rect 146024 8236 146076 8288
rect 149428 8236 149480 8288
rect 153016 8304 153068 8356
rect 151084 8236 151136 8288
rect 153476 8236 153528 8288
rect 153660 8279 153712 8288
rect 153660 8245 153669 8279
rect 153669 8245 153703 8279
rect 153703 8245 153712 8279
rect 153660 8236 153712 8245
rect 154212 8508 154264 8560
rect 155316 8585 155325 8619
rect 155325 8585 155359 8619
rect 155359 8585 155368 8619
rect 155316 8576 155368 8585
rect 155960 8576 156012 8628
rect 156788 8576 156840 8628
rect 156972 8576 157024 8628
rect 154304 8440 154356 8492
rect 156788 8483 156840 8492
rect 154212 8372 154264 8424
rect 154488 8347 154540 8356
rect 154488 8313 154497 8347
rect 154497 8313 154531 8347
rect 154531 8313 154540 8347
rect 154488 8304 154540 8313
rect 154764 8372 154816 8424
rect 155776 8372 155828 8424
rect 156788 8449 156797 8483
rect 156797 8449 156831 8483
rect 156831 8449 156840 8483
rect 156788 8440 156840 8449
rect 156972 8483 157024 8492
rect 156972 8449 156981 8483
rect 156981 8449 157015 8483
rect 157015 8449 157024 8483
rect 156972 8440 157024 8449
rect 158076 8483 158128 8492
rect 158076 8449 158085 8483
rect 158085 8449 158119 8483
rect 158119 8449 158128 8483
rect 158076 8440 158128 8449
rect 155960 8347 156012 8356
rect 154304 8236 154356 8288
rect 155408 8236 155460 8288
rect 155960 8313 155969 8347
rect 155969 8313 156003 8347
rect 156003 8313 156012 8347
rect 155960 8304 156012 8313
rect 156144 8304 156196 8356
rect 157340 8304 157392 8356
rect 157524 8304 157576 8356
rect 158076 8304 158128 8356
rect 158260 8347 158312 8356
rect 158260 8313 158269 8347
rect 158269 8313 158303 8347
rect 158303 8313 158312 8347
rect 158260 8304 158312 8313
rect 20672 8134 20724 8186
rect 20736 8134 20788 8186
rect 20800 8134 20852 8186
rect 20864 8134 20916 8186
rect 20928 8134 20980 8186
rect 60117 8134 60169 8186
rect 60181 8134 60233 8186
rect 60245 8134 60297 8186
rect 60309 8134 60361 8186
rect 60373 8134 60425 8186
rect 99562 8134 99614 8186
rect 99626 8134 99678 8186
rect 99690 8134 99742 8186
rect 99754 8134 99806 8186
rect 99818 8134 99870 8186
rect 139007 8134 139059 8186
rect 139071 8134 139123 8186
rect 139135 8134 139187 8186
rect 139199 8134 139251 8186
rect 139263 8134 139315 8186
rect 10692 8032 10744 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 13728 8032 13780 8084
rect 14280 8032 14332 8084
rect 17868 8032 17920 8084
rect 18604 8075 18656 8084
rect 18604 8041 18613 8075
rect 18613 8041 18647 8075
rect 18647 8041 18656 8075
rect 18604 8032 18656 8041
rect 22192 8032 22244 8084
rect 23388 8032 23440 8084
rect 27252 8032 27304 8084
rect 31024 8075 31076 8084
rect 31024 8041 31033 8075
rect 31033 8041 31067 8075
rect 31067 8041 31076 8075
rect 31024 8032 31076 8041
rect 31576 8075 31628 8084
rect 31576 8041 31585 8075
rect 31585 8041 31619 8075
rect 31619 8041 31628 8075
rect 31576 8032 31628 8041
rect 5448 7896 5500 7948
rect 15844 7896 15896 7948
rect 5632 7828 5684 7880
rect 6000 7828 6052 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14832 7828 14884 7880
rect 15016 7828 15068 7880
rect 16120 7871 16172 7880
rect 6644 7760 6696 7812
rect 8392 7760 8444 7812
rect 4804 7735 4856 7744
rect 4804 7701 4813 7735
rect 4813 7701 4847 7735
rect 4847 7701 4856 7735
rect 4804 7692 4856 7701
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13728 7760 13780 7812
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 15476 7760 15528 7812
rect 24216 7964 24268 8016
rect 32496 8007 32548 8016
rect 32496 7973 32505 8007
rect 32505 7973 32539 8007
rect 32539 7973 32548 8007
rect 32496 7964 32548 7973
rect 33232 7964 33284 8016
rect 18972 7896 19024 7948
rect 35900 8032 35952 8084
rect 36636 8032 36688 8084
rect 37280 8032 37332 8084
rect 38568 8032 38620 8084
rect 38936 7964 38988 8016
rect 39120 8007 39172 8016
rect 39120 7973 39129 8007
rect 39129 7973 39163 8007
rect 39163 7973 39172 8007
rect 39120 7964 39172 7973
rect 37556 7896 37608 7948
rect 37832 7896 37884 7948
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 14004 7692 14056 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 20076 7828 20128 7880
rect 21272 7828 21324 7880
rect 25872 7871 25924 7880
rect 25872 7837 25881 7871
rect 25881 7837 25915 7871
rect 25915 7837 25924 7871
rect 25872 7828 25924 7837
rect 33600 7828 33652 7880
rect 33784 7828 33836 7880
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 36912 7871 36964 7880
rect 36912 7837 36921 7871
rect 36921 7837 36955 7871
rect 36955 7837 36964 7871
rect 36912 7828 36964 7837
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 41696 8032 41748 8084
rect 42800 8075 42852 8084
rect 42800 8041 42809 8075
rect 42809 8041 42843 8075
rect 42843 8041 42852 8075
rect 42800 8032 42852 8041
rect 42984 8032 43036 8084
rect 45376 8075 45428 8084
rect 45376 8041 45385 8075
rect 45385 8041 45419 8075
rect 45419 8041 45428 8075
rect 45376 8032 45428 8041
rect 45468 8032 45520 8084
rect 46204 8032 46256 8084
rect 48136 8032 48188 8084
rect 49148 8032 49200 8084
rect 49516 8032 49568 8084
rect 49700 8032 49752 8084
rect 40776 7828 40828 7880
rect 42616 7828 42668 7880
rect 45468 7896 45520 7948
rect 44640 7871 44692 7880
rect 44640 7837 44649 7871
rect 44649 7837 44683 7871
rect 44683 7837 44692 7871
rect 45836 7871 45888 7880
rect 44640 7828 44692 7837
rect 45836 7837 45845 7871
rect 45845 7837 45879 7871
rect 45879 7837 45888 7871
rect 45836 7828 45888 7837
rect 46020 7873 46072 7880
rect 46020 7839 46029 7873
rect 46029 7839 46063 7873
rect 46063 7839 46072 7873
rect 49332 7964 49384 8016
rect 56140 8032 56192 8084
rect 56784 8032 56836 8084
rect 59544 8075 59596 8084
rect 59544 8041 59553 8075
rect 59553 8041 59587 8075
rect 59587 8041 59596 8075
rect 59544 8032 59596 8041
rect 47032 7896 47084 7948
rect 50344 7896 50396 7948
rect 51356 7896 51408 7948
rect 52552 7896 52604 7948
rect 58808 7964 58860 8016
rect 61200 8007 61252 8016
rect 61200 7973 61209 8007
rect 61209 7973 61243 8007
rect 61243 7973 61252 8007
rect 61200 7964 61252 7973
rect 46020 7828 46072 7839
rect 21088 7760 21140 7812
rect 27896 7760 27948 7812
rect 32864 7760 32916 7812
rect 34060 7803 34112 7812
rect 34060 7769 34078 7803
rect 34078 7769 34112 7803
rect 34060 7760 34112 7769
rect 36636 7760 36688 7812
rect 39120 7760 39172 7812
rect 18972 7692 19024 7744
rect 23020 7692 23072 7744
rect 30564 7692 30616 7744
rect 32496 7692 32548 7744
rect 32956 7735 33008 7744
rect 32956 7701 32965 7735
rect 32965 7701 32999 7735
rect 32999 7701 33008 7735
rect 32956 7692 33008 7701
rect 33968 7692 34020 7744
rect 42892 7760 42944 7812
rect 51816 7828 51868 7880
rect 52460 7828 52512 7880
rect 54116 7871 54168 7880
rect 54116 7837 54125 7871
rect 54125 7837 54159 7871
rect 54159 7837 54168 7871
rect 54116 7828 54168 7837
rect 54208 7871 54260 7880
rect 54208 7837 54217 7871
rect 54217 7837 54251 7871
rect 54251 7837 54260 7871
rect 54944 7871 54996 7880
rect 54208 7828 54260 7837
rect 54944 7837 54953 7871
rect 54953 7837 54987 7871
rect 54987 7837 54996 7871
rect 54944 7828 54996 7837
rect 59544 7896 59596 7948
rect 61568 7896 61620 7948
rect 66720 8032 66772 8084
rect 68928 8075 68980 8084
rect 68928 8041 68937 8075
rect 68937 8041 68971 8075
rect 68971 8041 68980 8075
rect 68928 8032 68980 8041
rect 75276 8032 75328 8084
rect 76564 8032 76616 8084
rect 80612 8075 80664 8084
rect 80612 8041 80621 8075
rect 80621 8041 80655 8075
rect 80655 8041 80664 8075
rect 80612 8032 80664 8041
rect 83924 8032 83976 8084
rect 64972 7964 65024 8016
rect 65892 8007 65944 8016
rect 65892 7973 65901 8007
rect 65901 7973 65935 8007
rect 65935 7973 65944 8007
rect 65892 7964 65944 7973
rect 73620 7964 73672 8016
rect 112076 8032 112128 8084
rect 112168 8032 112220 8084
rect 49516 7760 49568 7812
rect 46664 7692 46716 7744
rect 47952 7692 48004 7744
rect 49792 7735 49844 7744
rect 49792 7701 49801 7735
rect 49801 7701 49835 7735
rect 49835 7701 49844 7735
rect 49792 7692 49844 7701
rect 50620 7760 50672 7812
rect 52276 7760 52328 7812
rect 59084 7828 59136 7880
rect 62672 7828 62724 7880
rect 65248 7828 65300 7880
rect 59268 7760 59320 7812
rect 60924 7760 60976 7812
rect 51908 7692 51960 7744
rect 53748 7692 53800 7744
rect 54760 7735 54812 7744
rect 54760 7701 54769 7735
rect 54769 7701 54803 7735
rect 54803 7701 54812 7735
rect 54760 7692 54812 7701
rect 60832 7692 60884 7744
rect 66904 7828 66956 7880
rect 80428 7896 80480 7948
rect 73252 7828 73304 7880
rect 74356 7828 74408 7880
rect 74632 7871 74684 7880
rect 74632 7837 74641 7871
rect 74641 7837 74675 7871
rect 74675 7837 74684 7871
rect 74632 7828 74684 7837
rect 75552 7828 75604 7880
rect 76288 7871 76340 7880
rect 76288 7837 76297 7871
rect 76297 7837 76331 7871
rect 76331 7837 76340 7871
rect 76288 7828 76340 7837
rect 80612 7828 80664 7880
rect 86408 7896 86460 7948
rect 87880 7896 87932 7948
rect 90088 7964 90140 8016
rect 90640 7964 90692 8016
rect 90732 7964 90784 8016
rect 92940 7964 92992 8016
rect 98276 7964 98328 8016
rect 100116 7964 100168 8016
rect 110420 7964 110472 8016
rect 112536 7964 112588 8016
rect 117136 7964 117188 8016
rect 119436 7964 119488 8016
rect 91376 7896 91428 7948
rect 93768 7896 93820 7948
rect 67088 7760 67140 7812
rect 81440 7760 81492 7812
rect 85580 7803 85632 7812
rect 75552 7692 75604 7744
rect 76012 7692 76064 7744
rect 81256 7692 81308 7744
rect 85580 7769 85598 7803
rect 85598 7769 85632 7803
rect 85580 7760 85632 7769
rect 87696 7871 87748 7880
rect 87696 7837 87705 7871
rect 87705 7837 87739 7871
rect 87739 7837 87748 7871
rect 87696 7828 87748 7837
rect 89628 7828 89680 7880
rect 90824 7828 90876 7880
rect 91008 7871 91060 7880
rect 91008 7837 91017 7871
rect 91017 7837 91051 7871
rect 91051 7837 91060 7871
rect 91008 7828 91060 7837
rect 92388 7828 92440 7880
rect 93032 7828 93084 7880
rect 95332 7871 95384 7880
rect 95332 7837 95341 7871
rect 95341 7837 95375 7871
rect 95375 7837 95384 7871
rect 95332 7828 95384 7837
rect 98092 7828 98144 7880
rect 105360 7828 105412 7880
rect 109132 7871 109184 7880
rect 109132 7837 109141 7871
rect 109141 7837 109175 7871
rect 109175 7837 109184 7871
rect 109132 7828 109184 7837
rect 117596 7896 117648 7948
rect 118608 7939 118660 7948
rect 118608 7905 118617 7939
rect 118617 7905 118651 7939
rect 118651 7905 118660 7939
rect 118608 7896 118660 7905
rect 121276 8032 121328 8084
rect 124036 8032 124088 8084
rect 124956 8032 125008 8084
rect 127164 8032 127216 8084
rect 121828 7964 121880 8016
rect 123024 7964 123076 8016
rect 123300 7964 123352 8016
rect 110972 7828 111024 7880
rect 111064 7828 111116 7880
rect 112720 7828 112772 7880
rect 112904 7871 112956 7880
rect 112904 7837 112913 7871
rect 112913 7837 112947 7871
rect 112947 7837 112956 7871
rect 112904 7828 112956 7837
rect 113088 7828 113140 7880
rect 117136 7828 117188 7880
rect 117412 7828 117464 7880
rect 118700 7828 118752 7880
rect 90732 7760 90784 7812
rect 92664 7803 92716 7812
rect 92664 7769 92682 7803
rect 92682 7769 92716 7803
rect 92664 7760 92716 7769
rect 98460 7760 98512 7812
rect 90824 7692 90876 7744
rect 91376 7692 91428 7744
rect 92480 7692 92532 7744
rect 92940 7692 92992 7744
rect 94044 7735 94096 7744
rect 94044 7701 94053 7735
rect 94053 7701 94087 7735
rect 94087 7701 94096 7735
rect 94044 7692 94096 7701
rect 95056 7692 95108 7744
rect 95148 7735 95200 7744
rect 95148 7701 95157 7735
rect 95157 7701 95191 7735
rect 95191 7701 95200 7735
rect 97816 7735 97868 7744
rect 95148 7692 95200 7701
rect 97816 7701 97825 7735
rect 97825 7701 97859 7735
rect 97859 7701 97868 7735
rect 97816 7692 97868 7701
rect 99196 7760 99248 7812
rect 104900 7760 104952 7812
rect 106740 7760 106792 7812
rect 107292 7760 107344 7812
rect 100300 7735 100352 7744
rect 100300 7701 100309 7735
rect 100309 7701 100343 7735
rect 100343 7701 100352 7735
rect 100300 7692 100352 7701
rect 107200 7692 107252 7744
rect 109776 7760 109828 7812
rect 109868 7760 109920 7812
rect 110696 7692 110748 7744
rect 112996 7760 113048 7812
rect 115480 7760 115532 7812
rect 116216 7803 116268 7812
rect 116216 7769 116225 7803
rect 116225 7769 116259 7803
rect 116259 7769 116268 7803
rect 116216 7760 116268 7769
rect 116308 7760 116360 7812
rect 114836 7692 114888 7744
rect 117044 7692 117096 7744
rect 121460 7760 121512 7812
rect 121644 7760 121696 7812
rect 122472 7760 122524 7812
rect 124220 7871 124272 7880
rect 124220 7837 124229 7871
rect 124229 7837 124263 7871
rect 124263 7837 124272 7871
rect 124220 7828 124272 7837
rect 124404 7896 124456 7948
rect 127072 7896 127124 7948
rect 130292 8032 130344 8084
rect 129648 7964 129700 8016
rect 130384 7964 130436 8016
rect 134340 7964 134392 8016
rect 124036 7760 124088 7812
rect 122840 7692 122892 7744
rect 123208 7735 123260 7744
rect 123208 7701 123217 7735
rect 123217 7701 123251 7735
rect 123251 7701 123260 7735
rect 123208 7692 123260 7701
rect 125876 7735 125928 7744
rect 125876 7701 125885 7735
rect 125885 7701 125919 7735
rect 125919 7701 125928 7735
rect 125876 7692 125928 7701
rect 126244 7692 126296 7744
rect 127072 7735 127124 7744
rect 127072 7701 127081 7735
rect 127081 7701 127115 7735
rect 127115 7701 127124 7735
rect 127072 7692 127124 7701
rect 129280 7760 129332 7812
rect 129924 7871 129976 7880
rect 129924 7837 129933 7871
rect 129933 7837 129967 7871
rect 129967 7837 129976 7871
rect 130108 7871 130160 7880
rect 129924 7828 129976 7837
rect 130108 7837 130117 7871
rect 130117 7837 130151 7871
rect 130151 7837 130160 7871
rect 130108 7828 130160 7837
rect 130660 7871 130712 7880
rect 130660 7837 130669 7871
rect 130669 7837 130703 7871
rect 130703 7837 130712 7871
rect 130660 7828 130712 7837
rect 132868 7896 132920 7948
rect 132960 7896 133012 7948
rect 133144 7896 133196 7948
rect 133604 7896 133656 7948
rect 134800 7896 134852 7948
rect 136456 8032 136508 8084
rect 137836 8032 137888 8084
rect 138204 8032 138256 8084
rect 138572 8032 138624 8084
rect 138664 7896 138716 7948
rect 142988 8032 143040 8084
rect 140228 7964 140280 8016
rect 141424 8007 141476 8016
rect 130568 7760 130620 7812
rect 133512 7828 133564 7880
rect 133788 7828 133840 7880
rect 135720 7828 135772 7880
rect 141056 7896 141108 7948
rect 140688 7828 140740 7880
rect 141424 7973 141433 8007
rect 141433 7973 141467 8007
rect 141467 7973 141476 8007
rect 141424 7964 141476 7973
rect 141332 7896 141384 7948
rect 144736 8032 144788 8084
rect 142988 7828 143040 7880
rect 143080 7871 143132 7880
rect 143080 7837 143089 7871
rect 143089 7837 143123 7871
rect 143123 7837 143132 7871
rect 143080 7828 143132 7837
rect 135352 7760 135404 7812
rect 136364 7803 136416 7812
rect 136364 7769 136373 7803
rect 136373 7769 136407 7803
rect 136407 7769 136416 7803
rect 136364 7760 136416 7769
rect 137744 7760 137796 7812
rect 132960 7692 133012 7744
rect 133696 7692 133748 7744
rect 134432 7735 134484 7744
rect 134432 7701 134441 7735
rect 134441 7701 134475 7735
rect 134475 7701 134484 7735
rect 134432 7692 134484 7701
rect 137376 7692 137428 7744
rect 139860 7803 139912 7812
rect 139860 7769 139878 7803
rect 139878 7769 139912 7803
rect 139860 7760 139912 7769
rect 140412 7760 140464 7812
rect 139768 7692 139820 7744
rect 141056 7760 141108 7812
rect 144368 7828 144420 7880
rect 145196 7964 145248 8016
rect 147220 7964 147272 8016
rect 148140 7964 148192 8016
rect 146760 7896 146812 7948
rect 147036 7896 147088 7948
rect 149888 8032 149940 8084
rect 150164 8032 150216 8084
rect 151820 8032 151872 8084
rect 152280 8032 152332 8084
rect 152372 8032 152424 8084
rect 154764 8032 154816 8084
rect 155868 8032 155920 8084
rect 149244 7964 149296 8016
rect 154304 7964 154356 8016
rect 150900 7896 150952 7948
rect 145748 7760 145800 7812
rect 146392 7828 146444 7880
rect 147312 7871 147364 7880
rect 147312 7837 147321 7871
rect 147321 7837 147355 7871
rect 147355 7837 147364 7871
rect 147312 7828 147364 7837
rect 142252 7692 142304 7744
rect 142436 7735 142488 7744
rect 142436 7701 142445 7735
rect 142445 7701 142479 7735
rect 142479 7701 142488 7735
rect 142436 7692 142488 7701
rect 142988 7692 143040 7744
rect 144644 7692 144696 7744
rect 146300 7692 146352 7744
rect 147128 7760 147180 7812
rect 147956 7828 148008 7880
rect 148232 7871 148284 7880
rect 148232 7837 148241 7871
rect 148241 7837 148275 7871
rect 148275 7837 148284 7871
rect 148232 7828 148284 7837
rect 148968 7828 149020 7880
rect 148324 7760 148376 7812
rect 148876 7760 148928 7812
rect 148140 7692 148192 7744
rect 149336 7760 149388 7812
rect 150164 7803 150216 7812
rect 150164 7769 150173 7803
rect 150173 7769 150207 7803
rect 150207 7769 150216 7803
rect 150164 7760 150216 7769
rect 150532 7828 150584 7880
rect 151176 7828 151228 7880
rect 152280 7871 152332 7880
rect 152280 7837 152289 7871
rect 152289 7837 152323 7871
rect 152323 7837 152332 7871
rect 152280 7828 152332 7837
rect 152372 7871 152424 7880
rect 152372 7837 152381 7871
rect 152381 7837 152415 7871
rect 152415 7837 152424 7871
rect 152924 7896 152976 7948
rect 152372 7828 152424 7837
rect 153752 7871 153804 7880
rect 153752 7837 153761 7871
rect 153761 7837 153795 7871
rect 153795 7837 153804 7871
rect 153752 7828 153804 7837
rect 154028 7828 154080 7880
rect 155776 7896 155828 7948
rect 156052 7828 156104 7880
rect 156604 7871 156656 7880
rect 156604 7837 156613 7871
rect 156613 7837 156647 7871
rect 156647 7837 156656 7871
rect 156604 7828 156656 7837
rect 155500 7760 155552 7812
rect 151544 7692 151596 7744
rect 151820 7692 151872 7744
rect 152188 7692 152240 7744
rect 153384 7735 153436 7744
rect 153384 7701 153393 7735
rect 153393 7701 153427 7735
rect 153427 7701 153436 7735
rect 153384 7692 153436 7701
rect 154028 7692 154080 7744
rect 155868 7735 155920 7744
rect 155868 7701 155877 7735
rect 155877 7701 155911 7735
rect 155911 7701 155920 7735
rect 155868 7692 155920 7701
rect 156144 7692 156196 7744
rect 157524 7692 157576 7744
rect 158260 7692 158312 7744
rect 40394 7590 40446 7642
rect 40458 7590 40510 7642
rect 40522 7590 40574 7642
rect 40586 7590 40638 7642
rect 40650 7590 40702 7642
rect 79839 7590 79891 7642
rect 79903 7590 79955 7642
rect 79967 7590 80019 7642
rect 80031 7590 80083 7642
rect 80095 7590 80147 7642
rect 119284 7590 119336 7642
rect 119348 7590 119400 7642
rect 119412 7590 119464 7642
rect 119476 7590 119528 7642
rect 119540 7590 119592 7642
rect 158729 7590 158781 7642
rect 158793 7590 158845 7642
rect 158857 7590 158909 7642
rect 158921 7590 158973 7642
rect 158985 7590 159037 7642
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 6000 7531 6052 7540
rect 6000 7497 6009 7531
rect 6009 7497 6043 7531
rect 6043 7497 6052 7531
rect 6000 7488 6052 7497
rect 6736 7488 6788 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 23296 7488 23348 7540
rect 32864 7531 32916 7540
rect 16396 7420 16448 7472
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5080 7352 5132 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 16856 7352 16908 7404
rect 17868 7352 17920 7404
rect 11152 7284 11204 7336
rect 17776 7284 17828 7336
rect 18604 7420 18656 7472
rect 12716 7216 12768 7268
rect 15844 7216 15896 7268
rect 21640 7352 21692 7404
rect 21824 7352 21876 7404
rect 26608 7352 26660 7404
rect 30564 7420 30616 7472
rect 31024 7420 31076 7472
rect 32864 7497 32873 7531
rect 32873 7497 32907 7531
rect 32907 7497 32916 7531
rect 32864 7488 32916 7497
rect 38568 7531 38620 7540
rect 33784 7420 33836 7472
rect 38568 7497 38577 7531
rect 38577 7497 38611 7531
rect 38611 7497 38620 7531
rect 38568 7488 38620 7497
rect 40316 7488 40368 7540
rect 42064 7488 42116 7540
rect 43168 7488 43220 7540
rect 45376 7488 45428 7540
rect 49608 7488 49660 7540
rect 49792 7488 49844 7540
rect 57704 7488 57756 7540
rect 57796 7488 57848 7540
rect 58532 7488 58584 7540
rect 59176 7488 59228 7540
rect 59728 7531 59780 7540
rect 59728 7497 59737 7531
rect 59737 7497 59771 7531
rect 59771 7497 59780 7531
rect 59728 7488 59780 7497
rect 63224 7531 63276 7540
rect 63224 7497 63233 7531
rect 63233 7497 63267 7531
rect 63267 7497 63276 7531
rect 63224 7488 63276 7497
rect 64788 7531 64840 7540
rect 64788 7497 64797 7531
rect 64797 7497 64831 7531
rect 64831 7497 64840 7531
rect 64788 7488 64840 7497
rect 65248 7531 65300 7540
rect 65248 7497 65257 7531
rect 65257 7497 65291 7531
rect 65291 7497 65300 7531
rect 65248 7488 65300 7497
rect 67088 7531 67140 7540
rect 67088 7497 67097 7531
rect 67097 7497 67131 7531
rect 67131 7497 67140 7531
rect 67088 7488 67140 7497
rect 45560 7420 45612 7472
rect 45836 7420 45888 7472
rect 49516 7420 49568 7472
rect 54760 7420 54812 7472
rect 64236 7420 64288 7472
rect 23940 7284 23992 7336
rect 26332 7327 26384 7336
rect 26332 7293 26341 7327
rect 26341 7293 26375 7327
rect 26375 7293 26384 7327
rect 26332 7284 26384 7293
rect 18880 7216 18932 7268
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 18328 7148 18380 7200
rect 19156 7216 19208 7268
rect 33968 7395 34020 7404
rect 33968 7361 33986 7395
rect 33986 7361 34020 7395
rect 34244 7395 34296 7404
rect 33968 7352 34020 7361
rect 34244 7361 34253 7395
rect 34253 7361 34287 7395
rect 34287 7361 34296 7395
rect 34244 7352 34296 7361
rect 34888 7352 34940 7404
rect 36452 7352 36504 7404
rect 37832 7352 37884 7404
rect 40776 7352 40828 7404
rect 41236 7395 41288 7404
rect 33140 7284 33192 7336
rect 37188 7284 37240 7336
rect 38476 7284 38528 7336
rect 41236 7361 41245 7395
rect 41245 7361 41279 7395
rect 41279 7361 41288 7395
rect 41236 7352 41288 7361
rect 42432 7352 42484 7404
rect 49700 7352 49752 7404
rect 53104 7352 53156 7404
rect 53840 7395 53892 7404
rect 53840 7361 53849 7395
rect 53849 7361 53883 7395
rect 53883 7361 53892 7395
rect 53840 7352 53892 7361
rect 54300 7352 54352 7404
rect 60004 7352 60056 7404
rect 60556 7395 60608 7404
rect 60556 7361 60565 7395
rect 60565 7361 60599 7395
rect 60599 7361 60608 7395
rect 60556 7352 60608 7361
rect 61568 7352 61620 7404
rect 63408 7395 63460 7404
rect 45836 7284 45888 7336
rect 52368 7327 52420 7336
rect 52368 7293 52377 7327
rect 52377 7293 52411 7327
rect 52411 7293 52420 7327
rect 52368 7284 52420 7293
rect 62672 7284 62724 7336
rect 63408 7361 63417 7395
rect 63417 7361 63451 7395
rect 63451 7361 63460 7395
rect 63408 7352 63460 7361
rect 64604 7395 64656 7404
rect 64604 7361 64613 7395
rect 64613 7361 64647 7395
rect 64647 7361 64656 7395
rect 64604 7352 64656 7361
rect 66996 7352 67048 7404
rect 73620 7488 73672 7540
rect 74724 7488 74776 7540
rect 72884 7352 72936 7404
rect 83464 7420 83516 7472
rect 85304 7488 85356 7540
rect 86224 7488 86276 7540
rect 93492 7488 93544 7540
rect 96896 7488 96948 7540
rect 97356 7531 97408 7540
rect 97356 7497 97365 7531
rect 97365 7497 97399 7531
rect 97399 7497 97408 7531
rect 97356 7488 97408 7497
rect 97448 7488 97500 7540
rect 108856 7488 108908 7540
rect 89352 7420 89404 7472
rect 89812 7420 89864 7472
rect 116768 7488 116820 7540
rect 83096 7352 83148 7404
rect 84660 7395 84712 7404
rect 84660 7361 84669 7395
rect 84669 7361 84703 7395
rect 84703 7361 84712 7395
rect 84660 7352 84712 7361
rect 73160 7284 73212 7336
rect 75920 7327 75972 7336
rect 75920 7293 75929 7327
rect 75929 7293 75963 7327
rect 75963 7293 75972 7327
rect 75920 7284 75972 7293
rect 79048 7327 79100 7336
rect 79048 7293 79057 7327
rect 79057 7293 79091 7327
rect 79091 7293 79100 7327
rect 79048 7284 79100 7293
rect 81072 7284 81124 7336
rect 90824 7352 90876 7404
rect 90916 7352 90968 7404
rect 93492 7352 93544 7404
rect 96528 7395 96580 7404
rect 96528 7361 96546 7395
rect 96546 7361 96580 7395
rect 96804 7395 96856 7404
rect 96528 7352 96580 7361
rect 96804 7361 96813 7395
rect 96813 7361 96847 7395
rect 96847 7361 96856 7395
rect 96804 7352 96856 7361
rect 97356 7352 97408 7404
rect 110604 7420 110656 7472
rect 111616 7463 111668 7472
rect 111616 7429 111650 7463
rect 111650 7429 111668 7463
rect 111616 7420 111668 7429
rect 110696 7395 110748 7404
rect 110696 7361 110705 7395
rect 110705 7361 110739 7395
rect 110739 7361 110748 7395
rect 110696 7352 110748 7361
rect 114100 7395 114152 7404
rect 114100 7361 114109 7395
rect 114109 7361 114143 7395
rect 114143 7361 114152 7395
rect 114100 7352 114152 7361
rect 116952 7352 117004 7404
rect 19248 7148 19300 7200
rect 22560 7148 22612 7200
rect 35348 7148 35400 7200
rect 42892 7216 42944 7268
rect 50804 7216 50856 7268
rect 60832 7216 60884 7268
rect 86224 7284 86276 7336
rect 44364 7148 44416 7200
rect 45744 7148 45796 7200
rect 47032 7148 47084 7200
rect 61108 7148 61160 7200
rect 68376 7191 68428 7200
rect 68376 7157 68385 7191
rect 68385 7157 68419 7191
rect 68419 7157 68428 7191
rect 68376 7148 68428 7157
rect 80428 7191 80480 7200
rect 80428 7157 80437 7191
rect 80437 7157 80471 7191
rect 80471 7157 80480 7191
rect 80428 7148 80480 7157
rect 82636 7216 82688 7268
rect 82452 7148 82504 7200
rect 83096 7191 83148 7200
rect 83096 7157 83105 7191
rect 83105 7157 83139 7191
rect 83139 7157 83148 7191
rect 83096 7148 83148 7157
rect 83648 7148 83700 7200
rect 85580 7148 85632 7200
rect 86408 7148 86460 7200
rect 86776 7148 86828 7200
rect 87696 7148 87748 7200
rect 91376 7148 91428 7200
rect 92940 7191 92992 7200
rect 92940 7157 92949 7191
rect 92949 7157 92983 7191
rect 92983 7157 92992 7191
rect 93492 7191 93544 7200
rect 92940 7148 92992 7157
rect 93492 7157 93501 7191
rect 93501 7157 93535 7191
rect 93535 7157 93544 7191
rect 93492 7148 93544 7157
rect 93584 7148 93636 7200
rect 96896 7284 96948 7336
rect 99196 7284 99248 7336
rect 107016 7284 107068 7336
rect 96988 7216 97040 7268
rect 110328 7216 110380 7268
rect 97448 7148 97500 7200
rect 97540 7148 97592 7200
rect 109868 7148 109920 7200
rect 110052 7191 110104 7200
rect 110052 7157 110061 7191
rect 110061 7157 110095 7191
rect 110095 7157 110104 7191
rect 110052 7148 110104 7157
rect 110972 7284 111024 7336
rect 111340 7327 111392 7336
rect 111340 7293 111349 7327
rect 111349 7293 111383 7327
rect 111383 7293 111392 7327
rect 111340 7284 111392 7293
rect 112444 7284 112496 7336
rect 112904 7284 112956 7336
rect 113272 7284 113324 7336
rect 118424 7420 118476 7472
rect 123116 7420 123168 7472
rect 124404 7420 124456 7472
rect 125416 7420 125468 7472
rect 126336 7420 126388 7472
rect 119068 7395 119120 7404
rect 119068 7361 119097 7395
rect 119097 7361 119120 7395
rect 119068 7352 119120 7361
rect 112720 7191 112772 7200
rect 112720 7157 112729 7191
rect 112729 7157 112763 7191
rect 112763 7157 112772 7191
rect 112720 7148 112772 7157
rect 112904 7148 112956 7200
rect 114928 7148 114980 7200
rect 117412 7191 117464 7200
rect 117412 7157 117421 7191
rect 117421 7157 117455 7191
rect 117455 7157 117464 7191
rect 117412 7148 117464 7157
rect 118976 7148 119028 7200
rect 119988 7191 120040 7200
rect 119988 7157 119997 7191
rect 119997 7157 120031 7191
rect 120031 7157 120040 7191
rect 119988 7148 120040 7157
rect 124312 7352 124364 7404
rect 127808 7488 127860 7540
rect 127072 7420 127124 7472
rect 128912 7488 128964 7540
rect 129372 7531 129424 7540
rect 129372 7497 129381 7531
rect 129381 7497 129415 7531
rect 129415 7497 129424 7531
rect 129372 7488 129424 7497
rect 130200 7531 130252 7540
rect 130200 7497 130209 7531
rect 130209 7497 130243 7531
rect 130243 7497 130252 7531
rect 130200 7488 130252 7497
rect 130844 7531 130896 7540
rect 130844 7497 130853 7531
rect 130853 7497 130887 7531
rect 130887 7497 130896 7531
rect 130844 7488 130896 7497
rect 131212 7488 131264 7540
rect 132040 7488 132092 7540
rect 121644 7284 121696 7336
rect 121736 7216 121788 7268
rect 122012 7148 122064 7200
rect 123300 7284 123352 7336
rect 123668 7284 123720 7336
rect 125416 7284 125468 7336
rect 126428 7284 126480 7336
rect 126612 7327 126664 7336
rect 126612 7293 126621 7327
rect 126621 7293 126655 7327
rect 126655 7293 126664 7327
rect 126612 7284 126664 7293
rect 127256 7284 127308 7336
rect 127808 7284 127860 7336
rect 128912 7352 128964 7404
rect 129280 7420 129332 7472
rect 131948 7420 132000 7472
rect 137560 7488 137612 7540
rect 139216 7488 139268 7540
rect 141792 7488 141844 7540
rect 141976 7488 142028 7540
rect 142436 7488 142488 7540
rect 146208 7488 146260 7540
rect 129832 7352 129884 7404
rect 130844 7352 130896 7404
rect 134800 7395 134852 7404
rect 129556 7284 129608 7336
rect 134800 7361 134809 7395
rect 134809 7361 134843 7395
rect 134843 7361 134852 7395
rect 134800 7352 134852 7361
rect 135352 7395 135404 7404
rect 135352 7361 135361 7395
rect 135361 7361 135395 7395
rect 135395 7361 135404 7395
rect 135352 7352 135404 7361
rect 137284 7420 137336 7472
rect 138020 7352 138072 7404
rect 131304 7284 131356 7336
rect 132500 7284 132552 7336
rect 122472 7148 122524 7200
rect 133788 7216 133840 7268
rect 139216 7395 139268 7404
rect 139216 7361 139225 7395
rect 139225 7361 139259 7395
rect 139259 7361 139268 7395
rect 140872 7395 140924 7404
rect 139216 7352 139268 7361
rect 140872 7361 140881 7395
rect 140881 7361 140915 7395
rect 140915 7361 140924 7395
rect 140872 7352 140924 7361
rect 144000 7463 144052 7472
rect 144000 7429 144034 7463
rect 144034 7429 144052 7463
rect 144000 7420 144052 7429
rect 145288 7420 145340 7472
rect 144368 7352 144420 7404
rect 146944 7420 146996 7472
rect 148140 7420 148192 7472
rect 148324 7488 148376 7540
rect 150440 7488 150492 7540
rect 150808 7531 150860 7540
rect 150808 7497 150817 7531
rect 150817 7497 150851 7531
rect 150851 7497 150860 7531
rect 150808 7488 150860 7497
rect 151084 7488 151136 7540
rect 154580 7488 154632 7540
rect 155592 7488 155644 7540
rect 155868 7488 155920 7540
rect 156328 7488 156380 7540
rect 157616 7531 157668 7540
rect 157616 7497 157625 7531
rect 157625 7497 157659 7531
rect 157659 7497 157668 7531
rect 157616 7488 157668 7497
rect 146392 7352 146444 7404
rect 148600 7420 148652 7472
rect 149336 7420 149388 7472
rect 149520 7420 149572 7472
rect 148968 7352 149020 7404
rect 155684 7420 155736 7472
rect 155776 7420 155828 7472
rect 143264 7327 143316 7336
rect 124220 7148 124272 7200
rect 126152 7191 126204 7200
rect 126152 7157 126161 7191
rect 126161 7157 126195 7191
rect 126195 7157 126204 7191
rect 126152 7148 126204 7157
rect 126336 7148 126388 7200
rect 132040 7148 132092 7200
rect 132500 7148 132552 7200
rect 136824 7216 136876 7268
rect 135628 7148 135680 7200
rect 136640 7191 136692 7200
rect 136640 7157 136649 7191
rect 136649 7157 136683 7191
rect 136683 7157 136692 7191
rect 136640 7148 136692 7157
rect 138480 7148 138532 7200
rect 138940 7148 138992 7200
rect 140504 7216 140556 7268
rect 139492 7148 139544 7200
rect 140044 7148 140096 7200
rect 140136 7148 140188 7200
rect 143264 7293 143273 7327
rect 143273 7293 143307 7327
rect 143307 7293 143316 7327
rect 143264 7284 143316 7293
rect 143448 7284 143500 7336
rect 145012 7284 145064 7336
rect 146576 7284 146628 7336
rect 149244 7284 149296 7336
rect 153660 7352 153712 7404
rect 154304 7395 154356 7404
rect 154304 7361 154313 7395
rect 154313 7361 154347 7395
rect 154347 7361 154356 7395
rect 154304 7352 154356 7361
rect 152188 7327 152240 7336
rect 152188 7293 152197 7327
rect 152197 7293 152231 7327
rect 152231 7293 152240 7327
rect 152188 7284 152240 7293
rect 153292 7284 153344 7336
rect 153568 7284 153620 7336
rect 153936 7284 153988 7336
rect 145380 7216 145432 7268
rect 145932 7216 145984 7268
rect 146024 7148 146076 7200
rect 146116 7148 146168 7200
rect 147864 7216 147916 7268
rect 148140 7148 148192 7200
rect 149796 7148 149848 7200
rect 153476 7216 153528 7268
rect 154764 7284 154816 7336
rect 155592 7352 155644 7404
rect 156052 7352 156104 7404
rect 156972 7395 157024 7404
rect 156972 7361 156981 7395
rect 156981 7361 157015 7395
rect 157015 7361 157024 7395
rect 156972 7352 157024 7361
rect 157800 7395 157852 7404
rect 157800 7361 157809 7395
rect 157809 7361 157843 7395
rect 157843 7361 157852 7395
rect 157800 7352 157852 7361
rect 156236 7284 156288 7336
rect 156696 7284 156748 7336
rect 155684 7216 155736 7268
rect 157524 7216 157576 7268
rect 154396 7148 154448 7200
rect 154764 7148 154816 7200
rect 155776 7148 155828 7200
rect 156972 7148 157024 7200
rect 20672 7046 20724 7098
rect 20736 7046 20788 7098
rect 20800 7046 20852 7098
rect 20864 7046 20916 7098
rect 20928 7046 20980 7098
rect 60117 7046 60169 7098
rect 60181 7046 60233 7098
rect 60245 7046 60297 7098
rect 60309 7046 60361 7098
rect 60373 7046 60425 7098
rect 99562 7046 99614 7098
rect 99626 7046 99678 7098
rect 99690 7046 99742 7098
rect 99754 7046 99806 7098
rect 99818 7046 99870 7098
rect 139007 7046 139059 7098
rect 139071 7046 139123 7098
rect 139135 7046 139187 7098
rect 139199 7046 139251 7098
rect 139263 7046 139315 7098
rect 13452 6944 13504 6996
rect 14832 6944 14884 6996
rect 17868 6876 17920 6928
rect 15108 6808 15160 6860
rect 20260 6944 20312 6996
rect 30380 6944 30432 6996
rect 34888 6987 34940 6996
rect 34888 6953 34897 6987
rect 34897 6953 34931 6987
rect 34931 6953 34940 6987
rect 34888 6944 34940 6953
rect 37648 6987 37700 6996
rect 37648 6953 37657 6987
rect 37657 6953 37691 6987
rect 37691 6953 37700 6987
rect 37648 6944 37700 6953
rect 40224 6944 40276 6996
rect 19892 6808 19944 6860
rect 20076 6851 20128 6860
rect 20076 6817 20085 6851
rect 20085 6817 20119 6851
rect 20119 6817 20128 6851
rect 20076 6808 20128 6817
rect 21732 6808 21784 6860
rect 26332 6808 26384 6860
rect 30196 6808 30248 6860
rect 32036 6808 32088 6860
rect 33968 6876 34020 6928
rect 37188 6876 37240 6928
rect 33232 6808 33284 6860
rect 33508 6851 33560 6860
rect 33508 6817 33517 6851
rect 33517 6817 33551 6851
rect 33551 6817 33560 6851
rect 33508 6808 33560 6817
rect 37832 6808 37884 6860
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 13268 6740 13320 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15292 6740 15344 6792
rect 16488 6783 16540 6792
rect 16488 6749 16522 6783
rect 16522 6749 16540 6783
rect 16488 6740 16540 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 13728 6715 13780 6724
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 4068 6604 4120 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16856 6604 16908 6656
rect 17224 6604 17276 6656
rect 19892 6672 19944 6724
rect 21180 6740 21232 6792
rect 27068 6783 27120 6792
rect 18880 6604 18932 6656
rect 21456 6647 21508 6656
rect 21456 6613 21465 6647
rect 21465 6613 21499 6647
rect 21499 6613 21508 6647
rect 21456 6604 21508 6613
rect 23572 6672 23624 6724
rect 22560 6604 22612 6656
rect 23848 6604 23900 6656
rect 27068 6749 27077 6783
rect 27077 6749 27111 6783
rect 27111 6749 27120 6783
rect 27068 6740 27120 6749
rect 33968 6740 34020 6792
rect 36544 6783 36596 6792
rect 36544 6749 36553 6783
rect 36553 6749 36587 6783
rect 36587 6749 36596 6783
rect 36544 6740 36596 6749
rect 37004 6783 37056 6792
rect 37004 6749 37013 6783
rect 37013 6749 37047 6783
rect 37047 6749 37056 6783
rect 37004 6740 37056 6749
rect 45008 6808 45060 6860
rect 52368 6944 52420 6996
rect 54208 6944 54260 6996
rect 63684 6987 63736 6996
rect 63684 6953 63693 6987
rect 63693 6953 63727 6987
rect 63727 6953 63736 6987
rect 63684 6944 63736 6953
rect 50528 6876 50580 6928
rect 55772 6876 55824 6928
rect 61660 6876 61712 6928
rect 119988 6944 120040 6996
rect 83004 6876 83056 6928
rect 86776 6876 86828 6928
rect 108948 6876 109000 6928
rect 110604 6919 110656 6928
rect 43536 6783 43588 6792
rect 30564 6672 30616 6724
rect 30656 6672 30708 6724
rect 43536 6749 43545 6783
rect 43545 6749 43579 6783
rect 43579 6749 43588 6783
rect 43536 6740 43588 6749
rect 44180 6740 44232 6792
rect 45100 6740 45152 6792
rect 50436 6808 50488 6860
rect 52092 6851 52144 6860
rect 52092 6817 52101 6851
rect 52101 6817 52135 6851
rect 52135 6817 52144 6851
rect 52092 6808 52144 6817
rect 38384 6715 38436 6724
rect 38384 6681 38418 6715
rect 38418 6681 38436 6715
rect 38384 6672 38436 6681
rect 45468 6672 45520 6724
rect 46204 6740 46256 6792
rect 52276 6740 52328 6792
rect 56324 6808 56376 6860
rect 58992 6808 59044 6860
rect 54300 6740 54352 6792
rect 57520 6740 57572 6792
rect 69112 6808 69164 6860
rect 46572 6672 46624 6724
rect 47032 6672 47084 6724
rect 50712 6672 50764 6724
rect 52184 6672 52236 6724
rect 57152 6672 57204 6724
rect 59728 6740 59780 6792
rect 64420 6740 64472 6792
rect 64512 6740 64564 6792
rect 66536 6783 66588 6792
rect 60464 6672 60516 6724
rect 66536 6749 66545 6783
rect 66545 6749 66579 6783
rect 66579 6749 66588 6783
rect 66536 6740 66588 6749
rect 73160 6740 73212 6792
rect 73804 6740 73856 6792
rect 75920 6740 75972 6792
rect 79048 6740 79100 6792
rect 79140 6740 79192 6792
rect 81164 6808 81216 6860
rect 25596 6604 25648 6656
rect 26240 6604 26292 6656
rect 26884 6647 26936 6656
rect 26884 6613 26893 6647
rect 26893 6613 26927 6647
rect 26927 6613 26936 6647
rect 26884 6604 26936 6613
rect 36360 6647 36412 6656
rect 36360 6613 36369 6647
rect 36369 6613 36403 6647
rect 36403 6613 36412 6647
rect 36360 6604 36412 6613
rect 36452 6604 36504 6656
rect 43536 6604 43588 6656
rect 44364 6647 44416 6656
rect 44364 6613 44373 6647
rect 44373 6613 44407 6647
rect 44407 6613 44416 6647
rect 44364 6604 44416 6613
rect 53380 6604 53432 6656
rect 58624 6604 58676 6656
rect 66628 6672 66680 6724
rect 66260 6604 66312 6656
rect 67916 6647 67968 6656
rect 67916 6613 67925 6647
rect 67925 6613 67959 6647
rect 67959 6613 67968 6647
rect 67916 6604 67968 6613
rect 72332 6647 72384 6656
rect 72332 6613 72341 6647
rect 72341 6613 72375 6647
rect 72375 6613 72384 6647
rect 72332 6604 72384 6613
rect 73344 6672 73396 6724
rect 75184 6672 75236 6724
rect 76012 6672 76064 6724
rect 81164 6672 81216 6724
rect 82636 6783 82688 6792
rect 82636 6749 82645 6783
rect 82645 6749 82679 6783
rect 82679 6749 82688 6783
rect 82636 6740 82688 6749
rect 88340 6740 88392 6792
rect 74632 6604 74684 6656
rect 75092 6604 75144 6656
rect 79324 6604 79376 6656
rect 80612 6604 80664 6656
rect 86408 6647 86460 6656
rect 86408 6613 86417 6647
rect 86417 6613 86451 6647
rect 86451 6613 86460 6647
rect 86408 6604 86460 6613
rect 92204 6740 92256 6792
rect 93308 6851 93360 6860
rect 93308 6817 93317 6851
rect 93317 6817 93351 6851
rect 93351 6817 93360 6851
rect 93308 6808 93360 6817
rect 96804 6808 96856 6860
rect 96896 6808 96948 6860
rect 101588 6808 101640 6860
rect 103612 6808 103664 6860
rect 106924 6808 106976 6860
rect 108396 6851 108448 6860
rect 108396 6817 108405 6851
rect 108405 6817 108439 6851
rect 108439 6817 108448 6851
rect 108856 6851 108908 6860
rect 108396 6808 108448 6817
rect 108856 6817 108865 6851
rect 108865 6817 108899 6851
rect 108899 6817 108908 6851
rect 108856 6808 108908 6817
rect 110604 6885 110613 6919
rect 110613 6885 110647 6919
rect 110647 6885 110656 6919
rect 110604 6876 110656 6885
rect 111064 6919 111116 6928
rect 111064 6885 111073 6919
rect 111073 6885 111107 6919
rect 111107 6885 111116 6919
rect 111064 6876 111116 6885
rect 111340 6876 111392 6928
rect 111524 6876 111576 6928
rect 112904 6876 112956 6928
rect 114468 6876 114520 6928
rect 105452 6740 105504 6792
rect 105728 6740 105780 6792
rect 92480 6672 92532 6724
rect 93216 6672 93268 6724
rect 99380 6672 99432 6724
rect 101588 6672 101640 6724
rect 107384 6672 107436 6724
rect 110604 6740 110656 6792
rect 110696 6740 110748 6792
rect 113088 6808 113140 6860
rect 114560 6851 114612 6860
rect 114560 6817 114569 6851
rect 114569 6817 114603 6851
rect 114603 6817 114612 6851
rect 114560 6808 114612 6817
rect 116676 6876 116728 6928
rect 120632 6944 120684 6996
rect 124220 6944 124272 6996
rect 122012 6876 122064 6928
rect 123116 6876 123168 6928
rect 115480 6808 115532 6860
rect 116308 6808 116360 6860
rect 116860 6808 116912 6860
rect 118608 6808 118660 6860
rect 121644 6851 121696 6860
rect 121644 6817 121653 6851
rect 121653 6817 121687 6851
rect 121687 6817 121696 6851
rect 121644 6808 121696 6817
rect 122564 6808 122616 6860
rect 124956 6808 125008 6860
rect 125232 6808 125284 6860
rect 126428 6944 126480 6996
rect 126336 6876 126388 6928
rect 128544 6876 128596 6928
rect 129924 6944 129976 6996
rect 130844 6987 130896 6996
rect 130844 6953 130853 6987
rect 130853 6953 130887 6987
rect 130887 6953 130896 6987
rect 130844 6944 130896 6953
rect 130936 6944 130988 6996
rect 133604 6944 133656 6996
rect 133788 6944 133840 6996
rect 134340 6944 134392 6996
rect 137928 6944 137980 6996
rect 138572 6944 138624 6996
rect 139492 6944 139544 6996
rect 139860 6944 139912 6996
rect 132868 6876 132920 6928
rect 135536 6876 135588 6928
rect 141148 6876 141200 6928
rect 111432 6783 111484 6792
rect 111432 6749 111441 6783
rect 111441 6749 111475 6783
rect 111475 6749 111484 6783
rect 111432 6740 111484 6749
rect 114836 6740 114888 6792
rect 115020 6740 115072 6792
rect 118700 6740 118752 6792
rect 120816 6740 120868 6792
rect 122656 6783 122708 6792
rect 111616 6672 111668 6724
rect 115388 6672 115440 6724
rect 122656 6749 122665 6783
rect 122665 6749 122699 6783
rect 122699 6749 122708 6783
rect 122656 6740 122708 6749
rect 123024 6740 123076 6792
rect 124864 6783 124916 6792
rect 124864 6749 124873 6783
rect 124873 6749 124907 6783
rect 124907 6749 124916 6783
rect 124864 6740 124916 6749
rect 125416 6740 125468 6792
rect 128728 6808 128780 6860
rect 129832 6808 129884 6860
rect 130936 6808 130988 6860
rect 132776 6808 132828 6860
rect 138204 6808 138256 6860
rect 128176 6740 128228 6792
rect 129096 6740 129148 6792
rect 130200 6740 130252 6792
rect 133052 6740 133104 6792
rect 133788 6740 133840 6792
rect 91928 6647 91980 6656
rect 91928 6613 91937 6647
rect 91937 6613 91971 6647
rect 91971 6613 91980 6647
rect 91928 6604 91980 6613
rect 92572 6604 92624 6656
rect 93400 6604 93452 6656
rect 96896 6604 96948 6656
rect 97356 6604 97408 6656
rect 106372 6604 106424 6656
rect 107016 6647 107068 6656
rect 107016 6613 107025 6647
rect 107025 6613 107059 6647
rect 107059 6613 107068 6647
rect 107016 6604 107068 6613
rect 115020 6604 115072 6656
rect 118148 6604 118200 6656
rect 120172 6604 120224 6656
rect 121092 6604 121144 6656
rect 121552 6604 121604 6656
rect 121644 6604 121696 6656
rect 123300 6604 123352 6656
rect 129372 6672 129424 6724
rect 125416 6647 125468 6656
rect 125416 6613 125425 6647
rect 125425 6613 125459 6647
rect 125459 6613 125468 6647
rect 125416 6604 125468 6613
rect 125968 6647 126020 6656
rect 125968 6613 125977 6647
rect 125977 6613 126011 6647
rect 126011 6613 126020 6647
rect 125968 6604 126020 6613
rect 126152 6604 126204 6656
rect 126520 6647 126572 6656
rect 126520 6613 126529 6647
rect 126529 6613 126563 6647
rect 126563 6613 126572 6647
rect 126520 6604 126572 6613
rect 127808 6604 127860 6656
rect 128360 6647 128412 6656
rect 128360 6613 128369 6647
rect 128369 6613 128403 6647
rect 128403 6613 128412 6647
rect 128360 6604 128412 6613
rect 129280 6604 129332 6656
rect 133236 6672 133288 6724
rect 133328 6672 133380 6724
rect 134156 6672 134208 6724
rect 133420 6604 133472 6656
rect 133696 6604 133748 6656
rect 135812 6740 135864 6792
rect 136640 6740 136692 6792
rect 139676 6740 139728 6792
rect 135076 6672 135128 6724
rect 135168 6647 135220 6656
rect 135168 6613 135177 6647
rect 135177 6613 135211 6647
rect 135211 6613 135220 6647
rect 135168 6604 135220 6613
rect 139584 6672 139636 6724
rect 142344 6808 142396 6860
rect 142620 6808 142672 6860
rect 147036 6944 147088 6996
rect 146484 6876 146536 6928
rect 148140 6876 148192 6928
rect 148508 6808 148560 6860
rect 150072 6944 150124 6996
rect 149704 6876 149756 6928
rect 151452 6919 151504 6928
rect 150440 6808 150492 6860
rect 151452 6885 151461 6919
rect 151461 6885 151495 6919
rect 151495 6885 151504 6919
rect 151452 6876 151504 6885
rect 152832 6876 152884 6928
rect 153752 6876 153804 6928
rect 152188 6808 152240 6860
rect 140136 6783 140188 6792
rect 140136 6749 140145 6783
rect 140145 6749 140179 6783
rect 140179 6749 140188 6783
rect 140136 6740 140188 6749
rect 142804 6740 142856 6792
rect 143080 6740 143132 6792
rect 143448 6740 143500 6792
rect 146392 6740 146444 6792
rect 146576 6740 146628 6792
rect 139492 6604 139544 6656
rect 139860 6604 139912 6656
rect 140780 6647 140832 6656
rect 140780 6613 140789 6647
rect 140789 6613 140823 6647
rect 140823 6613 140832 6647
rect 140780 6604 140832 6613
rect 143080 6604 143132 6656
rect 145288 6672 145340 6724
rect 146300 6672 146352 6724
rect 147312 6604 147364 6656
rect 147680 6740 147732 6792
rect 149704 6740 149756 6792
rect 150256 6740 150308 6792
rect 151268 6740 151320 6792
rect 151728 6740 151780 6792
rect 152096 6740 152148 6792
rect 152832 6740 152884 6792
rect 155224 6808 155276 6860
rect 155408 6808 155460 6860
rect 156788 6808 156840 6860
rect 155500 6783 155552 6792
rect 147588 6604 147640 6656
rect 147772 6604 147824 6656
rect 150164 6604 150216 6656
rect 150440 6604 150492 6656
rect 152188 6672 152240 6724
rect 152832 6647 152884 6656
rect 152832 6613 152841 6647
rect 152841 6613 152875 6647
rect 152875 6613 152884 6647
rect 152832 6604 152884 6613
rect 153476 6647 153528 6656
rect 153476 6613 153485 6647
rect 153485 6613 153519 6647
rect 153519 6613 153528 6647
rect 153476 6604 153528 6613
rect 154580 6715 154632 6724
rect 154580 6681 154620 6715
rect 154620 6681 154632 6715
rect 154580 6672 154632 6681
rect 155500 6749 155509 6783
rect 155509 6749 155543 6783
rect 155543 6749 155552 6783
rect 155500 6740 155552 6749
rect 156052 6740 156104 6792
rect 157064 6740 157116 6792
rect 157892 6740 157944 6792
rect 157708 6672 157760 6724
rect 155960 6604 156012 6656
rect 157616 6647 157668 6656
rect 157616 6613 157625 6647
rect 157625 6613 157659 6647
rect 157659 6613 157668 6647
rect 157616 6604 157668 6613
rect 40394 6502 40446 6554
rect 40458 6502 40510 6554
rect 40522 6502 40574 6554
rect 40586 6502 40638 6554
rect 40650 6502 40702 6554
rect 79839 6502 79891 6554
rect 79903 6502 79955 6554
rect 79967 6502 80019 6554
rect 80031 6502 80083 6554
rect 80095 6502 80147 6554
rect 119284 6502 119336 6554
rect 119348 6502 119400 6554
rect 119412 6502 119464 6554
rect 119476 6502 119528 6554
rect 119540 6502 119592 6554
rect 158729 6502 158781 6554
rect 158793 6502 158845 6554
rect 158857 6502 158909 6554
rect 158921 6502 158973 6554
rect 158985 6502 159037 6554
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 14924 6400 14976 6452
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 17500 6332 17552 6384
rect 18880 6400 18932 6452
rect 20076 6400 20128 6452
rect 20260 6400 20312 6452
rect 21272 6443 21324 6452
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 21456 6400 21508 6452
rect 23756 6400 23808 6452
rect 14004 6307 14056 6316
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 11152 6196 11204 6248
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 15016 6264 15068 6316
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 15660 6264 15712 6316
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 20996 6332 21048 6384
rect 17040 6264 17092 6273
rect 18052 6264 18104 6316
rect 18788 6264 18840 6316
rect 17500 6196 17552 6248
rect 18512 6196 18564 6248
rect 9312 6128 9364 6180
rect 15292 6128 15344 6180
rect 6000 6060 6052 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 12256 6060 12308 6112
rect 17040 6060 17092 6112
rect 17684 6060 17736 6112
rect 19340 6128 19392 6180
rect 20352 6196 20404 6248
rect 21640 6264 21692 6316
rect 23940 6332 23992 6384
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 37464 6400 37516 6452
rect 37556 6400 37608 6452
rect 38384 6400 38436 6452
rect 41236 6400 41288 6452
rect 27620 6332 27672 6384
rect 36360 6332 36412 6384
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 23296 6128 23348 6180
rect 30196 6264 30248 6316
rect 32404 6264 32456 6316
rect 38476 6264 38528 6316
rect 38660 6307 38712 6316
rect 38660 6273 38694 6307
rect 38694 6273 38712 6307
rect 40224 6307 40276 6316
rect 38660 6264 38712 6273
rect 40224 6273 40233 6307
rect 40233 6273 40267 6307
rect 40267 6273 40276 6307
rect 40224 6264 40276 6273
rect 40868 6332 40920 6384
rect 44732 6400 44784 6452
rect 46020 6400 46072 6452
rect 46572 6400 46624 6452
rect 52368 6400 52420 6452
rect 53196 6443 53248 6452
rect 53196 6409 53205 6443
rect 53205 6409 53239 6443
rect 53239 6409 53248 6443
rect 53196 6400 53248 6409
rect 26332 6196 26384 6248
rect 29368 6171 29420 6180
rect 29368 6137 29377 6171
rect 29377 6137 29411 6171
rect 29411 6137 29420 6171
rect 29368 6128 29420 6137
rect 33784 6239 33836 6248
rect 33784 6205 33793 6239
rect 33793 6205 33827 6239
rect 33827 6205 33836 6239
rect 33784 6196 33836 6205
rect 43536 6264 43588 6316
rect 40960 6196 41012 6248
rect 50712 6332 50764 6384
rect 33968 6128 34020 6180
rect 38016 6128 38068 6180
rect 19984 6060 20036 6112
rect 20260 6060 20312 6112
rect 22192 6060 22244 6112
rect 22376 6103 22428 6112
rect 22376 6069 22385 6103
rect 22385 6069 22419 6103
rect 22419 6069 22428 6103
rect 22376 6060 22428 6069
rect 23756 6060 23808 6112
rect 30840 6060 30892 6112
rect 33508 6060 33560 6112
rect 34980 6060 35032 6112
rect 41236 6128 41288 6180
rect 45928 6264 45980 6316
rect 46664 6307 46716 6316
rect 46020 6239 46072 6248
rect 46020 6205 46029 6239
rect 46029 6205 46063 6239
rect 46063 6205 46072 6239
rect 46020 6196 46072 6205
rect 46664 6273 46673 6307
rect 46673 6273 46707 6307
rect 46707 6273 46716 6307
rect 46664 6264 46716 6273
rect 50804 6264 50856 6316
rect 48596 6196 48648 6248
rect 51816 6332 51868 6384
rect 59728 6443 59780 6452
rect 59728 6409 59737 6443
rect 59737 6409 59771 6443
rect 59771 6409 59780 6443
rect 59728 6400 59780 6409
rect 63500 6400 63552 6452
rect 64052 6400 64104 6452
rect 64420 6400 64472 6452
rect 65892 6400 65944 6452
rect 66076 6443 66128 6452
rect 66076 6409 66085 6443
rect 66085 6409 66119 6443
rect 66119 6409 66128 6443
rect 66076 6400 66128 6409
rect 66536 6400 66588 6452
rect 69112 6400 69164 6452
rect 72884 6443 72936 6452
rect 53380 6307 53432 6316
rect 53380 6273 53389 6307
rect 53389 6273 53423 6307
rect 53423 6273 53432 6307
rect 53380 6264 53432 6273
rect 68928 6332 68980 6384
rect 54116 6264 54168 6316
rect 55404 6264 55456 6316
rect 50252 6128 50304 6180
rect 46204 6060 46256 6112
rect 50804 6060 50856 6112
rect 54208 6128 54260 6180
rect 54852 6060 54904 6112
rect 63960 6128 64012 6180
rect 63500 6060 63552 6112
rect 68376 6264 68428 6316
rect 72884 6409 72893 6443
rect 72893 6409 72927 6443
rect 72927 6409 72936 6443
rect 72884 6400 72936 6409
rect 73804 6443 73856 6452
rect 73804 6409 73813 6443
rect 73813 6409 73847 6443
rect 73847 6409 73856 6443
rect 73804 6400 73856 6409
rect 75000 6443 75052 6452
rect 75000 6409 75009 6443
rect 75009 6409 75043 6443
rect 75043 6409 75052 6443
rect 75000 6400 75052 6409
rect 78864 6443 78916 6452
rect 78864 6409 78873 6443
rect 78873 6409 78907 6443
rect 78907 6409 78916 6443
rect 78864 6400 78916 6409
rect 79324 6400 79376 6452
rect 80612 6400 80664 6452
rect 81072 6400 81124 6452
rect 82636 6400 82688 6452
rect 85580 6400 85632 6452
rect 89444 6400 89496 6452
rect 92204 6400 92256 6452
rect 94504 6400 94556 6452
rect 102140 6400 102192 6452
rect 106464 6443 106516 6452
rect 106464 6409 106473 6443
rect 106473 6409 106507 6443
rect 106507 6409 106516 6443
rect 106464 6400 106516 6409
rect 108764 6443 108816 6452
rect 108764 6409 108773 6443
rect 108773 6409 108807 6443
rect 108807 6409 108816 6443
rect 108764 6400 108816 6409
rect 108856 6400 108908 6452
rect 111340 6400 111392 6452
rect 111616 6400 111668 6452
rect 117136 6443 117188 6452
rect 73896 6264 73948 6316
rect 75092 6264 75144 6316
rect 89628 6264 89680 6316
rect 91468 6307 91520 6316
rect 91468 6273 91477 6307
rect 91477 6273 91511 6307
rect 91511 6273 91520 6307
rect 91468 6264 91520 6273
rect 76472 6196 76524 6248
rect 77116 6196 77168 6248
rect 80428 6196 80480 6248
rect 81072 6196 81124 6248
rect 73712 6060 73764 6112
rect 79140 6128 79192 6180
rect 80704 6128 80756 6180
rect 85580 6060 85632 6112
rect 88432 6196 88484 6248
rect 89536 6239 89588 6248
rect 89536 6205 89545 6239
rect 89545 6205 89579 6239
rect 89579 6205 89588 6239
rect 89536 6196 89588 6205
rect 90548 6196 90600 6248
rect 93216 6264 93268 6316
rect 97356 6307 97408 6316
rect 97356 6273 97390 6307
rect 97390 6273 97408 6307
rect 97356 6264 97408 6273
rect 101588 6307 101640 6316
rect 101588 6273 101597 6307
rect 101597 6273 101631 6307
rect 101631 6273 101640 6307
rect 101588 6264 101640 6273
rect 101864 6307 101916 6316
rect 101864 6273 101873 6307
rect 101873 6273 101907 6307
rect 101907 6273 101916 6307
rect 101864 6264 101916 6273
rect 105176 6264 105228 6316
rect 107200 6332 107252 6384
rect 107844 6332 107896 6384
rect 110696 6375 110748 6384
rect 107016 6264 107068 6316
rect 107384 6307 107436 6316
rect 107384 6273 107393 6307
rect 107393 6273 107427 6307
rect 107427 6273 107436 6307
rect 107384 6264 107436 6273
rect 91836 6196 91888 6248
rect 94044 6196 94096 6248
rect 96620 6196 96672 6248
rect 100760 6196 100812 6248
rect 100852 6196 100904 6248
rect 106096 6196 106148 6248
rect 107108 6196 107160 6248
rect 110696 6341 110705 6375
rect 110705 6341 110739 6375
rect 110739 6341 110748 6375
rect 110696 6332 110748 6341
rect 111432 6332 111484 6384
rect 111984 6332 112036 6384
rect 117136 6409 117145 6443
rect 117145 6409 117179 6443
rect 117179 6409 117188 6443
rect 117136 6400 117188 6409
rect 120540 6400 120592 6452
rect 121644 6400 121696 6452
rect 93124 6060 93176 6112
rect 93860 6060 93912 6112
rect 94320 6060 94372 6112
rect 96620 6103 96672 6112
rect 96620 6069 96629 6103
rect 96629 6069 96663 6103
rect 96663 6069 96672 6103
rect 96620 6060 96672 6069
rect 105084 6128 105136 6180
rect 100944 6060 100996 6112
rect 114560 6264 114612 6316
rect 114928 6264 114980 6316
rect 115848 6307 115900 6316
rect 115848 6273 115866 6307
rect 115866 6273 115900 6307
rect 119068 6332 119120 6384
rect 121920 6400 121972 6452
rect 121828 6332 121880 6384
rect 122748 6332 122800 6384
rect 123852 6400 123904 6452
rect 126152 6400 126204 6452
rect 126704 6400 126756 6452
rect 127992 6400 128044 6452
rect 128544 6400 128596 6452
rect 129556 6443 129608 6452
rect 115848 6264 115900 6273
rect 122564 6264 122616 6316
rect 116124 6239 116176 6248
rect 116124 6205 116133 6239
rect 116133 6205 116167 6239
rect 116167 6205 116176 6239
rect 116124 6196 116176 6205
rect 111892 6060 111944 6112
rect 114652 6128 114704 6180
rect 113824 6103 113876 6112
rect 113824 6069 113833 6103
rect 113833 6069 113867 6103
rect 113867 6069 113876 6103
rect 113824 6060 113876 6069
rect 115848 6060 115900 6112
rect 119896 6196 119948 6248
rect 121828 6196 121880 6248
rect 124864 6264 124916 6316
rect 125232 6264 125284 6316
rect 128268 6332 128320 6384
rect 129556 6409 129565 6443
rect 129565 6409 129599 6443
rect 129599 6409 129608 6443
rect 129556 6400 129608 6409
rect 130200 6443 130252 6452
rect 130200 6409 130209 6443
rect 130209 6409 130243 6443
rect 130243 6409 130252 6443
rect 130200 6400 130252 6409
rect 130568 6332 130620 6384
rect 131580 6332 131632 6384
rect 123300 6196 123352 6248
rect 123944 6196 123996 6248
rect 116768 6128 116820 6180
rect 118240 6103 118292 6112
rect 118240 6069 118249 6103
rect 118249 6069 118283 6103
rect 118283 6069 118292 6103
rect 118240 6060 118292 6069
rect 119712 6060 119764 6112
rect 123116 6128 123168 6180
rect 123852 6128 123904 6180
rect 124404 6171 124456 6180
rect 124404 6137 124413 6171
rect 124413 6137 124447 6171
rect 124447 6137 124456 6171
rect 124404 6128 124456 6137
rect 124220 6060 124272 6112
rect 127532 6264 127584 6316
rect 129280 6264 129332 6316
rect 129372 6264 129424 6316
rect 135076 6400 135128 6452
rect 136916 6400 136968 6452
rect 134248 6375 134300 6384
rect 134248 6341 134257 6375
rect 134257 6341 134291 6375
rect 134291 6341 134300 6375
rect 134248 6332 134300 6341
rect 135904 6332 135956 6384
rect 138204 6332 138256 6384
rect 128084 6196 128136 6248
rect 128268 6196 128320 6248
rect 130844 6196 130896 6248
rect 126520 6128 126572 6180
rect 132224 6196 132276 6248
rect 132776 6196 132828 6248
rect 132960 6196 133012 6248
rect 133052 6196 133104 6248
rect 138664 6264 138716 6316
rect 139676 6400 139728 6452
rect 139860 6400 139912 6452
rect 143356 6400 143408 6452
rect 143908 6400 143960 6452
rect 145012 6400 145064 6452
rect 145656 6443 145708 6452
rect 145656 6409 145665 6443
rect 145665 6409 145699 6443
rect 145699 6409 145708 6443
rect 145656 6400 145708 6409
rect 146300 6400 146352 6452
rect 147588 6400 147640 6452
rect 148232 6400 148284 6452
rect 149152 6400 149204 6452
rect 149796 6400 149848 6452
rect 149888 6400 149940 6452
rect 150440 6400 150492 6452
rect 152924 6400 152976 6452
rect 141240 6375 141292 6384
rect 131580 6128 131632 6180
rect 141240 6341 141249 6375
rect 141249 6341 141283 6375
rect 141283 6341 141292 6375
rect 141240 6332 141292 6341
rect 141332 6332 141384 6384
rect 143724 6332 143776 6384
rect 143816 6332 143868 6384
rect 147864 6332 147916 6384
rect 142804 6307 142856 6316
rect 142804 6273 142813 6307
rect 142813 6273 142847 6307
rect 142847 6273 142856 6307
rect 142804 6264 142856 6273
rect 142896 6264 142948 6316
rect 144092 6264 144144 6316
rect 144736 6264 144788 6316
rect 144920 6264 144972 6316
rect 145656 6264 145708 6316
rect 145932 6264 145984 6316
rect 146944 6264 146996 6316
rect 147128 6264 147180 6316
rect 149152 6264 149204 6316
rect 149336 6307 149388 6316
rect 149336 6273 149345 6307
rect 149345 6273 149379 6307
rect 149379 6273 149388 6307
rect 149336 6264 149388 6273
rect 150256 6307 150308 6316
rect 150256 6273 150265 6307
rect 150265 6273 150299 6307
rect 150299 6273 150308 6307
rect 150256 6264 150308 6273
rect 151084 6264 151136 6316
rect 152372 6264 152424 6316
rect 153384 6264 153436 6316
rect 153752 6264 153804 6316
rect 154028 6264 154080 6316
rect 154488 6264 154540 6316
rect 157800 6332 157852 6384
rect 139676 6196 139728 6248
rect 140688 6196 140740 6248
rect 147036 6239 147088 6248
rect 138940 6128 138992 6180
rect 127624 6060 127676 6112
rect 128544 6103 128596 6112
rect 128544 6069 128553 6103
rect 128553 6069 128587 6103
rect 128587 6069 128596 6103
rect 128544 6060 128596 6069
rect 128728 6060 128780 6112
rect 131212 6060 131264 6112
rect 131488 6103 131540 6112
rect 131488 6069 131497 6103
rect 131497 6069 131531 6103
rect 131531 6069 131540 6103
rect 131488 6060 131540 6069
rect 132316 6060 132368 6112
rect 132960 6060 133012 6112
rect 135260 6060 135312 6112
rect 136088 6060 136140 6112
rect 136640 6060 136692 6112
rect 137928 6060 137980 6112
rect 139860 6060 139912 6112
rect 140044 6060 140096 6112
rect 140412 6060 140464 6112
rect 140596 6060 140648 6112
rect 147036 6205 147045 6239
rect 147045 6205 147079 6239
rect 147079 6205 147088 6239
rect 147036 6196 147088 6205
rect 145932 6128 145984 6180
rect 146392 6060 146444 6112
rect 147404 6060 147456 6112
rect 148508 6196 148560 6248
rect 152924 6196 152976 6248
rect 153476 6196 153528 6248
rect 148784 6128 148836 6180
rect 150072 6128 150124 6180
rect 151636 6171 151688 6180
rect 147772 6060 147824 6112
rect 149244 6060 149296 6112
rect 149520 6103 149572 6112
rect 149520 6069 149529 6103
rect 149529 6069 149563 6103
rect 149563 6069 149572 6103
rect 149520 6060 149572 6069
rect 150256 6060 150308 6112
rect 151636 6137 151645 6171
rect 151645 6137 151679 6171
rect 151679 6137 151688 6171
rect 151636 6128 151688 6137
rect 153936 6128 153988 6180
rect 156420 6264 156472 6316
rect 158444 6332 158496 6384
rect 158168 6264 158220 6316
rect 155224 6196 155276 6248
rect 156788 6196 156840 6248
rect 155316 6128 155368 6180
rect 152648 6060 152700 6112
rect 153660 6060 153712 6112
rect 154304 6060 154356 6112
rect 155868 6060 155920 6112
rect 156328 6103 156380 6112
rect 156328 6069 156337 6103
rect 156337 6069 156371 6103
rect 156371 6069 156380 6103
rect 156328 6060 156380 6069
rect 156788 6103 156840 6112
rect 156788 6069 156797 6103
rect 156797 6069 156831 6103
rect 156831 6069 156840 6103
rect 156788 6060 156840 6069
rect 157064 6060 157116 6112
rect 20672 5958 20724 6010
rect 20736 5958 20788 6010
rect 20800 5958 20852 6010
rect 20864 5958 20916 6010
rect 20928 5958 20980 6010
rect 60117 5958 60169 6010
rect 60181 5958 60233 6010
rect 60245 5958 60297 6010
rect 60309 5958 60361 6010
rect 60373 5958 60425 6010
rect 99562 5958 99614 6010
rect 99626 5958 99678 6010
rect 99690 5958 99742 6010
rect 99754 5958 99806 6010
rect 99818 5958 99870 6010
rect 139007 5958 139059 6010
rect 139071 5958 139123 6010
rect 139135 5958 139187 6010
rect 139199 5958 139251 6010
rect 139263 5958 139315 6010
rect 4896 5856 4948 5908
rect 5724 5856 5776 5908
rect 15200 5856 15252 5908
rect 16580 5856 16632 5908
rect 18144 5856 18196 5908
rect 18880 5856 18932 5908
rect 19524 5856 19576 5908
rect 20352 5856 20404 5908
rect 22008 5856 22060 5908
rect 22468 5856 22520 5908
rect 24032 5856 24084 5908
rect 24860 5856 24912 5908
rect 28908 5856 28960 5908
rect 30380 5856 30432 5908
rect 32312 5899 32364 5908
rect 17316 5788 17368 5840
rect 17500 5788 17552 5840
rect 30472 5788 30524 5840
rect 30564 5788 30616 5840
rect 32036 5788 32088 5840
rect 32312 5865 32321 5899
rect 32321 5865 32355 5899
rect 32355 5865 32364 5899
rect 32312 5856 32364 5865
rect 33784 5856 33836 5908
rect 33968 5788 34020 5840
rect 3884 5652 3936 5704
rect 4620 5652 4672 5704
rect 6092 5652 6144 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 20260 5720 20312 5772
rect 22008 5720 22060 5772
rect 25228 5720 25280 5772
rect 25780 5720 25832 5772
rect 38660 5856 38712 5908
rect 43260 5899 43312 5908
rect 43260 5865 43269 5899
rect 43269 5865 43303 5899
rect 43303 5865 43312 5899
rect 43260 5856 43312 5865
rect 44456 5856 44508 5908
rect 37464 5788 37516 5840
rect 43628 5788 43680 5840
rect 44640 5763 44692 5772
rect 14372 5584 14424 5636
rect 14464 5584 14516 5636
rect 15016 5584 15068 5636
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 17776 5652 17828 5704
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 19984 5652 20036 5704
rect 9680 5516 9732 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 15568 5516 15620 5568
rect 21088 5584 21140 5636
rect 22376 5652 22428 5704
rect 29000 5652 29052 5704
rect 30380 5695 30432 5704
rect 30380 5661 30389 5695
rect 30389 5661 30423 5695
rect 30423 5661 30432 5695
rect 30380 5652 30432 5661
rect 30472 5652 30524 5704
rect 34428 5652 34480 5704
rect 37832 5695 37884 5704
rect 23940 5584 23992 5636
rect 24032 5584 24084 5636
rect 33968 5584 34020 5636
rect 34336 5584 34388 5636
rect 37188 5584 37240 5636
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 16764 5516 16816 5568
rect 17040 5516 17092 5568
rect 18604 5516 18656 5568
rect 18696 5516 18748 5568
rect 22100 5516 22152 5568
rect 22192 5516 22244 5568
rect 26056 5516 26108 5568
rect 30380 5516 30432 5568
rect 33048 5516 33100 5568
rect 41236 5652 41288 5704
rect 44640 5729 44649 5763
rect 44649 5729 44683 5763
rect 44683 5729 44692 5763
rect 44640 5720 44692 5729
rect 48504 5856 48556 5908
rect 48596 5856 48648 5908
rect 59912 5856 59964 5908
rect 66628 5899 66680 5908
rect 47124 5788 47176 5840
rect 47308 5831 47360 5840
rect 47308 5797 47317 5831
rect 47317 5797 47351 5831
rect 47351 5797 47360 5831
rect 47308 5788 47360 5797
rect 49056 5788 49108 5840
rect 45836 5763 45888 5772
rect 45836 5729 45845 5763
rect 45845 5729 45879 5763
rect 45879 5729 45888 5763
rect 45836 5720 45888 5729
rect 46020 5720 46072 5772
rect 54668 5763 54720 5772
rect 54668 5729 54677 5763
rect 54677 5729 54711 5763
rect 54711 5729 54720 5763
rect 54668 5720 54720 5729
rect 63316 5720 63368 5772
rect 66628 5865 66637 5899
rect 66637 5865 66671 5899
rect 66671 5865 66680 5899
rect 66628 5856 66680 5865
rect 68928 5899 68980 5908
rect 68928 5865 68937 5899
rect 68937 5865 68971 5899
rect 68971 5865 68980 5899
rect 68928 5856 68980 5865
rect 69296 5856 69348 5908
rect 75920 5856 75972 5908
rect 76748 5856 76800 5908
rect 90640 5856 90692 5908
rect 91836 5899 91888 5908
rect 91836 5865 91845 5899
rect 91845 5865 91879 5899
rect 91879 5865 91888 5899
rect 91836 5856 91888 5865
rect 67640 5788 67692 5840
rect 69112 5788 69164 5840
rect 72700 5831 72752 5840
rect 72700 5797 72709 5831
rect 72709 5797 72743 5831
rect 72743 5797 72752 5831
rect 72700 5788 72752 5797
rect 65892 5720 65944 5772
rect 76012 5720 76064 5772
rect 38016 5584 38068 5636
rect 38568 5559 38620 5568
rect 38568 5525 38577 5559
rect 38577 5525 38611 5559
rect 38611 5525 38620 5559
rect 38568 5516 38620 5525
rect 43628 5516 43680 5568
rect 47216 5516 47268 5568
rect 47308 5516 47360 5568
rect 54208 5695 54260 5704
rect 54208 5661 54217 5695
rect 54217 5661 54251 5695
rect 54251 5661 54260 5695
rect 58624 5695 58676 5704
rect 54208 5652 54260 5661
rect 58624 5661 58633 5695
rect 58633 5661 58667 5695
rect 58667 5661 58676 5695
rect 58624 5652 58676 5661
rect 63776 5652 63828 5704
rect 66076 5652 66128 5704
rect 66260 5652 66312 5704
rect 62028 5584 62080 5636
rect 69112 5584 69164 5636
rect 73160 5652 73212 5704
rect 74172 5652 74224 5704
rect 86408 5788 86460 5840
rect 93860 5788 93912 5840
rect 80428 5763 80480 5772
rect 80428 5729 80437 5763
rect 80437 5729 80471 5763
rect 80471 5729 80480 5763
rect 80428 5720 80480 5729
rect 76748 5695 76800 5704
rect 76748 5661 76757 5695
rect 76757 5661 76791 5695
rect 76791 5661 76800 5695
rect 76748 5652 76800 5661
rect 78864 5652 78916 5704
rect 81256 5695 81308 5704
rect 81256 5661 81265 5695
rect 81265 5661 81299 5695
rect 81299 5661 81308 5695
rect 81256 5652 81308 5661
rect 83280 5652 83332 5704
rect 96620 5856 96672 5908
rect 101312 5856 101364 5908
rect 103428 5856 103480 5908
rect 108856 5899 108908 5908
rect 99932 5788 99984 5840
rect 105084 5788 105136 5840
rect 106648 5788 106700 5840
rect 108856 5865 108865 5899
rect 108865 5865 108899 5899
rect 108899 5865 108908 5899
rect 108856 5856 108908 5865
rect 116768 5856 116820 5908
rect 117412 5899 117464 5908
rect 117412 5865 117421 5899
rect 117421 5865 117455 5899
rect 117455 5865 117464 5899
rect 117412 5856 117464 5865
rect 101496 5720 101548 5772
rect 106096 5720 106148 5772
rect 114560 5788 114612 5840
rect 115388 5831 115440 5840
rect 115388 5797 115397 5831
rect 115397 5797 115431 5831
rect 115431 5797 115440 5831
rect 115388 5788 115440 5797
rect 117044 5788 117096 5840
rect 120540 5856 120592 5908
rect 120816 5899 120868 5908
rect 120816 5865 120825 5899
rect 120825 5865 120859 5899
rect 120859 5865 120868 5899
rect 120816 5856 120868 5865
rect 121920 5856 121972 5908
rect 122472 5899 122524 5908
rect 122472 5865 122481 5899
rect 122481 5865 122515 5899
rect 122515 5865 122524 5899
rect 122472 5856 122524 5865
rect 122564 5856 122616 5908
rect 127532 5856 127584 5908
rect 108488 5720 108540 5772
rect 117136 5720 117188 5772
rect 95332 5695 95384 5704
rect 74448 5584 74500 5636
rect 77208 5584 77260 5636
rect 94136 5584 94188 5636
rect 95332 5661 95341 5695
rect 95341 5661 95375 5695
rect 95375 5661 95384 5695
rect 95332 5652 95384 5661
rect 101312 5695 101364 5704
rect 58440 5559 58492 5568
rect 58440 5525 58449 5559
rect 58449 5525 58483 5559
rect 58483 5525 58492 5559
rect 58440 5516 58492 5525
rect 65800 5559 65852 5568
rect 65800 5525 65809 5559
rect 65809 5525 65843 5559
rect 65843 5525 65852 5559
rect 65800 5516 65852 5525
rect 75368 5516 75420 5568
rect 76012 5516 76064 5568
rect 93400 5559 93452 5568
rect 93400 5525 93409 5559
rect 93409 5525 93443 5559
rect 93443 5525 93452 5559
rect 93400 5516 93452 5525
rect 93860 5516 93912 5568
rect 94044 5516 94096 5568
rect 100944 5584 100996 5636
rect 101312 5661 101321 5695
rect 101321 5661 101355 5695
rect 101355 5661 101364 5695
rect 101312 5652 101364 5661
rect 107660 5652 107712 5704
rect 113732 5652 113784 5704
rect 121736 5831 121788 5840
rect 121736 5797 121745 5831
rect 121745 5797 121779 5831
rect 121779 5797 121788 5831
rect 121736 5788 121788 5797
rect 126520 5788 126572 5840
rect 127072 5831 127124 5840
rect 127072 5797 127081 5831
rect 127081 5797 127115 5831
rect 127115 5797 127124 5831
rect 127072 5788 127124 5797
rect 123024 5720 123076 5772
rect 123944 5720 123996 5772
rect 124956 5720 125008 5772
rect 128360 5856 128412 5908
rect 129648 5856 129700 5908
rect 132868 5899 132920 5908
rect 132868 5865 132877 5899
rect 132877 5865 132911 5899
rect 132911 5865 132920 5899
rect 132868 5856 132920 5865
rect 133972 5856 134024 5908
rect 135260 5856 135312 5908
rect 135720 5899 135772 5908
rect 135720 5865 135729 5899
rect 135729 5865 135763 5899
rect 135763 5865 135772 5899
rect 135720 5856 135772 5865
rect 136272 5899 136324 5908
rect 136272 5865 136281 5899
rect 136281 5865 136315 5899
rect 136315 5865 136324 5899
rect 136272 5856 136324 5865
rect 137008 5856 137060 5908
rect 118608 5652 118660 5704
rect 118976 5695 119028 5704
rect 118976 5661 118985 5695
rect 118985 5661 119019 5695
rect 119019 5661 119028 5695
rect 118976 5652 119028 5661
rect 99932 5559 99984 5568
rect 99932 5525 99941 5559
rect 99941 5525 99975 5559
rect 99975 5525 99984 5559
rect 99932 5516 99984 5525
rect 101956 5559 102008 5568
rect 101956 5525 101965 5559
rect 101965 5525 101999 5559
rect 101999 5525 102008 5559
rect 101956 5516 102008 5525
rect 107384 5584 107436 5636
rect 112168 5584 112220 5636
rect 117412 5584 117464 5636
rect 108028 5516 108080 5568
rect 113548 5516 113600 5568
rect 113732 5516 113784 5568
rect 121184 5695 121236 5704
rect 121184 5661 121193 5695
rect 121193 5661 121227 5695
rect 121227 5661 121236 5695
rect 121184 5652 121236 5661
rect 121736 5652 121788 5704
rect 125784 5695 125836 5704
rect 121368 5516 121420 5568
rect 125784 5661 125793 5695
rect 125793 5661 125827 5695
rect 125827 5661 125836 5695
rect 125784 5652 125836 5661
rect 126060 5652 126112 5704
rect 127624 5695 127676 5704
rect 123024 5584 123076 5636
rect 122564 5516 122616 5568
rect 124588 5516 124640 5568
rect 125048 5559 125100 5568
rect 125048 5525 125057 5559
rect 125057 5525 125091 5559
rect 125091 5525 125100 5559
rect 125048 5516 125100 5525
rect 125416 5584 125468 5636
rect 127624 5661 127633 5695
rect 127633 5661 127667 5695
rect 127667 5661 127676 5695
rect 127624 5652 127676 5661
rect 127900 5695 127952 5704
rect 127900 5661 127934 5695
rect 127934 5661 127952 5695
rect 127900 5652 127952 5661
rect 129096 5788 129148 5840
rect 141332 5856 141384 5908
rect 144920 5856 144972 5908
rect 145288 5856 145340 5908
rect 137284 5831 137336 5840
rect 131212 5720 131264 5772
rect 132316 5720 132368 5772
rect 132960 5720 133012 5772
rect 137284 5797 137293 5831
rect 137293 5797 137327 5831
rect 137327 5797 137336 5831
rect 137284 5788 137336 5797
rect 138296 5788 138348 5840
rect 140044 5788 140096 5840
rect 144184 5788 144236 5840
rect 137008 5720 137060 5772
rect 138848 5720 138900 5772
rect 130108 5652 130160 5704
rect 130844 5652 130896 5704
rect 133972 5695 134024 5704
rect 133972 5661 133981 5695
rect 133981 5661 134015 5695
rect 134015 5661 134024 5695
rect 133972 5652 134024 5661
rect 134524 5695 134576 5704
rect 134524 5661 134533 5695
rect 134533 5661 134567 5695
rect 134567 5661 134576 5695
rect 134524 5652 134576 5661
rect 130200 5627 130252 5636
rect 125692 5516 125744 5568
rect 126244 5516 126296 5568
rect 126704 5516 126756 5568
rect 130200 5593 130209 5627
rect 130209 5593 130243 5627
rect 130243 5593 130252 5627
rect 130200 5584 130252 5593
rect 131304 5627 131356 5636
rect 131304 5593 131313 5627
rect 131313 5593 131347 5627
rect 131347 5593 131356 5627
rect 131304 5584 131356 5593
rect 131948 5627 132000 5636
rect 131948 5593 131957 5627
rect 131957 5593 131991 5627
rect 131991 5593 132000 5627
rect 131948 5584 132000 5593
rect 136640 5652 136692 5704
rect 137928 5652 137980 5704
rect 139308 5652 139360 5704
rect 140504 5695 140556 5704
rect 140504 5661 140513 5695
rect 140513 5661 140547 5695
rect 140547 5661 140556 5695
rect 140504 5652 140556 5661
rect 144092 5720 144144 5772
rect 147680 5856 147732 5908
rect 156788 5856 156840 5908
rect 149428 5788 149480 5840
rect 149888 5788 149940 5840
rect 150624 5788 150676 5840
rect 152372 5788 152424 5840
rect 153936 5788 153988 5840
rect 154120 5788 154172 5840
rect 142436 5652 142488 5704
rect 142804 5652 142856 5704
rect 149244 5720 149296 5772
rect 128544 5516 128596 5568
rect 131028 5516 131080 5568
rect 133052 5516 133104 5568
rect 135536 5584 135588 5636
rect 136916 5584 136968 5636
rect 140044 5584 140096 5636
rect 140780 5584 140832 5636
rect 143356 5627 143408 5636
rect 143356 5593 143390 5627
rect 143390 5593 143408 5627
rect 143356 5584 143408 5593
rect 146208 5584 146260 5636
rect 146392 5652 146444 5704
rect 146760 5695 146812 5704
rect 146760 5661 146769 5695
rect 146769 5661 146803 5695
rect 146803 5661 146812 5695
rect 146760 5652 146812 5661
rect 146944 5695 146996 5704
rect 146944 5661 146953 5695
rect 146953 5661 146987 5695
rect 146987 5661 146996 5695
rect 146944 5652 146996 5661
rect 147036 5652 147088 5704
rect 147404 5652 147456 5704
rect 148876 5652 148928 5704
rect 149520 5652 149572 5704
rect 153108 5720 153160 5772
rect 153200 5720 153252 5772
rect 151544 5652 151596 5704
rect 151912 5652 151964 5704
rect 153568 5652 153620 5704
rect 153660 5695 153712 5704
rect 153660 5661 153669 5695
rect 153669 5661 153703 5695
rect 153703 5661 153712 5695
rect 153660 5652 153712 5661
rect 154120 5652 154172 5704
rect 154488 5788 154540 5840
rect 154948 5788 155000 5840
rect 156696 5788 156748 5840
rect 157248 5788 157300 5840
rect 158260 5720 158312 5772
rect 133788 5516 133840 5568
rect 136272 5516 136324 5568
rect 138664 5516 138716 5568
rect 142620 5516 142672 5568
rect 143080 5516 143132 5568
rect 146668 5516 146720 5568
rect 147404 5516 147456 5568
rect 148324 5516 148376 5568
rect 151452 5584 151504 5636
rect 154672 5695 154724 5704
rect 154672 5661 154681 5695
rect 154681 5661 154715 5695
rect 154715 5661 154724 5695
rect 155500 5695 155552 5704
rect 154672 5652 154724 5661
rect 155500 5661 155509 5695
rect 155509 5661 155543 5695
rect 155543 5661 155552 5695
rect 155500 5652 155552 5661
rect 149428 5516 149480 5568
rect 149704 5516 149756 5568
rect 150164 5516 150216 5568
rect 151084 5516 151136 5568
rect 155408 5584 155460 5636
rect 155776 5652 155828 5704
rect 157156 5695 157208 5704
rect 155868 5584 155920 5636
rect 157156 5661 157165 5695
rect 157165 5661 157199 5695
rect 157199 5661 157208 5695
rect 157156 5652 157208 5661
rect 157524 5652 157576 5704
rect 158628 5516 158680 5568
rect 40394 5414 40446 5466
rect 40458 5414 40510 5466
rect 40522 5414 40574 5466
rect 40586 5414 40638 5466
rect 40650 5414 40702 5466
rect 79839 5414 79891 5466
rect 79903 5414 79955 5466
rect 79967 5414 80019 5466
rect 80031 5414 80083 5466
rect 80095 5414 80147 5466
rect 119284 5414 119336 5466
rect 119348 5414 119400 5466
rect 119412 5414 119464 5466
rect 119476 5414 119528 5466
rect 119540 5414 119592 5466
rect 158729 5414 158781 5466
rect 158793 5414 158845 5466
rect 158857 5414 158909 5466
rect 158921 5414 158973 5466
rect 158985 5414 159037 5466
rect 5908 5312 5960 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 13728 5312 13780 5364
rect 13820 5312 13872 5364
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 16764 5312 16816 5364
rect 18144 5355 18196 5364
rect 18144 5321 18153 5355
rect 18153 5321 18187 5355
rect 18187 5321 18196 5355
rect 18144 5312 18196 5321
rect 18696 5312 18748 5364
rect 19892 5355 19944 5364
rect 19892 5321 19901 5355
rect 19901 5321 19935 5355
rect 19935 5321 19944 5355
rect 19892 5312 19944 5321
rect 3884 5244 3936 5296
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6000 5176 6052 5228
rect 14280 5244 14332 5296
rect 16948 5244 17000 5296
rect 12992 5176 13044 5228
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 9680 5108 9732 5160
rect 13636 5108 13688 5160
rect 17224 5176 17276 5228
rect 21364 5244 21416 5296
rect 23020 5287 23072 5296
rect 23020 5253 23054 5287
rect 23054 5253 23072 5287
rect 25504 5312 25556 5364
rect 25964 5312 26016 5364
rect 23020 5244 23072 5253
rect 34520 5312 34572 5364
rect 35348 5355 35400 5364
rect 35348 5321 35357 5355
rect 35357 5321 35391 5355
rect 35391 5321 35400 5355
rect 35348 5312 35400 5321
rect 43352 5312 43404 5364
rect 55036 5312 55088 5364
rect 62396 5355 62448 5364
rect 62396 5321 62405 5355
rect 62405 5321 62439 5355
rect 62439 5321 62448 5355
rect 62396 5312 62448 5321
rect 63316 5355 63368 5364
rect 63316 5321 63325 5355
rect 63325 5321 63359 5355
rect 63359 5321 63368 5355
rect 63316 5312 63368 5321
rect 65892 5312 65944 5364
rect 73160 5312 73212 5364
rect 74356 5312 74408 5364
rect 75920 5355 75972 5364
rect 75920 5321 75929 5355
rect 75929 5321 75963 5355
rect 75963 5321 75972 5355
rect 75920 5312 75972 5321
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 12624 4972 12676 5024
rect 14280 4972 14332 5024
rect 14924 4972 14976 5024
rect 15568 5108 15620 5160
rect 15844 5108 15896 5160
rect 22468 5108 22520 5160
rect 24676 5176 24728 5228
rect 32312 5244 32364 5296
rect 33784 5244 33836 5296
rect 45376 5287 45428 5296
rect 30472 5176 30524 5228
rect 35992 5176 36044 5228
rect 36636 5176 36688 5228
rect 45376 5253 45385 5287
rect 45385 5253 45419 5287
rect 45419 5253 45428 5287
rect 45376 5244 45428 5253
rect 45836 5244 45888 5296
rect 48320 5244 48372 5296
rect 38568 5176 38620 5228
rect 48688 5219 48740 5228
rect 48688 5185 48697 5219
rect 48697 5185 48731 5219
rect 48731 5185 48740 5219
rect 48688 5176 48740 5185
rect 58808 5176 58860 5228
rect 63592 5244 63644 5296
rect 61108 5176 61160 5228
rect 61752 5176 61804 5228
rect 74816 5176 74868 5228
rect 76012 5244 76064 5296
rect 114100 5312 114152 5364
rect 116032 5312 116084 5364
rect 118424 5312 118476 5364
rect 118700 5312 118752 5364
rect 118884 5312 118936 5364
rect 122656 5312 122708 5364
rect 123116 5355 123168 5364
rect 123116 5321 123125 5355
rect 123125 5321 123159 5355
rect 123159 5321 123168 5355
rect 123116 5312 123168 5321
rect 125508 5312 125560 5364
rect 126796 5312 126848 5364
rect 127808 5312 127860 5364
rect 128084 5312 128136 5364
rect 128360 5312 128412 5364
rect 129188 5312 129240 5364
rect 129740 5312 129792 5364
rect 129832 5312 129884 5364
rect 137376 5312 137428 5364
rect 137836 5355 137888 5364
rect 137836 5321 137845 5355
rect 137845 5321 137879 5355
rect 137879 5321 137888 5355
rect 137836 5312 137888 5321
rect 138388 5355 138440 5364
rect 138388 5321 138397 5355
rect 138397 5321 138431 5355
rect 138431 5321 138440 5355
rect 138388 5312 138440 5321
rect 139308 5355 139360 5364
rect 139308 5321 139317 5355
rect 139317 5321 139351 5355
rect 139351 5321 139360 5355
rect 139308 5312 139360 5321
rect 141516 5312 141568 5364
rect 142712 5312 142764 5364
rect 144644 5355 144696 5364
rect 81256 5244 81308 5296
rect 81072 5176 81124 5228
rect 17224 5040 17276 5092
rect 21916 5040 21968 5092
rect 22560 5040 22612 5092
rect 30288 5108 30340 5160
rect 31760 5151 31812 5160
rect 31760 5117 31769 5151
rect 31769 5117 31803 5151
rect 31803 5117 31812 5151
rect 31760 5108 31812 5117
rect 34336 5108 34388 5160
rect 51080 5108 51132 5160
rect 52276 5108 52328 5160
rect 55404 5151 55456 5160
rect 34060 5083 34112 5092
rect 18236 4972 18288 5024
rect 22652 4972 22704 5024
rect 34060 5049 34069 5083
rect 34069 5049 34103 5083
rect 34103 5049 34112 5083
rect 34060 5040 34112 5049
rect 24676 4972 24728 5024
rect 25320 4972 25372 5024
rect 30380 5015 30432 5024
rect 30380 4981 30389 5015
rect 30389 4981 30423 5015
rect 30423 4981 30432 5015
rect 30380 4972 30432 4981
rect 55404 5117 55413 5151
rect 55413 5117 55447 5151
rect 55447 5117 55456 5151
rect 55404 5108 55456 5117
rect 75552 5108 75604 5160
rect 88340 5176 88392 5228
rect 92572 5176 92624 5228
rect 93400 5244 93452 5296
rect 95332 5244 95384 5296
rect 116952 5244 117004 5296
rect 117136 5244 117188 5296
rect 120172 5287 120224 5296
rect 93124 5219 93176 5228
rect 93124 5185 93133 5219
rect 93133 5185 93167 5219
rect 93167 5185 93176 5219
rect 93124 5176 93176 5185
rect 93216 5176 93268 5228
rect 96712 5176 96764 5228
rect 105176 5176 105228 5228
rect 109132 5176 109184 5228
rect 109776 5176 109828 5228
rect 113824 5176 113876 5228
rect 77208 5040 77260 5092
rect 83004 5108 83056 5160
rect 101312 5108 101364 5160
rect 104624 5151 104676 5160
rect 104624 5117 104633 5151
rect 104633 5117 104667 5151
rect 104667 5117 104676 5151
rect 104624 5108 104676 5117
rect 110880 5108 110932 5160
rect 88064 5040 88116 5092
rect 56784 5015 56836 5024
rect 56784 4981 56793 5015
rect 56793 4981 56827 5015
rect 56827 4981 56836 5015
rect 56784 4972 56836 4981
rect 81900 5015 81952 5024
rect 81900 4981 81909 5015
rect 81909 4981 81943 5015
rect 81943 4981 81952 5015
rect 81900 4972 81952 4981
rect 84292 4972 84344 5024
rect 91100 4972 91152 5024
rect 94136 5040 94188 5092
rect 111892 5040 111944 5092
rect 113548 5108 113600 5160
rect 118056 5176 118108 5228
rect 118332 5176 118384 5228
rect 120172 5253 120206 5287
rect 120206 5253 120224 5287
rect 120172 5244 120224 5253
rect 121828 5244 121880 5296
rect 125048 5244 125100 5296
rect 127072 5244 127124 5296
rect 132040 5287 132092 5296
rect 132040 5253 132049 5287
rect 132049 5253 132083 5287
rect 132083 5253 132092 5287
rect 132040 5244 132092 5253
rect 137192 5244 137244 5296
rect 137284 5244 137336 5296
rect 116032 5108 116084 5160
rect 117780 5108 117832 5160
rect 117872 5108 117924 5160
rect 124220 5176 124272 5228
rect 126704 5176 126756 5228
rect 127164 5219 127216 5228
rect 121736 5151 121788 5160
rect 121736 5117 121745 5151
rect 121745 5117 121779 5151
rect 121779 5117 121788 5151
rect 121736 5108 121788 5117
rect 125048 5151 125100 5160
rect 125048 5117 125057 5151
rect 125057 5117 125091 5151
rect 125091 5117 125100 5151
rect 125048 5108 125100 5117
rect 125140 5108 125192 5160
rect 127164 5185 127173 5219
rect 127173 5185 127207 5219
rect 127207 5185 127216 5219
rect 127164 5176 127216 5185
rect 128084 5219 128136 5228
rect 128084 5185 128093 5219
rect 128093 5185 128127 5219
rect 128127 5185 128136 5219
rect 128084 5176 128136 5185
rect 131396 5219 131448 5228
rect 131396 5185 131405 5219
rect 131405 5185 131439 5219
rect 131439 5185 131448 5219
rect 131396 5176 131448 5185
rect 131488 5176 131540 5228
rect 134800 5176 134852 5228
rect 136824 5219 136876 5228
rect 136824 5185 136833 5219
rect 136833 5185 136867 5219
rect 136867 5185 136876 5219
rect 136824 5176 136876 5185
rect 136916 5176 136968 5228
rect 140228 5244 140280 5296
rect 138572 5219 138624 5228
rect 138572 5185 138581 5219
rect 138581 5185 138615 5219
rect 138615 5185 138624 5219
rect 138572 5176 138624 5185
rect 139768 5219 139820 5228
rect 139768 5185 139777 5219
rect 139777 5185 139811 5219
rect 139811 5185 139820 5219
rect 139768 5176 139820 5185
rect 139860 5176 139912 5228
rect 140044 5176 140096 5228
rect 141148 5176 141200 5228
rect 115848 5040 115900 5092
rect 118148 5040 118200 5092
rect 119068 5040 119120 5092
rect 122840 5040 122892 5092
rect 125876 5040 125928 5092
rect 112168 5015 112220 5024
rect 112168 4981 112177 5015
rect 112177 4981 112211 5015
rect 112211 4981 112220 5015
rect 112168 4972 112220 4981
rect 115480 4972 115532 5024
rect 119252 5015 119304 5024
rect 119252 4981 119261 5015
rect 119261 4981 119295 5015
rect 119295 4981 119304 5015
rect 119252 4972 119304 4981
rect 124036 4972 124088 5024
rect 125416 4972 125468 5024
rect 126520 4972 126572 5024
rect 127992 5108 128044 5160
rect 126796 5040 126848 5092
rect 129740 5108 129792 5160
rect 131672 5108 131724 5160
rect 132500 5108 132552 5160
rect 140964 5108 141016 5160
rect 142804 5244 142856 5296
rect 142344 5176 142396 5228
rect 144644 5321 144653 5355
rect 144653 5321 144687 5355
rect 144687 5321 144696 5355
rect 144644 5312 144696 5321
rect 145564 5312 145616 5364
rect 146760 5312 146812 5364
rect 147588 5312 147640 5364
rect 144184 5244 144236 5296
rect 147312 5244 147364 5296
rect 147680 5244 147732 5296
rect 150256 5244 150308 5296
rect 150348 5244 150400 5296
rect 151820 5244 151872 5296
rect 155868 5312 155920 5364
rect 156788 5355 156840 5364
rect 156788 5321 156797 5355
rect 156797 5321 156831 5355
rect 156831 5321 156840 5355
rect 156788 5312 156840 5321
rect 157156 5312 157208 5364
rect 145288 5176 145340 5228
rect 146944 5176 146996 5228
rect 147036 5219 147088 5228
rect 147036 5185 147045 5219
rect 147045 5185 147079 5219
rect 147079 5185 147088 5219
rect 147036 5176 147088 5185
rect 135720 5083 135772 5092
rect 130844 5015 130896 5024
rect 130844 4981 130853 5015
rect 130853 4981 130887 5015
rect 130887 4981 130896 5015
rect 130844 4972 130896 4981
rect 132316 4972 132368 5024
rect 133052 5015 133104 5024
rect 133052 4981 133061 5015
rect 133061 4981 133095 5015
rect 133095 4981 133104 5015
rect 135720 5049 135729 5083
rect 135729 5049 135763 5083
rect 135763 5049 135772 5083
rect 135720 5040 135772 5049
rect 140596 5083 140648 5092
rect 133052 4972 133104 4981
rect 134800 5015 134852 5024
rect 134800 4981 134809 5015
rect 134809 4981 134843 5015
rect 134843 4981 134852 5015
rect 134800 4972 134852 4981
rect 136916 4972 136968 5024
rect 137560 4972 137612 5024
rect 140596 5049 140605 5083
rect 140605 5049 140639 5083
rect 140639 5049 140648 5083
rect 140596 5040 140648 5049
rect 139584 4972 139636 5024
rect 139768 4972 139820 5024
rect 142712 4972 142764 5024
rect 145932 5108 145984 5160
rect 148876 5219 148928 5228
rect 148876 5185 148885 5219
rect 148885 5185 148919 5219
rect 148919 5185 148928 5219
rect 148876 5176 148928 5185
rect 149336 5176 149388 5228
rect 149796 5176 149848 5228
rect 154304 5244 154356 5296
rect 152372 5176 152424 5228
rect 154028 5176 154080 5228
rect 147128 5040 147180 5092
rect 145288 4972 145340 5024
rect 145656 4972 145708 5024
rect 147312 4972 147364 5024
rect 150348 5040 150400 5092
rect 149704 4972 149756 5024
rect 150808 5015 150860 5024
rect 150808 4981 150817 5015
rect 150817 4981 150851 5015
rect 150851 4981 150860 5015
rect 150808 4972 150860 4981
rect 152188 5151 152240 5160
rect 152188 5117 152197 5151
rect 152197 5117 152231 5151
rect 152231 5117 152240 5151
rect 152648 5151 152700 5160
rect 152188 5108 152240 5117
rect 152648 5117 152657 5151
rect 152657 5117 152691 5151
rect 152691 5117 152700 5151
rect 152648 5108 152700 5117
rect 153384 5108 153436 5160
rect 154120 5108 154172 5160
rect 154672 5219 154724 5228
rect 154672 5185 154681 5219
rect 154681 5185 154715 5219
rect 154715 5185 154724 5219
rect 154672 5176 154724 5185
rect 159180 5244 159232 5296
rect 155776 5176 155828 5228
rect 152556 5040 152608 5092
rect 155316 5040 155368 5092
rect 155500 5040 155552 5092
rect 156604 5176 156656 5228
rect 157340 5176 157392 5228
rect 158536 5176 158588 5228
rect 153016 4972 153068 5024
rect 154120 4972 154172 5024
rect 154672 4972 154724 5024
rect 155408 4972 155460 5024
rect 157064 4972 157116 5024
rect 157248 4972 157300 5024
rect 20672 4870 20724 4922
rect 20736 4870 20788 4922
rect 20800 4870 20852 4922
rect 20864 4870 20916 4922
rect 20928 4870 20980 4922
rect 60117 4870 60169 4922
rect 60181 4870 60233 4922
rect 60245 4870 60297 4922
rect 60309 4870 60361 4922
rect 60373 4870 60425 4922
rect 99562 4870 99614 4922
rect 99626 4870 99678 4922
rect 99690 4870 99742 4922
rect 99754 4870 99806 4922
rect 99818 4870 99870 4922
rect 139007 4870 139059 4922
rect 139071 4870 139123 4922
rect 139135 4870 139187 4922
rect 139199 4870 139251 4922
rect 139263 4870 139315 4922
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 6000 4768 6052 4820
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 12624 4768 12676 4820
rect 13268 4768 13320 4820
rect 14372 4768 14424 4820
rect 14924 4768 14976 4820
rect 15108 4768 15160 4820
rect 5172 4700 5224 4752
rect 14464 4700 14516 4752
rect 18236 4768 18288 4820
rect 19708 4768 19760 4820
rect 24676 4811 24728 4820
rect 24676 4777 24685 4811
rect 24685 4777 24719 4811
rect 24719 4777 24728 4811
rect 24676 4768 24728 4777
rect 25228 4811 25280 4820
rect 25228 4777 25237 4811
rect 25237 4777 25271 4811
rect 25271 4777 25280 4811
rect 25228 4768 25280 4777
rect 27068 4768 27120 4820
rect 27804 4768 27856 4820
rect 30748 4811 30800 4820
rect 13636 4632 13688 4684
rect 19432 4700 19484 4752
rect 14832 4632 14884 4684
rect 5356 4564 5408 4616
rect 12164 4607 12216 4616
rect 12164 4573 12173 4607
rect 12173 4573 12207 4607
rect 12207 4573 12216 4607
rect 12164 4564 12216 4573
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 13820 4564 13872 4616
rect 12624 4496 12676 4548
rect 17040 4607 17092 4616
rect 17040 4573 17058 4607
rect 17058 4573 17092 4607
rect 17040 4564 17092 4573
rect 17868 4564 17920 4616
rect 17960 4564 18012 4616
rect 22468 4700 22520 4752
rect 30380 4700 30432 4752
rect 30748 4777 30757 4811
rect 30757 4777 30791 4811
rect 30791 4777 30800 4811
rect 30748 4768 30800 4777
rect 45192 4768 45244 4820
rect 46112 4811 46164 4820
rect 46112 4777 46121 4811
rect 46121 4777 46155 4811
rect 46155 4777 46164 4811
rect 46112 4768 46164 4777
rect 49240 4768 49292 4820
rect 73160 4768 73212 4820
rect 73344 4811 73396 4820
rect 73344 4777 73353 4811
rect 73353 4777 73387 4811
rect 73387 4777 73396 4811
rect 73344 4768 73396 4777
rect 81072 4768 81124 4820
rect 87972 4768 88024 4820
rect 88340 4811 88392 4820
rect 88340 4777 88349 4811
rect 88349 4777 88383 4811
rect 88383 4777 88392 4811
rect 88340 4768 88392 4777
rect 93676 4768 93728 4820
rect 95332 4768 95384 4820
rect 44180 4743 44232 4752
rect 44180 4709 44189 4743
rect 44189 4709 44223 4743
rect 44223 4709 44232 4743
rect 44180 4700 44232 4709
rect 50436 4743 50488 4752
rect 50436 4709 50445 4743
rect 50445 4709 50479 4743
rect 50479 4709 50488 4743
rect 50436 4700 50488 4709
rect 22652 4632 22704 4684
rect 23848 4632 23900 4684
rect 25228 4632 25280 4684
rect 30564 4632 30616 4684
rect 31024 4632 31076 4684
rect 21180 4564 21232 4616
rect 25320 4564 25372 4616
rect 30104 4607 30156 4616
rect 21640 4539 21692 4548
rect 13820 4428 13872 4480
rect 15016 4428 15068 4480
rect 17868 4471 17920 4480
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 21640 4505 21674 4539
rect 21674 4505 21692 4539
rect 21640 4496 21692 4505
rect 25780 4496 25832 4548
rect 30104 4573 30113 4607
rect 30113 4573 30147 4607
rect 30147 4573 30156 4607
rect 30104 4564 30156 4573
rect 38568 4564 38620 4616
rect 43996 4496 44048 4548
rect 45468 4564 45520 4616
rect 81900 4632 81952 4684
rect 98184 4768 98236 4820
rect 104624 4768 104676 4820
rect 108120 4768 108172 4820
rect 109500 4768 109552 4820
rect 117228 4768 117280 4820
rect 117780 4811 117832 4820
rect 117780 4777 117789 4811
rect 117789 4777 117823 4811
rect 117823 4777 117832 4811
rect 117780 4768 117832 4777
rect 115112 4700 115164 4752
rect 117872 4700 117924 4752
rect 118148 4700 118200 4752
rect 119068 4768 119120 4820
rect 121828 4768 121880 4820
rect 122472 4768 122524 4820
rect 125324 4700 125376 4752
rect 125416 4700 125468 4752
rect 125968 4700 126020 4752
rect 127992 4700 128044 4752
rect 131488 4700 131540 4752
rect 96620 4632 96672 4684
rect 52276 4564 52328 4616
rect 73528 4564 73580 4616
rect 84292 4607 84344 4616
rect 47216 4496 47268 4548
rect 76380 4539 76432 4548
rect 76380 4505 76389 4539
rect 76389 4505 76423 4539
rect 76423 4505 76432 4539
rect 76380 4496 76432 4505
rect 84292 4573 84301 4607
rect 84301 4573 84335 4607
rect 84335 4573 84344 4607
rect 84292 4564 84344 4573
rect 88892 4564 88944 4616
rect 92572 4564 92624 4616
rect 21824 4428 21876 4480
rect 21916 4428 21968 4480
rect 24768 4428 24820 4480
rect 26240 4428 26292 4480
rect 91928 4496 91980 4548
rect 98552 4539 98604 4548
rect 98552 4505 98561 4539
rect 98561 4505 98595 4539
rect 98595 4505 98604 4539
rect 98552 4496 98604 4505
rect 101680 4564 101732 4616
rect 105268 4564 105320 4616
rect 108488 4564 108540 4616
rect 113732 4632 113784 4684
rect 116124 4632 116176 4684
rect 116768 4632 116820 4684
rect 119252 4632 119304 4684
rect 122748 4632 122800 4684
rect 109776 4564 109828 4616
rect 114100 4564 114152 4616
rect 109224 4496 109276 4548
rect 114652 4539 114704 4548
rect 114652 4505 114670 4539
rect 114670 4505 114704 4539
rect 114652 4496 114704 4505
rect 115388 4496 115440 4548
rect 117688 4496 117740 4548
rect 118056 4496 118108 4548
rect 122840 4564 122892 4616
rect 124128 4632 124180 4684
rect 126980 4675 127032 4684
rect 126980 4641 126989 4675
rect 126989 4641 127023 4675
rect 127023 4641 127032 4675
rect 126980 4632 127032 4641
rect 129372 4632 129424 4684
rect 131764 4700 131816 4752
rect 134616 4768 134668 4820
rect 135076 4811 135128 4820
rect 135076 4777 135085 4811
rect 135085 4777 135119 4811
rect 135119 4777 135128 4811
rect 135076 4768 135128 4777
rect 135904 4768 135956 4820
rect 138572 4768 138624 4820
rect 143816 4768 143868 4820
rect 146024 4768 146076 4820
rect 132316 4632 132368 4684
rect 138296 4700 138348 4752
rect 139032 4743 139084 4752
rect 139032 4709 139041 4743
rect 139041 4709 139075 4743
rect 139075 4709 139084 4743
rect 139032 4700 139084 4709
rect 140780 4700 140832 4752
rect 145288 4700 145340 4752
rect 145564 4700 145616 4752
rect 145840 4700 145892 4752
rect 151268 4768 151320 4820
rect 151452 4768 151504 4820
rect 152832 4811 152884 4820
rect 152832 4777 152841 4811
rect 152841 4777 152875 4811
rect 152875 4777 152884 4811
rect 152832 4768 152884 4777
rect 152924 4768 152976 4820
rect 159272 4768 159324 4820
rect 150072 4743 150124 4752
rect 150072 4709 150081 4743
rect 150081 4709 150115 4743
rect 150115 4709 150124 4743
rect 150072 4700 150124 4709
rect 152188 4700 152240 4752
rect 152464 4700 152516 4752
rect 154304 4700 154356 4752
rect 123944 4564 123996 4616
rect 133052 4564 133104 4616
rect 133604 4564 133656 4616
rect 135720 4564 135772 4616
rect 142436 4675 142488 4684
rect 101772 4428 101824 4480
rect 112168 4428 112220 4480
rect 113548 4471 113600 4480
rect 113548 4437 113557 4471
rect 113557 4437 113591 4471
rect 113591 4437 113600 4471
rect 113548 4428 113600 4437
rect 115572 4428 115624 4480
rect 115848 4428 115900 4480
rect 118148 4428 118200 4480
rect 119252 4428 119304 4480
rect 120356 4428 120408 4480
rect 121184 4428 121236 4480
rect 125416 4496 125468 4548
rect 128912 4496 128964 4548
rect 129832 4496 129884 4548
rect 124128 4428 124180 4480
rect 124864 4471 124916 4480
rect 124864 4437 124873 4471
rect 124873 4437 124907 4471
rect 124907 4437 124916 4471
rect 124864 4428 124916 4437
rect 126520 4428 126572 4480
rect 127808 4428 127860 4480
rect 127992 4428 128044 4480
rect 131120 4471 131172 4480
rect 131120 4437 131129 4471
rect 131129 4437 131163 4471
rect 131163 4437 131172 4471
rect 131120 4428 131172 4437
rect 132500 4428 132552 4480
rect 138388 4564 138440 4616
rect 139952 4564 140004 4616
rect 140596 4607 140648 4616
rect 139032 4496 139084 4548
rect 140596 4573 140605 4607
rect 140605 4573 140639 4607
rect 140639 4573 140648 4607
rect 140596 4564 140648 4573
rect 142436 4641 142445 4675
rect 142445 4641 142479 4675
rect 142479 4641 142488 4675
rect 142436 4632 142488 4641
rect 147496 4675 147548 4684
rect 143080 4607 143132 4616
rect 143080 4573 143089 4607
rect 143089 4573 143123 4607
rect 143123 4573 143132 4607
rect 143080 4564 143132 4573
rect 147496 4641 147505 4675
rect 147505 4641 147539 4675
rect 147539 4641 147548 4675
rect 147496 4632 147548 4641
rect 157248 4700 157300 4752
rect 143356 4607 143408 4616
rect 143356 4573 143365 4607
rect 143365 4573 143399 4607
rect 143399 4573 143408 4607
rect 143356 4564 143408 4573
rect 144184 4564 144236 4616
rect 144276 4607 144328 4616
rect 144276 4573 144285 4607
rect 144285 4573 144319 4607
rect 144319 4573 144328 4607
rect 144276 4564 144328 4573
rect 145840 4564 145892 4616
rect 147680 4564 147732 4616
rect 159364 4632 159416 4684
rect 151820 4564 151872 4616
rect 152096 4607 152148 4616
rect 151084 4496 151136 4548
rect 141056 4471 141108 4480
rect 141056 4437 141065 4471
rect 141065 4437 141099 4471
rect 141099 4437 141108 4471
rect 141056 4428 141108 4437
rect 141424 4428 141476 4480
rect 145564 4428 145616 4480
rect 146760 4428 146812 4480
rect 146944 4428 146996 4480
rect 149428 4428 149480 4480
rect 149888 4428 149940 4480
rect 151636 4496 151688 4548
rect 152096 4573 152105 4607
rect 152105 4573 152139 4607
rect 152139 4573 152148 4607
rect 152096 4564 152148 4573
rect 153568 4607 153620 4616
rect 153568 4573 153577 4607
rect 153577 4573 153611 4607
rect 153611 4573 153620 4607
rect 153568 4564 153620 4573
rect 153660 4564 153712 4616
rect 154580 4607 154632 4616
rect 154580 4573 154589 4607
rect 154589 4573 154623 4607
rect 154623 4573 154632 4607
rect 154580 4564 154632 4573
rect 155132 4607 155184 4616
rect 155132 4573 155141 4607
rect 155141 4573 155175 4607
rect 155175 4573 155184 4607
rect 155132 4564 155184 4573
rect 155224 4564 155276 4616
rect 156144 4607 156196 4616
rect 156144 4573 156153 4607
rect 156153 4573 156187 4607
rect 156187 4573 156196 4607
rect 156144 4564 156196 4573
rect 156880 4564 156932 4616
rect 157984 4564 158036 4616
rect 154948 4496 155000 4548
rect 152280 4471 152332 4480
rect 152280 4437 152289 4471
rect 152289 4437 152323 4471
rect 152323 4437 152332 4471
rect 152280 4428 152332 4437
rect 155316 4428 155368 4480
rect 157248 4471 157300 4480
rect 157248 4437 157257 4471
rect 157257 4437 157291 4471
rect 157291 4437 157300 4471
rect 157248 4428 157300 4437
rect 40394 4326 40446 4378
rect 40458 4326 40510 4378
rect 40522 4326 40574 4378
rect 40586 4326 40638 4378
rect 40650 4326 40702 4378
rect 79839 4326 79891 4378
rect 79903 4326 79955 4378
rect 79967 4326 80019 4378
rect 80031 4326 80083 4378
rect 80095 4326 80147 4378
rect 119284 4326 119336 4378
rect 119348 4326 119400 4378
rect 119412 4326 119464 4378
rect 119476 4326 119528 4378
rect 119540 4326 119592 4378
rect 158729 4326 158781 4378
rect 158793 4326 158845 4378
rect 158857 4326 158909 4378
rect 158921 4326 158973 4378
rect 158985 4326 159037 4378
rect 10416 4224 10468 4276
rect 19524 4224 19576 4276
rect 20168 4224 20220 4276
rect 43076 4224 43128 4276
rect 56784 4224 56836 4276
rect 12624 4199 12676 4208
rect 12624 4165 12633 4199
rect 12633 4165 12667 4199
rect 12667 4165 12676 4199
rect 12624 4156 12676 4165
rect 14280 4156 14332 4208
rect 16764 4156 16816 4208
rect 18880 4156 18932 4208
rect 21180 4156 21232 4208
rect 23664 4156 23716 4208
rect 9128 4088 9180 4140
rect 9588 4088 9640 4140
rect 10968 4088 11020 4140
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 13912 4088 13964 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 17684 4131 17736 4140
rect 13728 4020 13780 4072
rect 6828 3952 6880 4004
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 17868 4088 17920 4140
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 18788 4131 18840 4140
rect 18788 4097 18822 4131
rect 18822 4097 18840 4131
rect 18788 4088 18840 4097
rect 20076 4088 20128 4140
rect 20444 4088 20496 4140
rect 24584 4088 24636 4140
rect 30564 4156 30616 4208
rect 42892 4088 42944 4140
rect 19524 4020 19576 4072
rect 30564 4020 30616 4072
rect 31852 4020 31904 4072
rect 37188 4020 37240 4072
rect 41972 4063 42024 4072
rect 41972 4029 41981 4063
rect 41981 4029 42015 4063
rect 42015 4029 42024 4063
rect 44180 4088 44232 4140
rect 44640 4088 44692 4140
rect 45284 4088 45336 4140
rect 47952 4131 48004 4140
rect 47952 4097 47961 4131
rect 47961 4097 47995 4131
rect 47995 4097 48004 4131
rect 47952 4088 48004 4097
rect 50988 4156 51040 4208
rect 41972 4020 42024 4029
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12624 3884 12676 3936
rect 13268 3884 13320 3936
rect 13544 3884 13596 3936
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 18420 3884 18472 3936
rect 30472 3952 30524 4004
rect 30840 3952 30892 4004
rect 34428 3952 34480 4004
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 21180 3884 21232 3893
rect 31116 3884 31168 3936
rect 31760 3884 31812 3936
rect 32864 3927 32916 3936
rect 32864 3893 32873 3927
rect 32873 3893 32907 3927
rect 32907 3893 32916 3927
rect 32864 3884 32916 3893
rect 49792 4020 49844 4072
rect 45468 3952 45520 4004
rect 47584 3884 47636 3936
rect 48964 3884 49016 3936
rect 54668 3884 54720 3936
rect 58532 4020 58584 4072
rect 62120 4088 62172 4140
rect 63316 4224 63368 4276
rect 98552 4224 98604 4276
rect 110328 4224 110380 4276
rect 113732 4224 113784 4276
rect 118792 4224 118844 4276
rect 125048 4267 125100 4276
rect 125048 4233 125057 4267
rect 125057 4233 125091 4267
rect 125091 4233 125100 4267
rect 125048 4224 125100 4233
rect 127532 4224 127584 4276
rect 76380 4088 76432 4140
rect 78956 4088 79008 4140
rect 105176 4156 105228 4208
rect 105268 4156 105320 4208
rect 106556 4088 106608 4140
rect 109316 4088 109368 4140
rect 111156 4088 111208 4140
rect 64880 4020 64932 4072
rect 76012 4020 76064 4072
rect 109040 4063 109092 4072
rect 109040 4029 109049 4063
rect 109049 4029 109083 4063
rect 109083 4029 109092 4063
rect 109040 4020 109092 4029
rect 110972 4063 111024 4072
rect 110972 4029 110981 4063
rect 110981 4029 111015 4063
rect 111015 4029 111024 4063
rect 110972 4020 111024 4029
rect 114192 4156 114244 4208
rect 114652 4088 114704 4140
rect 115572 4088 115624 4140
rect 115756 4088 115808 4140
rect 118240 4131 118292 4140
rect 55772 3952 55824 4004
rect 60464 3884 60516 3936
rect 66260 3884 66312 3936
rect 74816 3927 74868 3936
rect 74816 3893 74825 3927
rect 74825 3893 74859 3927
rect 74859 3893 74868 3927
rect 74816 3884 74868 3893
rect 93032 3952 93084 4004
rect 107660 3995 107712 4004
rect 84844 3884 84896 3936
rect 91560 3884 91612 3936
rect 102968 3884 103020 3936
rect 107660 3961 107669 3995
rect 107669 3961 107703 3995
rect 107703 3961 107712 3995
rect 107660 3952 107712 3961
rect 109684 3952 109736 4004
rect 106004 3927 106056 3936
rect 106004 3893 106013 3927
rect 106013 3893 106047 3927
rect 106047 3893 106056 3927
rect 106004 3884 106056 3893
rect 113732 4020 113784 4072
rect 116768 4020 116820 4072
rect 118240 4097 118249 4131
rect 118249 4097 118283 4131
rect 118283 4097 118292 4131
rect 118240 4088 118292 4097
rect 118424 4131 118476 4140
rect 118424 4097 118433 4131
rect 118433 4097 118467 4131
rect 118467 4097 118476 4131
rect 118424 4088 118476 4097
rect 118608 4131 118660 4140
rect 118608 4097 118617 4131
rect 118617 4097 118651 4131
rect 118651 4097 118660 4131
rect 118608 4088 118660 4097
rect 119160 4156 119212 4208
rect 128176 4156 128228 4208
rect 128268 4156 128320 4208
rect 122748 4088 122800 4140
rect 122840 4088 122892 4140
rect 123300 4088 123352 4140
rect 123944 4088 123996 4140
rect 125232 4131 125284 4140
rect 125232 4097 125241 4131
rect 125241 4097 125275 4131
rect 125275 4097 125284 4131
rect 125232 4088 125284 4097
rect 125324 4088 125376 4140
rect 126152 4088 126204 4140
rect 111616 3952 111668 4004
rect 117780 3884 117832 3936
rect 118976 3952 119028 4004
rect 121000 3952 121052 4004
rect 122748 3952 122800 4004
rect 119252 3884 119304 3936
rect 120080 3884 120132 3936
rect 121184 3884 121236 3936
rect 122012 3927 122064 3936
rect 122012 3893 122021 3927
rect 122021 3893 122055 3927
rect 122055 3893 122064 3927
rect 122012 3884 122064 3893
rect 125508 4020 125560 4072
rect 127992 4088 128044 4140
rect 131672 4156 131724 4208
rect 133236 4224 133288 4276
rect 140136 4224 140188 4276
rect 141148 4267 141200 4276
rect 141148 4233 141157 4267
rect 141157 4233 141191 4267
rect 141191 4233 141200 4267
rect 141148 4224 141200 4233
rect 137928 4156 137980 4208
rect 129924 4020 129976 4072
rect 126060 3952 126112 4004
rect 127440 3995 127492 4004
rect 127440 3961 127449 3995
rect 127449 3961 127483 3995
rect 127483 3961 127492 3995
rect 127440 3952 127492 3961
rect 127624 3884 127676 3936
rect 127992 3884 128044 3936
rect 129004 3884 129056 3936
rect 131764 4088 131816 4140
rect 132040 4020 132092 4072
rect 133604 4020 133656 4072
rect 133972 4020 134024 4072
rect 134248 4020 134300 4072
rect 134984 4020 135036 4072
rect 131764 3952 131816 4004
rect 135260 3884 135312 3936
rect 138296 4131 138348 4140
rect 138296 4097 138330 4131
rect 138330 4097 138348 4131
rect 138296 4088 138348 4097
rect 139860 4088 139912 4140
rect 140320 4088 140372 4140
rect 143356 4156 143408 4208
rect 157248 4224 157300 4276
rect 145564 4156 145616 4208
rect 146668 4156 146720 4208
rect 149244 4156 149296 4208
rect 142896 4131 142948 4140
rect 142896 4097 142914 4131
rect 142914 4097 142948 4131
rect 142896 4088 142948 4097
rect 135720 4020 135772 4072
rect 136088 4020 136140 4072
rect 137836 4020 137888 4072
rect 144184 4088 144236 4140
rect 145196 4088 145248 4140
rect 147220 4088 147272 4140
rect 148784 4088 148836 4140
rect 148048 4063 148100 4072
rect 137652 3952 137704 4004
rect 139400 3995 139452 4004
rect 139400 3961 139409 3995
rect 139409 3961 139443 3995
rect 139443 3961 139452 3995
rect 139400 3952 139452 3961
rect 139952 3995 140004 4004
rect 139952 3961 139961 3995
rect 139961 3961 139995 3995
rect 139995 3961 140004 3995
rect 139952 3952 140004 3961
rect 141056 3952 141108 4004
rect 141792 3995 141844 4004
rect 141792 3961 141801 3995
rect 141801 3961 141835 3995
rect 141835 3961 141844 3995
rect 141792 3952 141844 3961
rect 139768 3884 139820 3936
rect 140044 3884 140096 3936
rect 140504 3927 140556 3936
rect 140504 3893 140513 3927
rect 140513 3893 140547 3927
rect 140547 3893 140556 3927
rect 140504 3884 140556 3893
rect 141424 3884 141476 3936
rect 145564 3952 145616 4004
rect 143632 3927 143684 3936
rect 143632 3893 143641 3927
rect 143641 3893 143675 3927
rect 143675 3893 143684 3927
rect 146944 3952 146996 4004
rect 146668 3927 146720 3936
rect 143632 3884 143684 3893
rect 146668 3893 146677 3927
rect 146677 3893 146711 3927
rect 146711 3893 146720 3927
rect 146668 3884 146720 3893
rect 148048 4029 148057 4063
rect 148057 4029 148091 4063
rect 148091 4029 148100 4063
rect 148048 4020 148100 4029
rect 151820 4156 151872 4208
rect 149888 4131 149940 4140
rect 149888 4097 149897 4131
rect 149897 4097 149931 4131
rect 149931 4097 149940 4131
rect 149888 4088 149940 4097
rect 151544 4088 151596 4140
rect 152004 4131 152056 4140
rect 152004 4097 152022 4131
rect 152022 4097 152056 4131
rect 154672 4156 154724 4208
rect 152740 4131 152792 4140
rect 152004 4088 152056 4097
rect 150072 4020 150124 4072
rect 151268 4020 151320 4072
rect 152464 4020 152516 4072
rect 152740 4097 152749 4131
rect 152749 4097 152783 4131
rect 152783 4097 152792 4131
rect 152740 4088 152792 4097
rect 155224 4088 155276 4140
rect 154672 4063 154724 4072
rect 154672 4029 154681 4063
rect 154681 4029 154715 4063
rect 154715 4029 154724 4063
rect 154672 4020 154724 4029
rect 156420 4088 156472 4140
rect 156512 4088 156564 4140
rect 157708 4088 157760 4140
rect 158260 4131 158312 4140
rect 158260 4097 158269 4131
rect 158269 4097 158303 4131
rect 158303 4097 158312 4131
rect 158260 4088 158312 4097
rect 147680 3884 147732 3936
rect 147864 3884 147916 3936
rect 148508 3927 148560 3936
rect 148508 3893 148517 3927
rect 148517 3893 148551 3927
rect 148551 3893 148560 3927
rect 148508 3884 148560 3893
rect 150900 3927 150952 3936
rect 150900 3893 150909 3927
rect 150909 3893 150943 3927
rect 150943 3893 150952 3927
rect 150900 3884 150952 3893
rect 153292 3927 153344 3936
rect 153292 3893 153301 3927
rect 153301 3893 153335 3927
rect 153335 3893 153344 3927
rect 153292 3884 153344 3893
rect 155132 3995 155184 4004
rect 155132 3961 155141 3995
rect 155141 3961 155175 3995
rect 155175 3961 155184 3995
rect 155132 3952 155184 3961
rect 156052 3952 156104 4004
rect 154948 3884 155000 3936
rect 156420 3884 156472 3936
rect 156788 3927 156840 3936
rect 156788 3893 156797 3927
rect 156797 3893 156831 3927
rect 156831 3893 156840 3927
rect 156788 3884 156840 3893
rect 156880 3884 156932 3936
rect 20672 3782 20724 3834
rect 20736 3782 20788 3834
rect 20800 3782 20852 3834
rect 20864 3782 20916 3834
rect 20928 3782 20980 3834
rect 60117 3782 60169 3834
rect 60181 3782 60233 3834
rect 60245 3782 60297 3834
rect 60309 3782 60361 3834
rect 60373 3782 60425 3834
rect 99562 3782 99614 3834
rect 99626 3782 99678 3834
rect 99690 3782 99742 3834
rect 99754 3782 99806 3834
rect 99818 3782 99870 3834
rect 139007 3782 139059 3834
rect 139071 3782 139123 3834
rect 139135 3782 139187 3834
rect 139199 3782 139251 3834
rect 139263 3782 139315 3834
rect 14004 3680 14056 3732
rect 16120 3680 16172 3732
rect 20444 3680 20496 3732
rect 21824 3680 21876 3732
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 25228 3680 25280 3732
rect 25872 3680 25924 3732
rect 30564 3723 30616 3732
rect 30564 3689 30573 3723
rect 30573 3689 30607 3723
rect 30607 3689 30616 3723
rect 30564 3680 30616 3689
rect 16304 3612 16356 3664
rect 20720 3612 20772 3664
rect 21640 3612 21692 3664
rect 24768 3612 24820 3664
rect 36912 3680 36964 3732
rect 37188 3680 37240 3732
rect 45468 3680 45520 3732
rect 32588 3612 32640 3664
rect 37372 3612 37424 3664
rect 37740 3612 37792 3664
rect 45192 3655 45244 3664
rect 45192 3621 45201 3655
rect 45201 3621 45235 3655
rect 45235 3621 45244 3655
rect 45192 3612 45244 3621
rect 13268 3544 13320 3596
rect 31116 3587 31168 3596
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14004 3408 14056 3460
rect 16672 3476 16724 3528
rect 16304 3408 16356 3460
rect 13544 3340 13596 3392
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 17592 3408 17644 3460
rect 17960 3340 18012 3392
rect 18236 3476 18288 3528
rect 18512 3476 18564 3528
rect 20076 3476 20128 3528
rect 22560 3476 22612 3528
rect 18420 3408 18472 3460
rect 19892 3408 19944 3460
rect 25228 3476 25280 3528
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 31116 3553 31125 3587
rect 31125 3553 31159 3587
rect 31159 3553 31168 3587
rect 31116 3544 31168 3553
rect 50896 3680 50948 3732
rect 34336 3519 34388 3528
rect 34336 3485 34345 3519
rect 34345 3485 34379 3519
rect 34379 3485 34388 3519
rect 34336 3476 34388 3485
rect 37188 3519 37240 3528
rect 37188 3485 37197 3519
rect 37197 3485 37231 3519
rect 37231 3485 37240 3519
rect 37372 3519 37424 3528
rect 37188 3476 37240 3485
rect 37372 3485 37381 3519
rect 37381 3485 37415 3519
rect 37415 3485 37424 3519
rect 37372 3476 37424 3485
rect 46572 3519 46624 3528
rect 46572 3485 46581 3519
rect 46581 3485 46615 3519
rect 46615 3485 46624 3519
rect 46572 3476 46624 3485
rect 24400 3340 24452 3392
rect 30564 3340 30616 3392
rect 32864 3408 32916 3460
rect 33784 3340 33836 3392
rect 37924 3340 37976 3392
rect 49700 3408 49752 3460
rect 52368 3544 52420 3596
rect 57244 3544 57296 3596
rect 58532 3587 58584 3596
rect 58532 3553 58541 3587
rect 58541 3553 58575 3587
rect 58575 3553 58584 3587
rect 58532 3544 58584 3553
rect 58716 3544 58768 3596
rect 62120 3680 62172 3732
rect 63500 3680 63552 3732
rect 64604 3680 64656 3732
rect 64880 3723 64932 3732
rect 64880 3689 64889 3723
rect 64889 3689 64923 3723
rect 64923 3689 64932 3723
rect 64880 3680 64932 3689
rect 73160 3723 73212 3732
rect 73160 3689 73169 3723
rect 73169 3689 73203 3723
rect 73203 3689 73212 3723
rect 73160 3680 73212 3689
rect 77116 3680 77168 3732
rect 88432 3723 88484 3732
rect 59176 3612 59228 3664
rect 53748 3519 53800 3528
rect 53748 3485 53757 3519
rect 53757 3485 53791 3519
rect 53791 3485 53800 3519
rect 53748 3476 53800 3485
rect 58440 3476 58492 3528
rect 62028 3451 62080 3460
rect 46848 3340 46900 3392
rect 49608 3340 49660 3392
rect 62028 3417 62037 3451
rect 62037 3417 62071 3451
rect 62071 3417 62080 3451
rect 62028 3408 62080 3417
rect 65800 3476 65852 3528
rect 88432 3689 88441 3723
rect 88441 3689 88475 3723
rect 88475 3689 88484 3723
rect 94504 3723 94556 3732
rect 88432 3680 88484 3689
rect 80244 3612 80296 3664
rect 94504 3689 94513 3723
rect 94513 3689 94547 3723
rect 94547 3689 94556 3723
rect 94504 3680 94556 3689
rect 99012 3612 99064 3664
rect 102048 3680 102100 3732
rect 108212 3680 108264 3732
rect 113916 3680 113968 3732
rect 117964 3680 118016 3732
rect 74540 3519 74592 3528
rect 74540 3485 74549 3519
rect 74549 3485 74583 3519
rect 74583 3485 74592 3519
rect 74540 3476 74592 3485
rect 90548 3476 90600 3528
rect 105176 3544 105228 3596
rect 96252 3476 96304 3528
rect 109040 3476 109092 3528
rect 109592 3476 109644 3528
rect 110972 3544 111024 3596
rect 116768 3587 116820 3596
rect 116768 3553 116777 3587
rect 116777 3553 116811 3587
rect 116811 3553 116820 3587
rect 116768 3544 116820 3553
rect 126152 3680 126204 3732
rect 126888 3680 126940 3732
rect 127900 3680 127952 3732
rect 127992 3680 128044 3732
rect 138756 3680 138808 3732
rect 123024 3612 123076 3664
rect 121000 3587 121052 3596
rect 110052 3476 110104 3528
rect 117780 3519 117832 3528
rect 67548 3408 67600 3460
rect 74448 3408 74500 3460
rect 84844 3408 84896 3460
rect 51080 3340 51132 3392
rect 53564 3383 53616 3392
rect 53564 3349 53573 3383
rect 53573 3349 53607 3383
rect 53607 3349 53616 3383
rect 53564 3340 53616 3349
rect 57152 3383 57204 3392
rect 57152 3349 57161 3383
rect 57161 3349 57195 3383
rect 57195 3349 57204 3383
rect 57152 3340 57204 3349
rect 57612 3340 57664 3392
rect 66168 3340 66220 3392
rect 69204 3340 69256 3392
rect 76104 3383 76156 3392
rect 76104 3349 76113 3383
rect 76113 3349 76147 3383
rect 76147 3349 76156 3383
rect 76104 3340 76156 3349
rect 102968 3451 103020 3460
rect 102968 3417 102986 3451
rect 102986 3417 103020 3451
rect 102968 3408 103020 3417
rect 110144 3408 110196 3460
rect 116952 3408 117004 3460
rect 117780 3485 117789 3519
rect 117789 3485 117823 3519
rect 117823 3485 117832 3519
rect 117780 3476 117832 3485
rect 118792 3476 118844 3528
rect 117688 3408 117740 3460
rect 121000 3553 121009 3587
rect 121009 3553 121043 3587
rect 121043 3553 121052 3587
rect 121000 3544 121052 3553
rect 122932 3544 122984 3596
rect 123300 3544 123352 3596
rect 123484 3544 123536 3596
rect 123944 3544 123996 3596
rect 125600 3612 125652 3664
rect 129464 3655 129516 3664
rect 119896 3476 119948 3528
rect 106464 3340 106516 3392
rect 108304 3383 108356 3392
rect 108304 3349 108313 3383
rect 108313 3349 108347 3383
rect 108347 3349 108356 3383
rect 108304 3340 108356 3349
rect 110052 3340 110104 3392
rect 111616 3340 111668 3392
rect 114836 3340 114888 3392
rect 118240 3340 118292 3392
rect 121276 3408 121328 3460
rect 119712 3340 119764 3392
rect 122564 3340 122616 3392
rect 123024 3383 123076 3392
rect 123024 3349 123033 3383
rect 123033 3349 123067 3383
rect 123067 3349 123076 3383
rect 123024 3340 123076 3349
rect 125324 3476 125376 3528
rect 125968 3519 126020 3528
rect 125968 3485 125977 3519
rect 125977 3485 126011 3519
rect 126011 3485 126020 3519
rect 125968 3476 126020 3485
rect 127716 3544 127768 3596
rect 127072 3519 127124 3528
rect 127072 3485 127081 3519
rect 127081 3485 127115 3519
rect 127115 3485 127124 3519
rect 127072 3476 127124 3485
rect 129464 3621 129473 3655
rect 129473 3621 129507 3655
rect 129507 3621 129516 3655
rect 129464 3612 129516 3621
rect 131028 3612 131080 3664
rect 137928 3612 137980 3664
rect 138020 3612 138072 3664
rect 128360 3476 128412 3528
rect 129740 3544 129792 3596
rect 131212 3544 131264 3596
rect 140504 3680 140556 3732
rect 142344 3680 142396 3732
rect 142620 3680 142672 3732
rect 146300 3723 146352 3732
rect 144184 3587 144236 3596
rect 144184 3553 144193 3587
rect 144193 3553 144227 3587
rect 144227 3553 144236 3587
rect 144184 3544 144236 3553
rect 129188 3476 129240 3528
rect 132500 3476 132552 3528
rect 132684 3476 132736 3528
rect 132960 3519 133012 3528
rect 132960 3485 132969 3519
rect 132969 3485 133003 3519
rect 133003 3485 133012 3519
rect 132960 3476 133012 3485
rect 133236 3476 133288 3528
rect 133512 3476 133564 3528
rect 135352 3519 135404 3528
rect 135352 3485 135361 3519
rect 135361 3485 135395 3519
rect 135395 3485 135404 3519
rect 135352 3476 135404 3485
rect 137284 3476 137336 3528
rect 137652 3476 137704 3528
rect 139952 3476 140004 3528
rect 143632 3476 143684 3528
rect 143724 3476 143776 3528
rect 146300 3689 146309 3723
rect 146309 3689 146343 3723
rect 146343 3689 146352 3723
rect 146300 3680 146352 3689
rect 145380 3612 145432 3664
rect 149520 3680 149572 3732
rect 149612 3680 149664 3732
rect 150164 3680 150216 3732
rect 152832 3723 152884 3732
rect 148324 3612 148376 3664
rect 152832 3689 152841 3723
rect 152841 3689 152875 3723
rect 152875 3689 152884 3723
rect 152832 3680 152884 3689
rect 156880 3680 156932 3732
rect 155684 3612 155736 3664
rect 151820 3587 151872 3596
rect 151820 3553 151829 3587
rect 151829 3553 151863 3587
rect 151863 3553 151872 3587
rect 151820 3544 151872 3553
rect 152556 3544 152608 3596
rect 129096 3408 129148 3460
rect 129740 3408 129792 3460
rect 130476 3408 130528 3460
rect 131212 3408 131264 3460
rect 127624 3340 127676 3392
rect 127716 3340 127768 3392
rect 129464 3340 129516 3392
rect 129924 3340 129976 3392
rect 138296 3408 138348 3460
rect 138756 3408 138808 3460
rect 139492 3408 139544 3460
rect 140688 3408 140740 3460
rect 141056 3408 141108 3460
rect 147680 3519 147732 3528
rect 147680 3485 147689 3519
rect 147689 3485 147723 3519
rect 147723 3485 147732 3519
rect 147680 3476 147732 3485
rect 148048 3476 148100 3528
rect 134708 3383 134760 3392
rect 134708 3349 134717 3383
rect 134717 3349 134751 3383
rect 134751 3349 134760 3383
rect 134708 3340 134760 3349
rect 135352 3340 135404 3392
rect 136456 3383 136508 3392
rect 136456 3349 136465 3383
rect 136465 3349 136499 3383
rect 136499 3349 136508 3383
rect 136456 3340 136508 3349
rect 136916 3383 136968 3392
rect 136916 3349 136925 3383
rect 136925 3349 136959 3383
rect 136959 3349 136968 3383
rect 136916 3340 136968 3349
rect 137192 3340 137244 3392
rect 139860 3340 139912 3392
rect 140596 3340 140648 3392
rect 142988 3340 143040 3392
rect 143724 3383 143776 3392
rect 143724 3349 143733 3383
rect 143733 3349 143767 3383
rect 143767 3349 143776 3383
rect 143724 3340 143776 3349
rect 145012 3408 145064 3460
rect 147312 3408 147364 3460
rect 147588 3408 147640 3460
rect 148232 3408 148284 3460
rect 149060 3476 149112 3528
rect 152464 3519 152516 3528
rect 149888 3408 149940 3460
rect 149980 3408 150032 3460
rect 150624 3408 150676 3460
rect 151544 3451 151596 3460
rect 151544 3417 151562 3451
rect 151562 3417 151596 3451
rect 151544 3408 151596 3417
rect 152464 3485 152473 3519
rect 152473 3485 152507 3519
rect 152507 3485 152516 3519
rect 152464 3476 152516 3485
rect 153108 3476 153160 3528
rect 154304 3476 154356 3528
rect 155132 3519 155184 3528
rect 155132 3485 155141 3519
rect 155141 3485 155175 3519
rect 155175 3485 155184 3519
rect 155132 3476 155184 3485
rect 155776 3519 155828 3528
rect 155776 3485 155785 3519
rect 155785 3485 155819 3519
rect 155819 3485 155828 3519
rect 155776 3476 155828 3485
rect 156972 3519 157024 3528
rect 154672 3408 154724 3460
rect 155040 3408 155092 3460
rect 155224 3408 155276 3460
rect 156972 3485 156981 3519
rect 156981 3485 157015 3519
rect 157015 3485 157024 3519
rect 156972 3476 157024 3485
rect 157616 3519 157668 3528
rect 157616 3485 157625 3519
rect 157625 3485 157659 3519
rect 157659 3485 157668 3519
rect 157616 3476 157668 3485
rect 146208 3340 146260 3392
rect 146576 3340 146628 3392
rect 149152 3340 149204 3392
rect 149244 3340 149296 3392
rect 151268 3340 151320 3392
rect 153384 3340 153436 3392
rect 153752 3383 153804 3392
rect 153752 3349 153761 3383
rect 153761 3349 153795 3383
rect 153795 3349 153804 3383
rect 153752 3340 153804 3349
rect 153936 3340 153988 3392
rect 157432 3383 157484 3392
rect 157432 3349 157441 3383
rect 157441 3349 157475 3383
rect 157475 3349 157484 3383
rect 157432 3340 157484 3349
rect 40394 3238 40446 3290
rect 40458 3238 40510 3290
rect 40522 3238 40574 3290
rect 40586 3238 40638 3290
rect 40650 3238 40702 3290
rect 79839 3238 79891 3290
rect 79903 3238 79955 3290
rect 79967 3238 80019 3290
rect 80031 3238 80083 3290
rect 80095 3238 80147 3290
rect 119284 3238 119336 3290
rect 119348 3238 119400 3290
rect 119412 3238 119464 3290
rect 119476 3238 119528 3290
rect 119540 3238 119592 3290
rect 158729 3238 158781 3290
rect 158793 3238 158845 3290
rect 158857 3238 158909 3290
rect 158921 3238 158973 3290
rect 158985 3238 159037 3290
rect 11060 3179 11112 3188
rect 11060 3145 11069 3179
rect 11069 3145 11103 3179
rect 11103 3145 11112 3179
rect 11060 3136 11112 3145
rect 11428 3136 11480 3188
rect 13912 3136 13964 3188
rect 14004 3136 14056 3188
rect 18788 3136 18840 3188
rect 20076 3179 20128 3188
rect 20076 3145 20085 3179
rect 20085 3145 20119 3179
rect 20119 3145 20128 3179
rect 20076 3136 20128 3145
rect 23940 3179 23992 3188
rect 13360 3068 13412 3120
rect 15108 3068 15160 3120
rect 18328 3068 18380 3120
rect 18604 3068 18656 3120
rect 20536 3068 20588 3120
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 13820 2932 13872 2984
rect 14464 2932 14516 2984
rect 19340 3000 19392 3052
rect 22468 3068 22520 3120
rect 23940 3145 23949 3179
rect 23949 3145 23983 3179
rect 23983 3145 23992 3179
rect 23940 3136 23992 3145
rect 24400 3136 24452 3188
rect 24676 3136 24728 3188
rect 24768 3136 24820 3188
rect 32772 3136 32824 3188
rect 32956 3136 33008 3188
rect 26792 3068 26844 3120
rect 26976 3068 27028 3120
rect 37924 3068 37976 3120
rect 50804 3136 50856 3188
rect 66260 3179 66312 3188
rect 47216 3111 47268 3120
rect 47216 3077 47225 3111
rect 47225 3077 47259 3111
rect 47259 3077 47268 3111
rect 47216 3068 47268 3077
rect 20812 3000 20864 3052
rect 22560 3043 22612 3052
rect 22560 3009 22569 3043
rect 22569 3009 22603 3043
rect 22603 3009 22612 3043
rect 22560 3000 22612 3009
rect 15200 2864 15252 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 17960 2796 18012 2848
rect 23940 2932 23992 2984
rect 31024 3000 31076 3052
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 33048 3000 33100 3052
rect 20720 2864 20772 2916
rect 22468 2864 22520 2916
rect 44180 3000 44232 3052
rect 46572 3000 46624 3052
rect 56416 3111 56468 3120
rect 48044 3043 48096 3052
rect 48044 3009 48078 3043
rect 48078 3009 48096 3043
rect 48044 3000 48096 3009
rect 49792 3000 49844 3052
rect 51080 3000 51132 3052
rect 56416 3077 56450 3111
rect 56450 3077 56468 3111
rect 56416 3068 56468 3077
rect 66260 3145 66269 3179
rect 66269 3145 66303 3179
rect 66303 3145 66312 3179
rect 66260 3136 66312 3145
rect 69112 3136 69164 3188
rect 69204 3136 69256 3188
rect 76104 3136 76156 3188
rect 81164 3136 81216 3188
rect 81348 3136 81400 3188
rect 83096 3136 83148 3188
rect 96252 3179 96304 3188
rect 96252 3145 96261 3179
rect 96261 3145 96295 3179
rect 96295 3145 96304 3179
rect 96252 3136 96304 3145
rect 109316 3136 109368 3188
rect 110144 3179 110196 3188
rect 110144 3145 110153 3179
rect 110153 3145 110187 3179
rect 110187 3145 110196 3179
rect 110144 3136 110196 3145
rect 114836 3179 114888 3188
rect 114836 3145 114845 3179
rect 114845 3145 114879 3179
rect 114879 3145 114888 3179
rect 114836 3136 114888 3145
rect 115664 3179 115716 3188
rect 115664 3145 115673 3179
rect 115673 3145 115707 3179
rect 115707 3145 115716 3179
rect 115664 3136 115716 3145
rect 116952 3179 117004 3188
rect 116952 3145 116961 3179
rect 116961 3145 116995 3179
rect 116995 3145 117004 3179
rect 116952 3136 117004 3145
rect 62028 3000 62080 3052
rect 64604 3043 64656 3052
rect 64604 3009 64613 3043
rect 64613 3009 64647 3043
rect 64647 3009 64656 3043
rect 64604 3000 64656 3009
rect 42892 2932 42944 2984
rect 19340 2796 19392 2848
rect 38844 2796 38896 2848
rect 40316 2796 40368 2848
rect 49700 2864 49752 2916
rect 57244 2864 57296 2916
rect 51724 2796 51776 2848
rect 57612 2796 57664 2848
rect 67548 3000 67600 3052
rect 108304 3068 108356 3120
rect 108396 3068 108448 3120
rect 118516 3068 118568 3120
rect 119160 3136 119212 3188
rect 126612 3136 126664 3188
rect 126796 3179 126848 3188
rect 126796 3145 126805 3179
rect 126805 3145 126839 3179
rect 126839 3145 126848 3179
rect 126796 3136 126848 3145
rect 127072 3136 127124 3188
rect 127900 3179 127952 3188
rect 127900 3145 127909 3179
rect 127909 3145 127943 3179
rect 127943 3145 127952 3179
rect 127900 3136 127952 3145
rect 129096 3179 129148 3188
rect 129096 3145 129105 3179
rect 129105 3145 129139 3179
rect 129139 3145 129148 3179
rect 129096 3136 129148 3145
rect 131948 3136 132000 3188
rect 132500 3136 132552 3188
rect 134708 3179 134760 3188
rect 134708 3145 134717 3179
rect 134717 3145 134751 3179
rect 134751 3145 134760 3179
rect 134708 3136 134760 3145
rect 135444 3179 135496 3188
rect 135444 3145 135453 3179
rect 135453 3145 135487 3179
rect 135487 3145 135496 3179
rect 135444 3136 135496 3145
rect 121092 3111 121144 3120
rect 121092 3077 121101 3111
rect 121101 3077 121135 3111
rect 121135 3077 121144 3111
rect 121092 3068 121144 3077
rect 122012 3068 122064 3120
rect 125968 3068 126020 3120
rect 69112 2932 69164 2984
rect 74540 2932 74592 2984
rect 96988 3000 97040 3052
rect 107660 3000 107712 3052
rect 88524 2932 88576 2984
rect 100852 2864 100904 2916
rect 106464 2932 106516 2984
rect 110052 2864 110104 2916
rect 83004 2839 83056 2848
rect 83004 2805 83013 2839
rect 83013 2805 83047 2839
rect 83047 2805 83056 2839
rect 83004 2796 83056 2805
rect 98644 2796 98696 2848
rect 114836 3000 114888 3052
rect 115480 3043 115532 3052
rect 115480 3009 115489 3043
rect 115489 3009 115523 3043
rect 115523 3009 115532 3043
rect 115480 3000 115532 3009
rect 118424 3000 118476 3052
rect 120080 2975 120132 2984
rect 120080 2941 120089 2975
rect 120089 2941 120123 2975
rect 120123 2941 120132 2975
rect 120080 2932 120132 2941
rect 120632 2975 120684 2984
rect 120632 2941 120641 2975
rect 120641 2941 120675 2975
rect 120675 2941 120684 2975
rect 120632 2932 120684 2941
rect 120908 2932 120960 2984
rect 122196 2975 122248 2984
rect 122196 2941 122205 2975
rect 122205 2941 122239 2975
rect 122239 2941 122248 2975
rect 122196 2932 122248 2941
rect 125600 2932 125652 2984
rect 125968 2932 126020 2984
rect 131580 3111 131632 3120
rect 131580 3077 131589 3111
rect 131589 3077 131623 3111
rect 131623 3077 131632 3111
rect 131580 3068 131632 3077
rect 131856 3068 131908 3120
rect 136364 3136 136416 3188
rect 136456 3136 136508 3188
rect 137560 3111 137612 3120
rect 137560 3077 137594 3111
rect 137594 3077 137612 3111
rect 137560 3068 137612 3077
rect 139676 3136 139728 3188
rect 139860 3179 139912 3188
rect 139860 3145 139869 3179
rect 139869 3145 139903 3179
rect 139903 3145 139912 3179
rect 139860 3136 139912 3145
rect 139952 3136 140004 3188
rect 141424 3179 141476 3188
rect 141424 3145 141433 3179
rect 141433 3145 141467 3179
rect 141467 3145 141476 3179
rect 141424 3136 141476 3145
rect 141976 3136 142028 3188
rect 141700 3068 141752 3120
rect 142620 3136 142672 3188
rect 142896 3136 142948 3188
rect 146484 3136 146536 3188
rect 147036 3179 147088 3188
rect 147036 3145 147045 3179
rect 147045 3145 147079 3179
rect 147079 3145 147088 3179
rect 147036 3136 147088 3145
rect 127532 3000 127584 3052
rect 126612 2932 126664 2984
rect 129372 3000 129424 3052
rect 130200 3000 130252 3052
rect 136916 3000 136968 3052
rect 137284 3043 137336 3052
rect 137284 3009 137293 3043
rect 137293 3009 137327 3043
rect 137327 3009 137336 3043
rect 137284 3000 137336 3009
rect 127808 2932 127860 2984
rect 110328 2864 110380 2916
rect 129924 2864 129976 2916
rect 111524 2796 111576 2848
rect 117596 2839 117648 2848
rect 117596 2805 117605 2839
rect 117605 2805 117639 2839
rect 117639 2805 117648 2839
rect 117596 2796 117648 2805
rect 117688 2796 117740 2848
rect 119160 2796 119212 2848
rect 119344 2839 119396 2848
rect 119344 2805 119353 2839
rect 119353 2805 119387 2839
rect 119387 2805 119396 2839
rect 119344 2796 119396 2805
rect 123392 2839 123444 2848
rect 123392 2805 123401 2839
rect 123401 2805 123435 2839
rect 123435 2805 123444 2839
rect 123392 2796 123444 2805
rect 123852 2839 123904 2848
rect 123852 2805 123861 2839
rect 123861 2805 123895 2839
rect 123895 2805 123904 2839
rect 123852 2796 123904 2805
rect 123944 2796 123996 2848
rect 125232 2796 125284 2848
rect 125876 2796 125928 2848
rect 126060 2796 126112 2848
rect 127900 2796 127952 2848
rect 128820 2796 128872 2848
rect 130200 2907 130252 2916
rect 130200 2873 130209 2907
rect 130209 2873 130243 2907
rect 130243 2873 130252 2907
rect 130200 2864 130252 2873
rect 142988 3068 143040 3120
rect 145472 3068 145524 3120
rect 147680 3136 147732 3188
rect 131120 2796 131172 2848
rect 133144 2796 133196 2848
rect 143816 2932 143868 2984
rect 136916 2796 136968 2848
rect 140688 2796 140740 2848
rect 145564 3000 145616 3052
rect 147588 3068 147640 3120
rect 150164 3136 150216 3188
rect 150716 3136 150768 3188
rect 147864 3068 147916 3120
rect 145288 2932 145340 2984
rect 145656 2975 145708 2984
rect 145656 2941 145665 2975
rect 145665 2941 145699 2975
rect 145699 2941 145708 2975
rect 145656 2932 145708 2941
rect 146944 2796 146996 2848
rect 149428 3000 149480 3052
rect 149520 3043 149572 3052
rect 149520 3009 149529 3043
rect 149529 3009 149563 3043
rect 149563 3009 149572 3043
rect 149520 3000 149572 3009
rect 150532 3000 150584 3052
rect 150624 3000 150676 3052
rect 149152 2932 149204 2984
rect 151452 3068 151504 3120
rect 152004 3111 152056 3120
rect 152004 3077 152013 3111
rect 152013 3077 152047 3111
rect 152047 3077 152056 3111
rect 152004 3068 152056 3077
rect 152280 3068 152332 3120
rect 151360 3000 151412 3052
rect 151820 2932 151872 2984
rect 151912 2932 151964 2984
rect 153016 2932 153068 2984
rect 153844 3000 153896 3052
rect 154396 3136 154448 3188
rect 154580 3179 154632 3188
rect 154580 3145 154589 3179
rect 154589 3145 154623 3179
rect 154623 3145 154632 3179
rect 154580 3136 154632 3145
rect 156604 3136 156656 3188
rect 158168 3136 158220 3188
rect 154488 3000 154540 3052
rect 155132 3000 155184 3052
rect 155408 3000 155460 3052
rect 157064 3043 157116 3052
rect 157064 3009 157073 3043
rect 157073 3009 157107 3043
rect 157107 3009 157116 3043
rect 157064 3000 157116 3009
rect 148600 2864 148652 2916
rect 148692 2796 148744 2848
rect 151268 2864 151320 2916
rect 153200 2864 153252 2916
rect 153476 2907 153528 2916
rect 153476 2873 153485 2907
rect 153485 2873 153519 2907
rect 153519 2873 153528 2907
rect 153476 2864 153528 2873
rect 154028 2932 154080 2984
rect 154948 2932 155000 2984
rect 156236 2932 156288 2984
rect 156328 2932 156380 2984
rect 155592 2864 155644 2916
rect 155960 2864 156012 2916
rect 154212 2796 154264 2848
rect 155776 2796 155828 2848
rect 156420 2839 156472 2848
rect 156420 2805 156429 2839
rect 156429 2805 156463 2839
rect 156463 2805 156472 2839
rect 156420 2796 156472 2805
rect 156512 2796 156564 2848
rect 157156 2796 157208 2848
rect 20672 2694 20724 2746
rect 20736 2694 20788 2746
rect 20800 2694 20852 2746
rect 20864 2694 20916 2746
rect 20928 2694 20980 2746
rect 60117 2694 60169 2746
rect 60181 2694 60233 2746
rect 60245 2694 60297 2746
rect 60309 2694 60361 2746
rect 60373 2694 60425 2746
rect 99562 2694 99614 2746
rect 99626 2694 99678 2746
rect 99690 2694 99742 2746
rect 99754 2694 99806 2746
rect 99818 2694 99870 2746
rect 139007 2694 139059 2746
rect 139071 2694 139123 2746
rect 139135 2694 139187 2746
rect 139199 2694 139251 2746
rect 139263 2694 139315 2746
rect 4712 2592 4764 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 13820 2592 13872 2644
rect 17960 2592 18012 2644
rect 18788 2592 18840 2644
rect 19616 2592 19668 2644
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 13636 2524 13688 2576
rect 19892 2524 19944 2576
rect 5816 2388 5868 2440
rect 11152 2456 11204 2508
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 24400 2456 24452 2508
rect 41328 2592 41380 2644
rect 49700 2592 49752 2644
rect 59820 2592 59872 2644
rect 63316 2592 63368 2644
rect 25964 2567 26016 2576
rect 25964 2533 25973 2567
rect 25973 2533 26007 2567
rect 26007 2533 26016 2567
rect 25964 2524 26016 2533
rect 33784 2499 33836 2508
rect 33784 2465 33793 2499
rect 33793 2465 33827 2499
rect 33827 2465 33836 2499
rect 33784 2456 33836 2465
rect 11060 2388 11112 2440
rect 17408 2388 17460 2440
rect 21088 2388 21140 2440
rect 23572 2388 23624 2440
rect 47308 2456 47360 2508
rect 58716 2499 58768 2508
rect 58716 2465 58725 2499
rect 58725 2465 58759 2499
rect 58759 2465 58768 2499
rect 58716 2456 58768 2465
rect 71044 2592 71096 2644
rect 81440 2635 81492 2644
rect 81440 2601 81449 2635
rect 81449 2601 81483 2635
rect 81483 2601 81492 2635
rect 81440 2592 81492 2601
rect 107292 2592 107344 2644
rect 109592 2635 109644 2644
rect 109592 2601 109601 2635
rect 109601 2601 109635 2635
rect 109635 2601 109644 2635
rect 109592 2592 109644 2601
rect 112720 2592 112772 2644
rect 113640 2635 113692 2644
rect 65984 2524 66036 2576
rect 11704 2320 11756 2372
rect 45376 2320 45428 2372
rect 56600 2388 56652 2440
rect 59268 2388 59320 2440
rect 74540 2388 74592 2440
rect 81348 2388 81400 2440
rect 111248 2388 111300 2440
rect 113640 2601 113649 2635
rect 113649 2601 113683 2635
rect 113683 2601 113692 2635
rect 113640 2592 113692 2601
rect 114468 2592 114520 2644
rect 123300 2592 123352 2644
rect 125140 2592 125192 2644
rect 126336 2592 126388 2644
rect 127072 2635 127124 2644
rect 127072 2601 127081 2635
rect 127081 2601 127115 2635
rect 127115 2601 127124 2635
rect 127072 2592 127124 2601
rect 130200 2635 130252 2644
rect 130200 2601 130209 2635
rect 130209 2601 130243 2635
rect 130243 2601 130252 2635
rect 130200 2592 130252 2601
rect 131580 2592 131632 2644
rect 134616 2635 134668 2644
rect 122196 2524 122248 2576
rect 126428 2567 126480 2576
rect 126428 2533 126437 2567
rect 126437 2533 126471 2567
rect 126471 2533 126480 2567
rect 126428 2524 126480 2533
rect 134616 2601 134625 2635
rect 134625 2601 134659 2635
rect 134659 2601 134668 2635
rect 134616 2592 134668 2601
rect 137284 2635 137336 2644
rect 137284 2601 137293 2635
rect 137293 2601 137327 2635
rect 137327 2601 137336 2635
rect 137284 2592 137336 2601
rect 138664 2592 138716 2644
rect 139768 2592 139820 2644
rect 141608 2592 141660 2644
rect 142528 2635 142580 2644
rect 142528 2601 142537 2635
rect 142537 2601 142571 2635
rect 142571 2601 142580 2635
rect 142528 2592 142580 2601
rect 144184 2592 144236 2644
rect 143724 2567 143776 2576
rect 143724 2533 143733 2567
rect 143733 2533 143767 2567
rect 143767 2533 143776 2567
rect 143724 2524 143776 2533
rect 129556 2499 129608 2508
rect 129556 2465 129565 2499
rect 129565 2465 129599 2499
rect 129599 2465 129608 2499
rect 129556 2456 129608 2465
rect 118792 2431 118844 2440
rect 118792 2397 118801 2431
rect 118801 2397 118835 2431
rect 118835 2397 118844 2431
rect 118792 2388 118844 2397
rect 120540 2388 120592 2440
rect 126336 2388 126388 2440
rect 131120 2456 131172 2508
rect 133144 2456 133196 2508
rect 135352 2499 135404 2508
rect 135352 2465 135361 2499
rect 135361 2465 135395 2499
rect 135395 2465 135404 2499
rect 135352 2456 135404 2465
rect 135628 2431 135680 2440
rect 135628 2397 135662 2431
rect 135662 2397 135680 2431
rect 75460 2320 75512 2372
rect 83004 2320 83056 2372
rect 119344 2320 119396 2372
rect 129004 2363 129056 2372
rect 129004 2329 129013 2363
rect 129013 2329 129047 2363
rect 129047 2329 129056 2363
rect 129004 2320 129056 2329
rect 135628 2388 135680 2397
rect 133144 2320 133196 2372
rect 138480 2456 138532 2508
rect 141976 2499 142028 2508
rect 141976 2465 141985 2499
rect 141985 2465 142019 2499
rect 142019 2465 142028 2499
rect 141976 2456 142028 2465
rect 148876 2592 148928 2644
rect 148968 2592 149020 2644
rect 152188 2635 152240 2644
rect 152188 2601 152197 2635
rect 152197 2601 152231 2635
rect 152231 2601 152240 2635
rect 152188 2592 152240 2601
rect 152740 2635 152792 2644
rect 152740 2601 152749 2635
rect 152749 2601 152783 2635
rect 152783 2601 152792 2635
rect 152740 2592 152792 2601
rect 159088 2592 159140 2644
rect 149428 2524 149480 2576
rect 150256 2524 150308 2576
rect 150440 2524 150492 2576
rect 145656 2499 145708 2508
rect 145656 2465 145665 2499
rect 145665 2465 145699 2499
rect 145699 2465 145708 2499
rect 145656 2456 145708 2465
rect 146944 2456 146996 2508
rect 138664 2431 138716 2440
rect 138664 2397 138673 2431
rect 138673 2397 138707 2431
rect 138707 2397 138716 2431
rect 138664 2388 138716 2397
rect 138020 2363 138072 2372
rect 138020 2329 138029 2363
rect 138029 2329 138063 2363
rect 138063 2329 138072 2363
rect 141884 2388 141936 2440
rect 138020 2320 138072 2329
rect 31760 2295 31812 2304
rect 31760 2261 31769 2295
rect 31769 2261 31803 2295
rect 31803 2261 31812 2295
rect 31760 2252 31812 2261
rect 32404 2295 32456 2304
rect 32404 2261 32413 2295
rect 32413 2261 32447 2295
rect 32447 2261 32456 2295
rect 32404 2252 32456 2261
rect 117412 2295 117464 2304
rect 117412 2261 117421 2295
rect 117421 2261 117455 2295
rect 117455 2261 117464 2295
rect 117412 2252 117464 2261
rect 120816 2295 120868 2304
rect 120816 2261 120825 2295
rect 120825 2261 120859 2295
rect 120859 2261 120868 2295
rect 120816 2252 120868 2261
rect 121368 2295 121420 2304
rect 121368 2261 121377 2295
rect 121377 2261 121411 2295
rect 121411 2261 121420 2295
rect 121368 2252 121420 2261
rect 123852 2295 123904 2304
rect 123852 2261 123861 2295
rect 123861 2261 123895 2295
rect 123895 2261 123904 2295
rect 123852 2252 123904 2261
rect 124404 2295 124456 2304
rect 124404 2261 124413 2295
rect 124413 2261 124447 2295
rect 124447 2261 124456 2295
rect 124404 2252 124456 2261
rect 125324 2295 125376 2304
rect 125324 2261 125333 2295
rect 125333 2261 125367 2295
rect 125367 2261 125376 2295
rect 125324 2252 125376 2261
rect 128544 2295 128596 2304
rect 128544 2261 128553 2295
rect 128553 2261 128587 2295
rect 128587 2261 128596 2295
rect 128544 2252 128596 2261
rect 135260 2252 135312 2304
rect 140872 2320 140924 2372
rect 141700 2363 141752 2372
rect 141700 2329 141740 2363
rect 141740 2329 141752 2363
rect 141700 2320 141752 2329
rect 141976 2320 142028 2372
rect 145932 2363 145984 2372
rect 145932 2329 145966 2363
rect 145966 2329 145984 2363
rect 145932 2320 145984 2329
rect 147680 2431 147732 2440
rect 147680 2397 147689 2431
rect 147689 2397 147723 2431
rect 147723 2397 147732 2431
rect 147680 2388 147732 2397
rect 140596 2295 140648 2304
rect 140596 2261 140605 2295
rect 140605 2261 140639 2295
rect 140639 2261 140648 2295
rect 140596 2252 140648 2261
rect 147496 2295 147548 2304
rect 147496 2261 147505 2295
rect 147505 2261 147539 2295
rect 147539 2261 147548 2295
rect 147496 2252 147548 2261
rect 147864 2252 147916 2304
rect 148048 2456 148100 2508
rect 149704 2456 149756 2508
rect 154120 2499 154172 2508
rect 154120 2465 154129 2499
rect 154129 2465 154163 2499
rect 154163 2465 154172 2499
rect 154120 2456 154172 2465
rect 155776 2524 155828 2576
rect 155960 2524 156012 2576
rect 157432 2524 157484 2576
rect 157156 2456 157208 2508
rect 148784 2388 148836 2440
rect 150348 2388 150400 2440
rect 154304 2431 154356 2440
rect 154304 2397 154313 2431
rect 154313 2397 154347 2431
rect 154347 2397 154356 2431
rect 154304 2388 154356 2397
rect 155132 2431 155184 2440
rect 155132 2397 155141 2431
rect 155141 2397 155175 2431
rect 155175 2397 155184 2431
rect 155132 2388 155184 2397
rect 155868 2388 155920 2440
rect 149152 2320 149204 2372
rect 151084 2320 151136 2372
rect 149612 2295 149664 2304
rect 149612 2261 149621 2295
rect 149621 2261 149655 2295
rect 149655 2261 149664 2295
rect 149612 2252 149664 2261
rect 151728 2252 151780 2304
rect 155868 2252 155920 2304
rect 156604 2295 156656 2304
rect 156604 2261 156613 2295
rect 156613 2261 156647 2295
rect 156647 2261 156656 2295
rect 156604 2252 156656 2261
rect 157800 2295 157852 2304
rect 157800 2261 157809 2295
rect 157809 2261 157843 2295
rect 157843 2261 157852 2295
rect 157800 2252 157852 2261
rect 40394 2150 40446 2202
rect 40458 2150 40510 2202
rect 40522 2150 40574 2202
rect 40586 2150 40638 2202
rect 40650 2150 40702 2202
rect 79839 2150 79891 2202
rect 79903 2150 79955 2202
rect 79967 2150 80019 2202
rect 80031 2150 80083 2202
rect 80095 2150 80147 2202
rect 119284 2150 119336 2202
rect 119348 2150 119400 2202
rect 119412 2150 119464 2202
rect 119476 2150 119528 2202
rect 119540 2150 119592 2202
rect 158729 2150 158781 2202
rect 158793 2150 158845 2202
rect 158857 2150 158909 2202
rect 158921 2150 158973 2202
rect 158985 2150 159037 2202
rect 10968 2048 11020 2100
rect 32404 2048 32456 2100
rect 120172 2048 120224 2100
rect 124404 2048 124456 2100
rect 128544 2048 128596 2100
rect 145932 2048 145984 2100
rect 146668 2048 146720 2100
rect 149060 2048 149112 2100
rect 150256 2048 150308 2100
rect 156604 2048 156656 2100
rect 15568 1980 15620 2032
rect 31760 1980 31812 2032
rect 121368 1980 121420 2032
rect 134064 1980 134116 2032
rect 136640 1980 136692 2032
rect 150348 1980 150400 2032
rect 106556 1912 106608 1964
rect 123852 1912 123904 1964
rect 124864 1912 124916 1964
rect 147496 1912 147548 1964
rect 149152 1912 149204 1964
rect 159180 1912 159232 1964
rect 146116 1844 146168 1896
rect 146668 1844 146720 1896
rect 114468 1776 114520 1828
rect 115572 1640 115624 1692
rect 124404 1776 124456 1828
rect 130844 1776 130896 1828
rect 141976 1776 142028 1828
rect 147772 1776 147824 1828
rect 147864 1776 147916 1828
rect 156052 1776 156104 1828
rect 123024 1708 123076 1760
rect 140596 1708 140648 1760
rect 143632 1708 143684 1760
rect 154948 1708 155000 1760
rect 125324 1640 125376 1692
rect 142804 1640 142856 1692
rect 146208 1640 146260 1692
rect 155132 1640 155184 1692
rect 120816 1572 120868 1624
rect 136088 1572 136140 1624
rect 144000 1572 144052 1624
rect 155960 1572 156012 1624
rect 126980 1504 127032 1556
rect 147772 1504 147824 1556
rect 156972 1504 157024 1556
rect 125324 1436 125376 1488
rect 110236 1300 110288 1352
rect 152004 1300 152056 1352
rect 115204 1232 115256 1284
rect 150900 1232 150952 1284
rect 121184 1164 121236 1216
rect 155408 1164 155460 1216
rect 119804 1096 119856 1148
rect 150808 1096 150860 1148
rect 101956 1028 102008 1080
rect 128452 1028 128504 1080
rect 129188 1028 129240 1080
rect 151176 1028 151228 1080
rect 113548 960 113600 1012
rect 138112 960 138164 1012
<< metal2 >>
rect 9586 15314 9642 16000
rect 9232 15286 9642 15314
rect 4068 13864 4120 13870
rect 4066 13832 4068 13841
rect 4120 13832 4122 13841
rect 4066 13767 4122 13776
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13530 7880 13670
rect 9232 13530 9260 15286
rect 9586 15200 9642 15286
rect 10138 15200 10194 16000
rect 10690 15314 10746 16000
rect 10520 15286 10746 15314
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 10060 13462 10088 13942
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12986 9444 13262
rect 10152 12986 10180 15200
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10428 13326 10456 13738
rect 10232 13320 10284 13326
rect 10230 13288 10232 13297
rect 10416 13320 10468 13326
rect 10284 13288 10286 13297
rect 10416 13262 10468 13268
rect 10230 13223 10286 13232
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12306 10088 12650
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 5724 12232 5776 12238
rect 9864 12232 9916 12238
rect 5724 12174 5776 12180
rect 9862 12200 9864 12209
rect 9916 12200 9918 12209
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 10606 3832 11630
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10062 3832 10542
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9897 1624 9930
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 1596 9722 1624 9823
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 3804 9586 3832 9998
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4080 6662 4108 11698
rect 4172 10742 4200 12038
rect 4448 11354 4476 12174
rect 5736 11558 5764 12174
rect 6828 12164 6880 12170
rect 9862 12135 9918 12144
rect 6828 12106 6880 12112
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7410 4844 7686
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 5953 1624 6258
rect 1582 5944 1638 5953
rect 1582 5879 1638 5888
rect 4632 5710 4660 7142
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 3896 5302 3924 5646
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 2446 1716 2790
rect 4724 2650 4752 6734
rect 4908 5914 4936 11154
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 4826 5028 9930
rect 5184 9654 5212 10406
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5184 8634 5212 9590
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7410 5120 8230
rect 5276 7546 5304 8842
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5184 4758 5212 4966
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5368 4622 5396 8298
rect 5460 7954 5488 9862
rect 5552 8498 5580 11494
rect 5736 10810 5764 11494
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5736 10266 5764 10746
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5736 10062 5764 10202
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9722 5764 9998
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5644 7886 5672 8366
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5736 5914 5764 9522
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5828 8634 5856 8910
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 7546 6040 7822
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5920 5234 5948 5306
rect 6012 5234 6040 6054
rect 6104 5710 6132 11562
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6656 5370 6684 7754
rect 6748 7546 6776 8298
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 4826 6040 5170
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 6840 4010 6868 12106
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11150 7788 11494
rect 8404 11286 8432 11698
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 9600 11150 9628 12038
rect 10060 11558 10088 12242
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11626 10364 12174
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 8220 10470 8248 11086
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 9994 8248 10406
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 6458 8064 9318
rect 8220 8362 8248 9930
rect 8404 9926 8432 10610
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8404 7818 8432 9862
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8680 6254 8708 8230
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 9324 6186 9352 10610
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 4146 9168 6054
rect 9600 4146 9628 11086
rect 10060 10470 10088 11494
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 9654 10088 10406
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10336 6225 10364 11562
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5166 9720 5510
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 10428 4282 10456 12786
rect 10520 12442 10548 15286
rect 10690 15200 10746 15286
rect 11242 15200 11298 16000
rect 11794 15200 11850 16000
rect 12346 15200 12402 16000
rect 12898 15314 12954 16000
rect 12636 15286 12954 15314
rect 11256 14006 11284 15200
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12782 10824 13126
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10690 11656 10746 11665
rect 10690 11591 10746 11600
rect 10506 11248 10562 11257
rect 10704 11218 10732 11591
rect 10506 11183 10508 11192
rect 10560 11183 10562 11192
rect 10692 11212 10744 11218
rect 10508 11154 10560 11160
rect 10692 11154 10744 11160
rect 10704 9110 10732 11154
rect 10888 11150 10916 12786
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12306 11008 12718
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11072 11082 11100 12174
rect 11164 11082 11192 13262
rect 11808 12986 11836 15200
rect 12360 13530 12388 15200
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12544 13394 12572 13874
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12646 11928 13262
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11992 12850 12020 12922
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11256 11354 11284 11698
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11072 10810 11100 11018
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10704 8294 10732 9046
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 8090 10732 8230
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5828 2446 5856 2790
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 1688 2009 1716 2382
rect 10980 2106 11008 4082
rect 11072 3194 11100 9114
rect 11440 8974 11468 10950
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 6254 11192 7278
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11072 2446 11100 3130
rect 11164 2650 11192 6190
rect 11440 3194 11468 8910
rect 11716 6662 11744 12106
rect 11886 11792 11942 11801
rect 11886 11727 11888 11736
rect 11940 11727 11942 11736
rect 11888 11698 11940 11704
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11808 5710 11836 9862
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11164 2514 11192 2586
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11716 2378 11744 3878
rect 11900 2650 11928 11086
rect 11992 8362 12020 12786
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12084 12345 12112 12378
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 10742 12112 11494
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12176 9330 12204 13262
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12268 10810 12296 11086
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12360 9586 12388 12582
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 10577 12480 12271
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12438 10568 12494 10577
rect 12438 10503 12494 10512
rect 12544 9994 12572 11698
rect 12636 11694 12664 15286
rect 12898 15200 12954 15286
rect 13450 15200 13506 16000
rect 14002 15200 14058 16000
rect 14554 15200 14610 16000
rect 15106 15200 15162 16000
rect 15658 15200 15714 16000
rect 16210 15200 16266 16000
rect 16762 15200 16818 16000
rect 17314 15314 17370 16000
rect 17314 15286 17540 15314
rect 17314 15200 17370 15286
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13326 12756 13670
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12176 9302 12296 9330
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12176 4622 12204 8774
rect 12268 6118 12296 9302
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12360 4826 12388 8774
rect 12452 8634 12480 8910
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12728 7274 12756 13262
rect 13464 12714 13492 15200
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13924 12986 13952 13194
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 12900 11688 12952 11694
rect 12898 11656 12900 11665
rect 12952 11656 12954 11665
rect 12898 11591 12954 11600
rect 13096 10062 13124 12582
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 11898 13216 12174
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13372 11762 13400 12582
rect 14016 12442 14044 15200
rect 14568 13462 14596 15200
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 15120 13258 15148 15200
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 13802 15332 13874
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13358 10568 13414 10577
rect 13358 10503 13414 10512
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12912 8090 12940 8570
rect 13280 8566 13308 9862
rect 13372 8922 13400 10503
rect 13556 10010 13584 12174
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13648 11014 13676 11290
rect 14108 11257 14136 12378
rect 14292 11898 14320 13126
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15028 12782 15056 12922
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14832 12232 14884 12238
rect 14830 12200 14832 12209
rect 14884 12200 14886 12209
rect 14464 12164 14516 12170
rect 14830 12135 14886 12144
rect 14464 12106 14516 12112
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14476 11762 14504 12106
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11830 14964 12038
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15212 11762 15240 13738
rect 15672 13530 15700 15200
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 14094 11248 14150 11257
rect 14094 11183 14150 11192
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10470 13676 10610
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 10198 13676 10406
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 13556 9982 13676 10010
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13464 9042 13492 9590
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13372 8894 13492 8922
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5234 13032 5510
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4826 12664 4966
rect 13280 4826 13308 6734
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12636 4554 12664 4762
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12636 3942 12664 4150
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3602 13308 3878
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13372 3126 13400 7686
rect 13464 7410 13492 8894
rect 13556 7886 13584 9862
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 7002 13492 7346
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13648 5166 13676 9982
rect 14200 9586 14228 10066
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9654 14320 9998
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 8090 13768 8434
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 6730 13768 7754
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 5370 13768 6666
rect 14016 6322 14044 7686
rect 14108 7546 14136 9522
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14278 9072 14334 9081
rect 14278 9007 14280 9016
rect 14332 9007 14334 9016
rect 14280 8978 14332 8984
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 8090 14320 8230
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14384 6798 14412 8774
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 3942 13584 4558
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13556 3058 13584 3334
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 13648 2582 13676 4626
rect 13832 4622 13860 5306
rect 14292 5302 14320 5646
rect 14476 5642 14504 9318
rect 14568 6662 14596 11698
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10554 15240 11086
rect 15304 10810 15332 13194
rect 15764 12986 15792 13262
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15580 12238 15608 12922
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15120 10526 15240 10554
rect 15120 10062 15148 10526
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7002 14872 7822
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14292 5030 14320 5238
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13820 4616 13872 4622
rect 13872 4576 14044 4604
rect 13820 4558 13872 4564
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4298 13860 4422
rect 13740 4270 13860 4298
rect 13740 4078 13768 4270
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13832 2990 13860 4082
rect 13924 3194 13952 4082
rect 14016 3738 14044 4576
rect 14292 4214 14320 4966
rect 14384 4826 14412 5578
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14016 3466 14044 3674
rect 14476 3534 14504 4694
rect 14844 4690 14872 6938
rect 14936 6458 14964 8434
rect 15028 7886 15056 9454
rect 15120 9042 15148 9998
rect 15396 9654 15424 10610
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15120 7546 15148 8978
rect 15488 7818 15516 11698
rect 15580 9586 15608 11766
rect 15672 10538 15700 12106
rect 15856 11558 15884 12854
rect 16224 12322 16252 15200
rect 16394 13288 16450 13297
rect 16394 13223 16450 13232
rect 16408 13190 16436 13223
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16776 12986 16804 15200
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13326 17448 13670
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17512 12986 17540 15286
rect 17866 15200 17922 16000
rect 18418 15200 18474 16000
rect 18970 15314 19026 16000
rect 18708 15286 19026 15314
rect 17880 13530 17908 15200
rect 18432 13530 18460 15200
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17696 12850 17724 13194
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17236 12434 17264 12718
rect 16132 12294 16252 12322
rect 17052 12406 17264 12434
rect 18616 12434 18644 13262
rect 18708 12986 18736 15286
rect 18970 15200 19026 15286
rect 19522 15200 19578 16000
rect 20074 15200 20130 16000
rect 20626 15314 20682 16000
rect 20548 15286 20682 15314
rect 19536 13530 19564 15200
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 18616 12406 18828 12434
rect 16132 12102 16160 12294
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15934 11792 15990 11801
rect 15934 11727 15990 11736
rect 16120 11756 16172 11762
rect 15948 11558 15976 11727
rect 16120 11698 16172 11704
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15028 6322 15056 6734
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15028 5642 15056 6258
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15028 5234 15056 5578
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4826 14964 4966
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 15028 4486 15056 5170
rect 15120 4826 15148 6802
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15212 5914 15240 6258
rect 15304 6186 15332 6734
rect 15672 6458 15700 8842
rect 15764 8294 15792 9522
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15856 7954 15884 11494
rect 16132 8838 16160 11698
rect 16224 11218 16252 12174
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15580 5166 15608 5510
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14016 3194 14044 3402
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14476 2990 14504 3470
rect 15120 3126 15148 4762
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 13832 2650 13860 2926
rect 15212 2922 15240 3878
rect 15580 3398 15608 5102
rect 15672 4146 15700 6258
rect 15856 5166 15884 7210
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 16132 3738 16160 7822
rect 16316 7750 16344 12106
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16960 10742 16988 12038
rect 17052 11694 17080 12406
rect 17958 12200 18014 12209
rect 17958 12135 18014 12144
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11762 17264 12038
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8514 16528 8774
rect 16408 8498 16528 8514
rect 16408 8492 16540 8498
rect 16408 8486 16488 8492
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16408 7478 16436 8486
rect 16488 8434 16540 8440
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16500 6798 16528 8298
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16592 5914 16620 10610
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10062 16712 10406
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16684 9586 16712 9998
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16776 9058 16804 10134
rect 16960 10130 16988 10678
rect 17052 10674 17080 11630
rect 17592 11280 17644 11286
rect 17592 11222 17644 11228
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17222 10704 17278 10713
rect 17040 10668 17092 10674
rect 17222 10639 17278 10648
rect 17040 10610 17092 10616
rect 17052 10130 17080 10610
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16684 9030 16804 9058
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16302 5400 16358 5409
rect 16302 5335 16304 5344
rect 16356 5335 16358 5344
rect 16304 5306 16356 5312
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16316 3670 16344 5306
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16316 3466 16344 3606
rect 16684 3534 16712 9030
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8430 16804 8910
rect 16868 8430 16896 9930
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16946 9072 17002 9081
rect 16946 9007 16948 9016
rect 17000 9007 17002 9016
rect 16948 8978 17000 8984
rect 16764 8424 16816 8430
rect 16762 8392 16764 8401
rect 16856 8424 16908 8430
rect 16816 8392 16818 8401
rect 16856 8366 16908 8372
rect 16762 8327 16818 8336
rect 16868 7410 16896 8366
rect 16960 8294 16988 8978
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16868 6746 16896 7346
rect 16776 6718 17080 6746
rect 16776 5574 16804 6718
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5370 16804 5510
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16776 4214 16804 5306
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 15580 2038 15608 3334
rect 16868 3058 16896 6598
rect 17052 6322 17080 6718
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16960 5302 16988 6258
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5574 17080 6054
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17040 4616 17092 4622
rect 17144 4604 17172 9862
rect 17236 9586 17264 10639
rect 17328 10198 17356 11154
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 6662 17264 9522
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17328 5846 17356 8230
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17328 5409 17356 5646
rect 17314 5400 17370 5409
rect 17314 5335 17370 5344
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17236 5098 17264 5170
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 17092 4576 17172 4604
rect 17040 4558 17092 4564
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17420 2446 17448 9318
rect 17512 6390 17540 9318
rect 17604 8906 17632 11222
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17696 9042 17724 9114
rect 17788 9110 17816 9590
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17696 8786 17724 8978
rect 17788 8974 17816 9046
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17604 8758 17724 8786
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17512 5846 17540 6190
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17604 3466 17632 8758
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17696 8378 17724 8434
rect 17696 8362 17816 8378
rect 17696 8356 17828 8362
rect 17696 8350 17776 8356
rect 17776 8298 17828 8304
rect 17880 8090 17908 8434
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 4146 17724 6054
rect 17788 5710 17816 7278
rect 17880 6934 17908 7346
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17972 4622 18000 12135
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18156 10130 18184 11630
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18340 11206 18552 11234
rect 18340 11082 18368 11206
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18432 11014 18460 11086
rect 18524 11082 18552 11206
rect 18616 11150 18644 11562
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10810 18644 10950
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 6322 18092 8774
rect 18156 7886 18184 10066
rect 18524 9994 18552 10474
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18248 8498 18276 8570
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18616 8090 18644 9046
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8634 18736 8774
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18616 7478 18644 8026
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18156 5370 18184 5850
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4826 18276 4966
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17880 4486 17908 4558
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4146 17908 4422
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 2854 18000 3334
rect 18248 3058 18276 3470
rect 18340 3126 18368 7142
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18524 6254 18552 6734
rect 18800 6322 18828 12406
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 7274 18920 12038
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18984 7954 19012 8230
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6458 18920 6598
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18892 5914 18920 6394
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18432 3466 18460 3878
rect 18524 3534 18552 4082
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18616 3126 18644 5510
rect 18708 5370 18736 5510
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18880 4480 18932 4486
rect 18984 4468 19012 7686
rect 19168 7274 19196 12718
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11694 19288 12038
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19352 11121 19380 11494
rect 19444 11218 19472 12174
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19444 10810 19472 11154
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19340 10056 19392 10062
rect 19392 10004 19472 10010
rect 19340 9998 19472 10004
rect 19352 9982 19472 9998
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9654 19380 9862
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19444 9586 19472 9982
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18932 4440 19012 4468
rect 18880 4422 18932 4428
rect 18892 4214 18920 4422
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 19260 4162 19288 7142
rect 19352 6186 19380 8842
rect 19444 8634 19472 8978
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19430 8392 19486 8401
rect 19430 8327 19486 8336
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19444 4758 19472 8327
rect 19536 5914 19564 9454
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19536 4282 19564 4422
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18800 3194 18828 4082
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17972 2650 18000 2790
rect 18892 2666 18920 4150
rect 19260 4134 19564 4162
rect 19536 4078 19564 4134
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2854 19380 2994
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 18800 2650 18920 2666
rect 19628 2650 19656 13738
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19812 12434 19840 12718
rect 19720 12406 19840 12434
rect 19720 4826 19748 12406
rect 19904 12374 19932 13262
rect 20088 12986 20116 15200
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19892 12368 19944 12374
rect 19812 12316 19892 12322
rect 19812 12310 19944 12316
rect 19812 12294 19932 12310
rect 19812 11830 19840 12294
rect 20180 11898 20208 12922
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 20364 11642 20392 13262
rect 20548 11898 20576 15286
rect 20626 15200 20682 15286
rect 21178 15200 21234 16000
rect 21730 15200 21786 16000
rect 22282 15200 22338 16000
rect 22834 15200 22890 16000
rect 23386 15200 23442 16000
rect 23938 15200 23994 16000
rect 24490 15200 24546 16000
rect 25042 15314 25098 16000
rect 25594 15314 25650 16000
rect 26146 15314 26202 16000
rect 26698 15314 26754 16000
rect 24872 15286 25098 15314
rect 20672 13628 20980 13637
rect 20672 13626 20678 13628
rect 20734 13626 20758 13628
rect 20814 13626 20838 13628
rect 20894 13626 20918 13628
rect 20974 13626 20980 13628
rect 20734 13574 20736 13626
rect 20916 13574 20918 13626
rect 20672 13572 20678 13574
rect 20734 13572 20758 13574
rect 20814 13572 20838 13574
rect 20894 13572 20918 13574
rect 20974 13572 20980 13574
rect 20672 13563 20980 13572
rect 21192 13462 21220 15200
rect 21744 13530 21772 15200
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21640 13456 21692 13462
rect 22008 13456 22060 13462
rect 21692 13404 22008 13410
rect 21640 13398 22060 13404
rect 21652 13382 22048 13398
rect 21456 13320 21508 13326
rect 21508 13280 21680 13308
rect 21456 13262 21508 13268
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21376 13161 21404 13194
rect 21548 13184 21600 13190
rect 21362 13152 21418 13161
rect 21548 13126 21600 13132
rect 21362 13087 21418 13096
rect 21456 12776 21508 12782
rect 21560 12753 21588 13126
rect 21456 12718 21508 12724
rect 21546 12744 21602 12753
rect 20672 12540 20980 12549
rect 20672 12538 20678 12540
rect 20734 12538 20758 12540
rect 20814 12538 20838 12540
rect 20894 12538 20918 12540
rect 20974 12538 20980 12540
rect 20734 12486 20736 12538
rect 20916 12486 20918 12538
rect 20672 12484 20678 12486
rect 20734 12484 20758 12486
rect 20814 12484 20838 12486
rect 20894 12484 20918 12486
rect 20974 12484 20980 12486
rect 20672 12475 20980 12484
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20640 11665 20668 12310
rect 21468 12238 21496 12718
rect 21546 12679 21602 12688
rect 21652 12434 21680 13280
rect 22204 13258 22232 13466
rect 22296 13462 22324 15200
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22112 12442 22140 12718
rect 22100 12436 22152 12442
rect 21652 12406 21772 12434
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 20732 12102 20760 12174
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 20180 11614 20392 11642
rect 20626 11656 20682 11665
rect 20180 11558 20208 11614
rect 20626 11591 20682 11600
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19798 9480 19854 9489
rect 19798 9415 19800 9424
rect 19852 9415 19854 9424
rect 19800 9386 19852 9392
rect 19904 9382 19932 9522
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19996 8430 20024 10406
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20088 9926 20116 10202
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20088 9518 20116 9862
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19812 5710 19840 8366
rect 20088 7970 20116 9454
rect 19996 7942 20116 7970
rect 19996 7154 20024 7942
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19904 7126 20024 7154
rect 19904 6866 19932 7126
rect 20088 6866 20116 7822
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19904 5370 19932 6666
rect 20088 6458 20116 6802
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5710 20024 6054
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 20088 4146 20116 6394
rect 20180 4282 20208 11494
rect 20272 11082 20300 11494
rect 20672 11452 20980 11461
rect 20672 11450 20678 11452
rect 20734 11450 20758 11452
rect 20814 11450 20838 11452
rect 20894 11450 20918 11452
rect 20974 11450 20980 11452
rect 20734 11398 20736 11450
rect 20916 11398 20918 11450
rect 20672 11396 20678 11398
rect 20734 11396 20758 11398
rect 20814 11396 20838 11398
rect 20894 11396 20918 11398
rect 20974 11396 20980 11398
rect 20672 11387 20980 11396
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20548 10810 20576 11154
rect 21100 11150 21128 11698
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20548 9654 20576 10746
rect 21376 10470 21404 11018
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 20672 10364 20980 10373
rect 20672 10362 20678 10364
rect 20734 10362 20758 10364
rect 20814 10362 20838 10364
rect 20894 10362 20918 10364
rect 20974 10362 20980 10364
rect 20734 10310 20736 10362
rect 20916 10310 20918 10362
rect 20672 10308 20678 10310
rect 20734 10308 20758 10310
rect 20814 10308 20838 10310
rect 20894 10308 20918 10310
rect 20974 10308 20980 10310
rect 20672 10299 20980 10308
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20672 9276 20980 9285
rect 20672 9274 20678 9276
rect 20734 9274 20758 9276
rect 20814 9274 20838 9276
rect 20894 9274 20918 9276
rect 20974 9274 20980 9276
rect 20734 9222 20736 9274
rect 20916 9222 20918 9274
rect 20672 9220 20678 9222
rect 20734 9220 20758 9222
rect 20814 9220 20838 9222
rect 20894 9220 20918 9222
rect 20974 9220 20980 9222
rect 20672 9211 20980 9220
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20672 8188 20980 8197
rect 20672 8186 20678 8188
rect 20734 8186 20758 8188
rect 20814 8186 20838 8188
rect 20894 8186 20918 8188
rect 20974 8186 20980 8188
rect 20734 8134 20736 8186
rect 20916 8134 20918 8186
rect 20672 8132 20678 8134
rect 20734 8132 20758 8134
rect 20814 8132 20838 8134
rect 20894 8132 20918 8134
rect 20974 8132 20980 8134
rect 20672 8123 20980 8132
rect 21008 7426 21036 8774
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7546 21128 7754
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21008 7398 21128 7426
rect 20672 7100 20980 7109
rect 20672 7098 20678 7100
rect 20734 7098 20758 7100
rect 20814 7098 20838 7100
rect 20894 7098 20918 7100
rect 20974 7098 20980 7100
rect 20734 7046 20736 7098
rect 20916 7046 20918 7098
rect 20672 7044 20678 7046
rect 20734 7044 20758 7046
rect 20814 7044 20838 7046
rect 20894 7044 20918 7046
rect 20974 7044 20980 7046
rect 20672 7035 20980 7044
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20272 6458 20300 6938
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20272 6202 20300 6394
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20352 6248 20404 6254
rect 20272 6196 20352 6202
rect 20272 6190 20404 6196
rect 20272 6174 20392 6190
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 5778 20300 6054
rect 20364 5914 20392 6174
rect 20672 6012 20980 6021
rect 20672 6010 20678 6012
rect 20734 6010 20758 6012
rect 20814 6010 20838 6012
rect 20894 6010 20918 6012
rect 20974 6010 20980 6012
rect 20734 5958 20736 6010
rect 20916 5958 20918 6010
rect 20672 5956 20678 5958
rect 20734 5956 20758 5958
rect 20814 5956 20838 5958
rect 20894 5956 20918 5958
rect 20974 5956 20980 5958
rect 20672 5947 20980 5956
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20672 4924 20980 4933
rect 20672 4922 20678 4924
rect 20734 4922 20758 4924
rect 20814 4922 20838 4924
rect 20894 4922 20918 4924
rect 20974 4922 20980 4924
rect 20734 4870 20736 4922
rect 20916 4870 20918 4922
rect 20672 4868 20678 4870
rect 20734 4868 20758 4870
rect 20814 4868 20838 4870
rect 20894 4868 20918 4870
rect 20974 4868 20980 4870
rect 20672 4859 20980 4868
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20088 3534 20116 4082
rect 20456 3738 20484 4082
rect 20672 3836 20980 3845
rect 20672 3834 20678 3836
rect 20734 3834 20758 3836
rect 20814 3834 20838 3836
rect 20894 3834 20918 3836
rect 20974 3834 20980 3836
rect 20734 3782 20736 3834
rect 20916 3782 20918 3834
rect 20672 3780 20678 3782
rect 20734 3780 20758 3782
rect 20814 3780 20838 3782
rect 20894 3780 20918 3782
rect 20974 3780 20980 3782
rect 20672 3771 20980 3780
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18788 2644 18920 2650
rect 18840 2638 18920 2644
rect 19616 2644 19668 2650
rect 18788 2586 18840 2592
rect 19616 2586 19668 2592
rect 19904 2582 19932 3402
rect 20088 3194 20116 3470
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20536 3120 20588 3126
rect 20534 3088 20536 3097
rect 20588 3088 20590 3097
rect 20534 3023 20590 3032
rect 20732 2922 20760 3606
rect 21008 3074 21036 6326
rect 21100 5642 21128 7398
rect 21192 6798 21220 8910
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21284 6458 21312 7822
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 20824 3058 21036 3074
rect 20812 3052 21036 3058
rect 20864 3046 21036 3052
rect 20812 2994 20864 3000
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20672 2748 20980 2757
rect 20672 2746 20678 2748
rect 20734 2746 20758 2748
rect 20814 2746 20838 2748
rect 20894 2746 20918 2748
rect 20974 2746 20980 2748
rect 20734 2694 20736 2746
rect 20916 2694 20918 2746
rect 20672 2692 20678 2694
rect 20734 2692 20758 2694
rect 20814 2692 20838 2694
rect 20894 2692 20918 2694
rect 20974 2692 20980 2694
rect 20672 2683 20980 2692
rect 19892 2576 19944 2582
rect 19892 2518 19944 2524
rect 21100 2446 21128 5578
rect 21376 5302 21404 10406
rect 21652 7410 21680 11834
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 6866 21772 12406
rect 22100 12378 22152 12384
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21928 11082 21956 11766
rect 22204 11762 22232 12786
rect 22388 12714 22416 13670
rect 22742 12880 22798 12889
rect 22742 12815 22744 12824
rect 22796 12815 22798 12824
rect 22744 12786 22796 12792
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22848 12442 22876 15200
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 11082 22140 11494
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10810 22048 10950
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22204 10606 22232 11698
rect 22466 11656 22522 11665
rect 22466 11591 22522 11600
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21914 8528 21970 8537
rect 21914 8463 21970 8472
rect 21928 8362 21956 8463
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 22296 8242 22324 11494
rect 22112 8214 22324 8242
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 6458 21496 6598
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21192 4214 21220 4558
rect 21652 4554 21680 6258
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21180 4208 21232 4214
rect 21180 4150 21232 4156
rect 21192 3942 21220 4150
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21192 2514 21220 3878
rect 21652 3670 21680 4490
rect 21836 4486 21864 7346
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22020 5914 22048 6190
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22020 5778 22048 5850
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22112 5681 22140 8214
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22204 6322 22232 8026
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22098 5672 22154 5681
rect 22098 5607 22154 5616
rect 22112 5574 22140 5607
rect 22204 5574 22232 6054
rect 22388 5710 22416 6054
rect 22480 5914 22508 11591
rect 23032 10606 23060 12786
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 6662 22600 7142
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 21928 4486 21956 5034
rect 22480 4758 22508 5102
rect 22572 5098 22600 6598
rect 23032 5302 23060 7686
rect 23308 7546 23336 13262
rect 23400 12986 23428 15200
rect 23952 13530 23980 15200
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23768 12646 23796 13262
rect 24030 12744 24086 12753
rect 24030 12679 24032 12688
rect 24084 12679 24086 12688
rect 24032 12650 24084 12656
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23768 12434 23796 12582
rect 24504 12442 24532 15200
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24768 13796 24820 13802
rect 24768 13738 24820 13744
rect 24596 13530 24624 13738
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24780 13190 24808 13738
rect 24768 13184 24820 13190
rect 24688 13132 24768 13138
rect 24688 13126 24820 13132
rect 24688 13110 24808 13126
rect 23676 12406 23796 12434
rect 24492 12436 24544 12442
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 8090 23428 9590
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23296 6180 23348 6186
rect 23296 6122 23348 6128
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 22468 4752 22520 4758
rect 22468 4694 22520 4700
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21836 3738 21864 4422
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 22572 3534 22600 5034
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4690 22692 4966
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 23308 3738 23336 6122
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22480 2922 22508 3062
rect 22572 3058 22600 3470
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 23584 2446 23612 6666
rect 23676 4214 23704 12406
rect 24492 12378 24544 12384
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24136 11762 24164 12038
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23768 10470 23796 11630
rect 24412 11218 24440 12310
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 24596 11150 24624 12174
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23768 10266 23796 10406
rect 24596 10266 24624 11086
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24216 8288 24268 8294
rect 24216 8230 24268 8236
rect 24228 8022 24256 8230
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23768 6118 23796 6394
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23860 4690 23888 6598
rect 23952 6390 23980 7278
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24044 5642 24072 5850
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 24032 5636 24084 5642
rect 24032 5578 24084 5584
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 23952 3194 23980 5578
rect 24688 5386 24716 13110
rect 24872 13002 24900 15286
rect 25042 15200 25098 15286
rect 25240 15286 25650 15314
rect 25240 13462 25268 15286
rect 25594 15200 25650 15286
rect 25792 15286 26202 15314
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24964 13190 24992 13330
rect 25792 13326 25820 15286
rect 26146 15200 26202 15286
rect 26436 15286 26754 15314
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24780 12986 24900 13002
rect 25056 12986 25084 13262
rect 24768 12980 24900 12986
rect 24820 12974 24900 12980
rect 25044 12980 25096 12986
rect 24768 12922 24820 12928
rect 25044 12922 25096 12928
rect 25148 12434 25176 13262
rect 26436 12986 26464 15286
rect 26698 15200 26754 15286
rect 27250 15200 27306 16000
rect 27802 15200 27858 16000
rect 28354 15314 28410 16000
rect 28092 15286 28410 15314
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 26516 13184 26568 13190
rect 26700 13184 26752 13190
rect 26568 13132 26700 13138
rect 26516 13126 26752 13132
rect 26528 13110 26740 13126
rect 26804 12986 26832 13330
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25424 12434 25452 12718
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 24964 12406 25452 12434
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24872 5914 24900 12106
rect 24964 11762 24992 12406
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 25608 11354 25636 12650
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25148 10810 25176 11018
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25148 10062 25176 10746
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25608 6662 25636 10406
rect 25700 9926 25728 12786
rect 26148 12776 26200 12782
rect 26252 12753 26280 12922
rect 26148 12718 26200 12724
rect 26238 12744 26294 12753
rect 26160 12374 26188 12718
rect 26238 12679 26294 12688
rect 27264 12442 27292 15200
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27448 12646 27476 13466
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 26148 12368 26200 12374
rect 26148 12310 26200 12316
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26976 12164 27028 12170
rect 26976 12106 27028 12112
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 25792 5778 25820 12038
rect 26620 11694 26648 12106
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26608 11688 26660 11694
rect 26608 11630 26660 11636
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 24596 5358 24716 5386
rect 24596 4146 24624 5358
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24688 5030 24716 5170
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4826 24716 4966
rect 25240 4826 25268 5714
rect 25504 5364 25556 5370
rect 25504 5306 25556 5312
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 3194 24440 3334
rect 24688 3194 24716 4762
rect 25240 4690 25268 4762
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 3670 24808 4422
rect 25240 3738 25268 4626
rect 25332 4622 25360 4966
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 25240 3534 25268 3674
rect 25516 3534 25544 5306
rect 25792 4554 25820 5714
rect 25780 4548 25832 4554
rect 25780 4490 25832 4496
rect 25884 3738 25912 7822
rect 25976 5370 26004 11562
rect 26252 11082 26280 11630
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26056 8832 26108 8838
rect 26056 8774 26108 8780
rect 26068 5574 26096 8774
rect 26252 8378 26280 11018
rect 26620 10810 26648 11086
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26896 10985 26924 11018
rect 26882 10976 26938 10985
rect 26882 10911 26938 10920
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26344 9178 26372 9454
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26528 9178 26556 9318
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26344 8498 26372 9114
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26252 8350 26372 8378
rect 26344 7342 26372 8350
rect 26620 7410 26648 10746
rect 26988 10470 27016 12106
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26332 7336 26384 7342
rect 26332 7278 26384 7284
rect 26344 6866 26372 7278
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 23952 2990 23980 3130
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24412 2514 24440 3130
rect 24780 3097 24808 3130
rect 24766 3088 24822 3097
rect 24766 3023 24822 3032
rect 26068 2774 26096 5510
rect 26252 4486 26280 6598
rect 26344 6254 26372 6802
rect 26896 6662 26924 9522
rect 27080 9450 27108 11494
rect 27356 11082 27384 12174
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27344 11076 27396 11082
rect 27344 11018 27396 11024
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 27172 8974 27200 11018
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10742 27292 10950
rect 27540 10792 27568 13262
rect 27724 13002 27752 13330
rect 27632 12974 27752 13002
rect 27632 11898 27660 12974
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27620 11892 27672 11898
rect 27724 11880 27752 12650
rect 27816 12442 27844 15200
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27804 12436 27856 12442
rect 27804 12378 27856 12384
rect 27724 11852 27844 11880
rect 27620 11834 27672 11840
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27724 11150 27752 11698
rect 27712 11144 27764 11150
rect 27712 11086 27764 11092
rect 27724 10810 27752 11086
rect 27620 10804 27672 10810
rect 27540 10764 27620 10792
rect 27620 10746 27672 10752
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27252 10736 27304 10742
rect 27252 10678 27304 10684
rect 27264 10470 27292 10678
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27264 10266 27292 10406
rect 27356 10266 27384 10542
rect 27632 10418 27660 10746
rect 27816 10713 27844 11852
rect 27802 10704 27858 10713
rect 27802 10639 27858 10648
rect 27632 10390 27844 10418
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27724 9042 27752 9318
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27066 8392 27122 8401
rect 27066 8327 27068 8336
rect 27120 8327 27122 8336
rect 27068 8298 27120 8304
rect 27264 8090 27292 8434
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 27080 4826 27108 6734
rect 27632 6390 27660 8978
rect 27710 8528 27766 8537
rect 27710 8463 27712 8472
rect 27764 8463 27766 8472
rect 27712 8434 27764 8440
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27816 4826 27844 10390
rect 27908 7818 27936 13670
rect 28092 13530 28120 15286
rect 28354 15200 28410 15286
rect 28906 15200 28962 16000
rect 29458 15200 29514 16000
rect 30010 15314 30066 16000
rect 29840 15286 30066 15314
rect 28264 13796 28316 13802
rect 28264 13738 28316 13744
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 28276 13326 28304 13738
rect 28920 13530 28948 15200
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29276 13456 29328 13462
rect 29276 13398 29328 13404
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 27986 13152 28042 13161
rect 27986 13087 28042 13096
rect 28000 11898 28028 13087
rect 28816 12912 28868 12918
rect 28816 12854 28868 12860
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 28184 11354 28212 12174
rect 28172 11348 28224 11354
rect 28172 11290 28224 11296
rect 28368 10674 28396 12174
rect 28540 12164 28592 12170
rect 28540 12106 28592 12112
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28552 8634 28580 12106
rect 28828 11762 28856 12854
rect 29012 12850 29040 13262
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 29012 11694 29040 12786
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 29196 11830 29224 12038
rect 29184 11824 29236 11830
rect 29184 11766 29236 11772
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 28906 11112 28962 11121
rect 28906 11047 28962 11056
rect 28632 9648 28684 9654
rect 28632 9590 28684 9596
rect 28644 9489 28672 9590
rect 28630 9480 28686 9489
rect 28630 9415 28686 9424
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28172 8424 28224 8430
rect 28170 8392 28172 8401
rect 28224 8392 28226 8401
rect 28170 8327 28226 8336
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 28920 5914 28948 11047
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 29104 10810 29132 10950
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 29012 5710 29040 9862
rect 29104 9722 29132 10746
rect 29288 9926 29316 13398
rect 29472 12442 29500 15200
rect 29734 12744 29790 12753
rect 29734 12679 29736 12688
rect 29788 12679 29790 12688
rect 29736 12650 29788 12656
rect 29840 12646 29868 15286
rect 30010 15200 30066 15286
rect 30562 15200 30618 16000
rect 31114 15200 31170 16000
rect 31666 15200 31722 16000
rect 32218 15314 32274 16000
rect 32218 15286 32536 15314
rect 32218 15200 32274 15286
rect 30576 13530 30604 15200
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 30116 13297 30144 13330
rect 30102 13288 30158 13297
rect 30102 13223 30158 13232
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 29828 12640 29880 12646
rect 29828 12582 29880 12588
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 30484 11830 30512 13194
rect 30654 12880 30710 12889
rect 30654 12815 30710 12824
rect 30668 12442 30696 12815
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 29552 11824 29604 11830
rect 29552 11766 29604 11772
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 29564 11218 29592 11766
rect 30196 11756 30248 11762
rect 29748 11716 30196 11744
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 29656 11150 29684 11630
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29564 10062 29592 10610
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 29472 9722 29500 9998
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29104 8974 29132 9454
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29104 8566 29132 8910
rect 29564 8634 29592 9998
rect 29748 9110 29776 11716
rect 30196 11698 30248 11704
rect 30668 11626 30696 12038
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 30656 11620 30708 11626
rect 30656 11562 30708 11568
rect 30748 11552 30800 11558
rect 30748 11494 30800 11500
rect 30760 11286 30788 11494
rect 30748 11280 30800 11286
rect 30748 11222 30800 11228
rect 29920 11076 29972 11082
rect 29972 11036 30052 11064
rect 29920 11018 29972 11024
rect 30024 10606 30052 11036
rect 30378 10976 30434 10985
rect 30378 10911 30434 10920
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30116 10674 30144 10746
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30024 9382 30052 10542
rect 30208 10198 30236 10746
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29656 8430 29684 8570
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 29366 6216 29422 6225
rect 29366 6151 29368 6160
rect 29420 6151 29422 6160
rect 29368 6122 29420 6128
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 27068 4820 27120 4826
rect 27068 4762 27120 4768
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 30116 4622 30144 9862
rect 30392 7002 30420 10911
rect 30852 10266 30880 11630
rect 30944 11354 30972 12038
rect 31128 11898 31156 15200
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 31404 12730 31432 12922
rect 31404 12702 31524 12730
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31300 12436 31352 12442
rect 31300 12378 31352 12384
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 31116 11076 31168 11082
rect 31116 11018 31168 11024
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30484 8498 30512 8910
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30576 7750 30604 8366
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30576 7478 30604 7686
rect 30564 7472 30616 7478
rect 30564 7414 30616 7420
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30208 6322 30236 6802
rect 30668 6730 30696 9590
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30564 6724 30616 6730
rect 30564 6666 30616 6672
rect 30656 6724 30708 6730
rect 30656 6666 30708 6672
rect 30196 6316 30248 6322
rect 30248 6276 30328 6304
rect 30196 6258 30248 6264
rect 30300 5166 30328 6276
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30392 5710 30420 5850
rect 30576 5846 30604 6666
rect 30472 5840 30524 5846
rect 30472 5782 30524 5788
rect 30564 5840 30616 5846
rect 30564 5782 30616 5788
rect 30484 5710 30512 5782
rect 30380 5704 30432 5710
rect 30378 5672 30380 5681
rect 30472 5704 30524 5710
rect 30432 5672 30434 5681
rect 30472 5646 30524 5652
rect 30378 5607 30434 5616
rect 30392 5574 30420 5607
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26792 3120 26844 3126
rect 26976 3120 27028 3126
rect 26844 3080 26976 3108
rect 26792 3062 26844 3068
rect 26976 3062 27028 3068
rect 30300 2990 30328 5102
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30392 4758 30420 4966
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 30484 4010 30512 5170
rect 30760 4826 30788 9522
rect 30852 8482 30880 10202
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 31036 8566 31064 9454
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 30840 8476 30892 8482
rect 30840 8418 30892 8424
rect 31036 8090 31064 8502
rect 31128 8430 31156 11018
rect 31208 11008 31260 11014
rect 31208 10950 31260 10956
rect 31220 10606 31248 10950
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 31312 10554 31340 12378
rect 31404 11354 31432 12582
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31496 11014 31524 12702
rect 31680 12442 31708 15200
rect 31758 13288 31814 13297
rect 31758 13223 31814 13232
rect 31772 12918 31800 13223
rect 32508 12986 32536 15286
rect 32770 15200 32826 16000
rect 33322 15314 33378 16000
rect 33322 15286 33548 15314
rect 33322 15200 33378 15286
rect 32784 13530 32812 15200
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32588 13320 32640 13326
rect 32588 13262 32640 13268
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 31760 12912 31812 12918
rect 31760 12854 31812 12860
rect 32036 12776 32088 12782
rect 32036 12718 32088 12724
rect 31668 12436 31720 12442
rect 31668 12378 31720 12384
rect 32048 12306 32076 12718
rect 32036 12300 32088 12306
rect 32036 12242 32088 12248
rect 32048 11762 32076 12242
rect 32324 11898 32352 12922
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 32036 11756 32088 11762
rect 32036 11698 32088 11704
rect 31680 11150 31708 11698
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 31772 11150 31800 11494
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31760 11144 31812 11150
rect 31812 11104 31892 11132
rect 31760 11086 31812 11092
rect 31484 11008 31536 11014
rect 31484 10950 31536 10956
rect 31312 10526 31432 10554
rect 31300 10464 31352 10470
rect 31300 10406 31352 10412
rect 31312 10062 31340 10406
rect 31300 10056 31352 10062
rect 31300 9998 31352 10004
rect 31312 9722 31340 9998
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 31404 8294 31432 10526
rect 31576 9988 31628 9994
rect 31576 9930 31628 9936
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31588 8090 31616 9930
rect 31680 9722 31708 11086
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 31680 9042 31708 9658
rect 31668 9036 31720 9042
rect 31668 8978 31720 8984
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 30840 6112 30892 6118
rect 30840 6054 30892 6060
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 30564 4684 30616 4690
rect 30564 4626 30616 4632
rect 30576 4214 30604 4626
rect 30564 4208 30616 4214
rect 30564 4150 30616 4156
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 30472 4004 30524 4010
rect 30472 3946 30524 3952
rect 30576 3738 30604 4014
rect 30852 4010 30880 6054
rect 31036 4690 31064 7414
rect 31760 5160 31812 5166
rect 31760 5102 31812 5108
rect 31024 4684 31076 4690
rect 31024 4626 31076 4632
rect 30840 4004 30892 4010
rect 30840 3946 30892 3952
rect 30564 3732 30616 3738
rect 30564 3674 30616 3680
rect 30576 3398 30604 3674
rect 30564 3392 30616 3398
rect 30564 3334 30616 3340
rect 31036 3058 31064 4626
rect 31772 3942 31800 5102
rect 31864 4078 31892 11104
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32048 9761 32076 9862
rect 32034 9752 32090 9761
rect 32034 9687 32090 9696
rect 32048 9654 32076 9687
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32036 6860 32088 6866
rect 32036 6802 32088 6808
rect 32048 5846 32076 6802
rect 32416 6322 32444 8842
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32508 7750 32536 7958
rect 32496 7744 32548 7750
rect 32496 7686 32548 7692
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 32036 5840 32088 5846
rect 32036 5782 32088 5788
rect 32324 5302 32352 5850
rect 32312 5296 32364 5302
rect 32312 5238 32364 5244
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31760 3936 31812 3942
rect 31760 3878 31812 3884
rect 31128 3602 31156 3878
rect 32600 3670 32628 13262
rect 33520 12986 33548 15286
rect 33874 15200 33930 16000
rect 34426 15200 34482 16000
rect 34978 15314 35034 16000
rect 34978 15286 35204 15314
rect 34978 15200 35034 15286
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33704 12102 33732 12786
rect 33888 12442 33916 15200
rect 34440 13530 34468 15200
rect 34428 13524 34480 13530
rect 34428 13466 34480 13472
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34060 13252 34112 13258
rect 34060 13194 34112 13200
rect 34428 13252 34480 13258
rect 34428 13194 34480 13200
rect 33876 12436 33928 12442
rect 33876 12378 33928 12384
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 32864 11892 32916 11898
rect 32864 11834 32916 11840
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32588 3664 32640 3670
rect 32588 3606 32640 3612
rect 31116 3596 31168 3602
rect 31116 3538 31168 3544
rect 32784 3194 32812 9998
rect 32876 8974 32904 11834
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33600 11212 33652 11218
rect 33600 11154 33652 11160
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33508 11008 33560 11014
rect 33508 10950 33560 10956
rect 33336 10810 33364 10950
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33244 10198 33272 10746
rect 33520 10742 33548 10950
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33612 10606 33640 11154
rect 33784 11008 33836 11014
rect 33784 10950 33836 10956
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 33232 10192 33284 10198
rect 33232 10134 33284 10140
rect 33612 9926 33640 10542
rect 33796 10470 33824 10950
rect 33888 10674 33916 11494
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 33784 10464 33836 10470
rect 33784 10406 33836 10412
rect 33600 9920 33652 9926
rect 33600 9862 33652 9868
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32968 8294 32996 8910
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 32864 7812 32916 7818
rect 32864 7754 32916 7760
rect 32876 7546 32904 7754
rect 32968 7750 32996 8230
rect 32956 7744 33008 7750
rect 32956 7686 33008 7692
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 32876 3466 32904 3878
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32968 3194 32996 7686
rect 33060 5574 33088 9318
rect 33232 9036 33284 9042
rect 33232 8978 33284 8984
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 33152 7342 33180 8434
rect 33244 8022 33272 8978
rect 33336 8634 33364 9522
rect 33612 9042 33640 9862
rect 33888 9518 33916 10610
rect 33876 9512 33928 9518
rect 33704 9472 33876 9500
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33704 8906 33732 9472
rect 33876 9454 33928 9460
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 33324 8628 33376 8634
rect 33324 8570 33376 8576
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 33244 6866 33272 7958
rect 33612 7886 33640 8774
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33796 7478 33824 7822
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 33232 6860 33284 6866
rect 33232 6802 33284 6808
rect 33508 6860 33560 6866
rect 33508 6802 33560 6808
rect 33520 6118 33548 6802
rect 33796 6254 33824 7414
rect 33888 6746 33916 9318
rect 33980 7750 34008 12038
rect 34072 11762 34100 13194
rect 34152 12912 34204 12918
rect 34152 12854 34204 12860
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 34072 11150 34100 11698
rect 34060 11144 34112 11150
rect 34060 11086 34112 11092
rect 34164 8838 34192 12854
rect 34440 12646 34468 13194
rect 34428 12640 34480 12646
rect 34428 12582 34480 12588
rect 34336 12164 34388 12170
rect 34336 12106 34388 12112
rect 34244 11552 34296 11558
rect 34244 11494 34296 11500
rect 34256 9654 34284 11494
rect 34348 11218 34376 12106
rect 34808 11665 34836 13262
rect 35176 12442 35204 15286
rect 35530 15200 35586 16000
rect 36082 15200 36138 16000
rect 36634 15200 36690 16000
rect 37186 15200 37242 16000
rect 37738 15200 37794 16000
rect 38290 15200 38346 16000
rect 38842 15200 38898 16000
rect 39394 15200 39450 16000
rect 39946 15200 40002 16000
rect 40498 15314 40554 16000
rect 40498 15286 40816 15314
rect 40498 15200 40554 15286
rect 35544 13530 35572 15200
rect 35532 13524 35584 13530
rect 35532 13466 35584 13472
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 35452 12918 35480 13126
rect 35440 12912 35492 12918
rect 35440 12854 35492 12860
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 35164 12436 35216 12442
rect 35164 12378 35216 12384
rect 35360 12238 35388 12718
rect 36096 12442 36124 15200
rect 36268 13796 36320 13802
rect 36268 13738 36320 13744
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 36188 13326 36216 13670
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36280 12646 36308 13738
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 36556 12986 36584 13126
rect 36648 12986 36676 15200
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 36636 12980 36688 12986
rect 36636 12922 36688 12928
rect 36728 12844 36780 12850
rect 36728 12786 36780 12792
rect 36268 12640 36320 12646
rect 36268 12582 36320 12588
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 36176 12232 36228 12238
rect 36176 12174 36228 12180
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 34888 12096 34940 12102
rect 34888 12038 34940 12044
rect 34794 11656 34850 11665
rect 34794 11591 34796 11600
rect 34848 11591 34850 11600
rect 34796 11562 34848 11568
rect 34900 11286 34928 12038
rect 35900 11824 35952 11830
rect 35900 11766 35952 11772
rect 34888 11280 34940 11286
rect 34888 11222 34940 11228
rect 34336 11212 34388 11218
rect 34336 11154 34388 11160
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 34428 10600 34480 10606
rect 34426 10568 34428 10577
rect 34992 10588 35020 11086
rect 35912 11082 35940 11766
rect 36188 11354 36216 12174
rect 36372 11898 36400 12174
rect 36360 11892 36412 11898
rect 36360 11834 36412 11840
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35256 10600 35308 10606
rect 34480 10568 34482 10577
rect 34992 10560 35256 10588
rect 35256 10542 35308 10548
rect 34426 10503 34482 10512
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 34244 9648 34296 9654
rect 34244 9590 34296 9596
rect 34532 9586 34560 9930
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 34520 9580 34572 9586
rect 34520 9522 34572 9528
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34060 7812 34112 7818
rect 34060 7754 34112 7760
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33980 6934 34008 7346
rect 33968 6928 34020 6934
rect 33968 6870 34020 6876
rect 33968 6792 34020 6798
rect 33888 6740 33968 6746
rect 33888 6734 34020 6740
rect 33888 6718 34008 6734
rect 33784 6248 33836 6254
rect 33784 6190 33836 6196
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 33796 5914 33824 6190
rect 33980 6186 34008 6718
rect 33968 6180 34020 6186
rect 33968 6122 34020 6128
rect 33784 5908 33836 5914
rect 33784 5850 33836 5856
rect 33048 5568 33100 5574
rect 33048 5510 33100 5516
rect 32772 3188 32824 3194
rect 32772 3130 32824 3136
rect 32956 3188 33008 3194
rect 32956 3130 33008 3136
rect 33060 3058 33088 5510
rect 33796 5302 33824 5850
rect 33968 5840 34020 5846
rect 33968 5782 34020 5788
rect 33980 5642 34008 5782
rect 33968 5636 34020 5642
rect 33968 5578 34020 5584
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 34072 5098 34100 7754
rect 34256 7410 34284 8570
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34428 5704 34480 5710
rect 34428 5646 34480 5652
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 34348 5166 34376 5578
rect 34336 5160 34388 5166
rect 34336 5102 34388 5108
rect 34060 5092 34112 5098
rect 34060 5034 34112 5040
rect 34348 3534 34376 5102
rect 34440 4010 34468 5646
rect 34532 5370 34560 9522
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 34900 7002 34928 7346
rect 34888 6996 34940 7002
rect 34888 6938 34940 6944
rect 34992 6118 35020 9862
rect 35268 8634 35296 10542
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 35268 8498 35296 8570
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 35360 7886 35388 9998
rect 35912 9926 35940 9998
rect 35900 9920 35952 9926
rect 35900 9862 35952 9868
rect 35912 9722 35940 9862
rect 35900 9716 35952 9722
rect 35900 9658 35952 9664
rect 35912 8634 35940 9658
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35912 8090 35940 8570
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35348 7200 35400 7206
rect 35348 7142 35400 7148
rect 34980 6112 35032 6118
rect 34980 6054 35032 6060
rect 35360 5370 35388 7142
rect 34520 5364 34572 5370
rect 34520 5306 34572 5312
rect 35348 5364 35400 5370
rect 35348 5306 35400 5312
rect 36004 5234 36032 11018
rect 36452 10464 36504 10470
rect 36452 10406 36504 10412
rect 36268 10192 36320 10198
rect 36268 10134 36320 10140
rect 36280 6746 36308 10134
rect 36464 7410 36492 10406
rect 36556 8498 36584 11494
rect 36740 11354 36768 12786
rect 37200 12442 37228 15200
rect 37752 12986 37780 15200
rect 37832 13184 37884 13190
rect 37832 13126 37884 13132
rect 37740 12980 37792 12986
rect 37740 12922 37792 12928
rect 37844 12850 37872 13126
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 38304 12442 38332 15200
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 38384 12708 38436 12714
rect 38384 12650 38436 12656
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 38292 12436 38344 12442
rect 38292 12378 38344 12384
rect 38108 12368 38160 12374
rect 38108 12310 38160 12316
rect 38200 12368 38252 12374
rect 38200 12310 38252 12316
rect 38120 12170 38148 12310
rect 38212 12238 38240 12310
rect 38396 12238 38424 12650
rect 38764 12434 38792 13262
rect 38856 12986 38884 15200
rect 39408 13530 39436 15200
rect 39396 13524 39448 13530
rect 39396 13466 39448 13472
rect 39856 13524 39908 13530
rect 39856 13466 39908 13472
rect 39488 13320 39540 13326
rect 39488 13262 39540 13268
rect 38844 12980 38896 12986
rect 38844 12922 38896 12928
rect 38764 12406 38884 12434
rect 38200 12232 38252 12238
rect 38200 12174 38252 12180
rect 38384 12232 38436 12238
rect 38384 12174 38436 12180
rect 37648 12164 37700 12170
rect 37648 12106 37700 12112
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 37660 11898 37688 12106
rect 37648 11892 37700 11898
rect 37648 11834 37700 11840
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 36728 11348 36780 11354
rect 36728 11290 36780 11296
rect 36636 9988 36688 9994
rect 36636 9930 36688 9936
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36544 8356 36596 8362
rect 36544 8298 36596 8304
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36556 6798 36584 8298
rect 36648 8090 36676 9930
rect 37200 9761 37228 11630
rect 37660 11132 37688 11834
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 11354 37872 11494
rect 37832 11348 37884 11354
rect 37832 11290 37884 11296
rect 38568 11280 38620 11286
rect 38568 11222 38620 11228
rect 37740 11144 37792 11150
rect 37660 11104 37740 11132
rect 37556 11076 37608 11082
rect 37556 11018 37608 11024
rect 37186 9752 37242 9761
rect 36728 9716 36780 9722
rect 37186 9687 37242 9696
rect 36728 9658 36780 9664
rect 36740 9042 36768 9658
rect 36728 9036 36780 9042
rect 36728 8978 36780 8984
rect 37004 8424 37056 8430
rect 37004 8366 37056 8372
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36912 7880 36964 7886
rect 36912 7822 36964 7828
rect 36636 7812 36688 7818
rect 36636 7754 36688 7760
rect 36544 6792 36596 6798
rect 36280 6718 36492 6746
rect 36544 6734 36596 6740
rect 36464 6662 36492 6718
rect 36360 6656 36412 6662
rect 36360 6598 36412 6604
rect 36452 6656 36504 6662
rect 36452 6598 36504 6604
rect 36372 6390 36400 6598
rect 36360 6384 36412 6390
rect 36360 6326 36412 6332
rect 36648 5234 36676 7754
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36636 5228 36688 5234
rect 36636 5170 36688 5176
rect 34428 4004 34480 4010
rect 34428 3946 34480 3952
rect 36924 3738 36952 7822
rect 37016 6798 37044 8366
rect 37200 7342 37228 9687
rect 37568 9450 37596 11018
rect 37660 10810 37688 11104
rect 37740 11086 37792 11092
rect 37832 11008 37884 11014
rect 37832 10950 37884 10956
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 37556 9444 37608 9450
rect 37556 9386 37608 9392
rect 37280 8900 37332 8906
rect 37280 8842 37332 8848
rect 37292 8090 37320 8842
rect 37648 8560 37700 8566
rect 37648 8502 37700 8508
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37556 7948 37608 7954
rect 37556 7890 37608 7896
rect 37188 7336 37240 7342
rect 37188 7278 37240 7284
rect 37200 6934 37228 7278
rect 37188 6928 37240 6934
rect 37188 6870 37240 6876
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 37200 5642 37228 6870
rect 37568 6458 37596 7890
rect 37660 7002 37688 8502
rect 37844 8498 37872 10950
rect 38580 10130 38608 11222
rect 38568 10124 38620 10130
rect 38568 10066 38620 10072
rect 38580 10010 38608 10066
rect 38488 9982 38608 10010
rect 38016 8832 38068 8838
rect 38016 8774 38068 8780
rect 38028 8498 38056 8774
rect 38488 8566 38516 9982
rect 38580 9846 38792 9874
rect 38580 9654 38608 9846
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 38568 9648 38620 9654
rect 38568 9590 38620 9596
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38476 8560 38528 8566
rect 38476 8502 38528 8508
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 37844 7954 37872 8434
rect 38580 8090 38608 9318
rect 38672 9178 38700 9658
rect 38764 9382 38792 9846
rect 38752 9376 38804 9382
rect 38752 9318 38804 9324
rect 38660 9172 38712 9178
rect 38660 9114 38712 9120
rect 38672 8498 38700 9114
rect 38660 8492 38712 8498
rect 38660 8434 38712 8440
rect 38568 8084 38620 8090
rect 38568 8026 38620 8032
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 37844 7410 37872 7890
rect 38568 7540 38620 7546
rect 38672 7528 38700 8434
rect 38620 7500 38700 7528
rect 38568 7482 38620 7488
rect 37832 7404 37884 7410
rect 37832 7346 37884 7352
rect 37844 7018 37872 7346
rect 38476 7336 38528 7342
rect 38476 7278 38528 7284
rect 37648 6996 37700 7002
rect 37648 6938 37700 6944
rect 37752 6990 37872 7018
rect 37464 6452 37516 6458
rect 37464 6394 37516 6400
rect 37556 6452 37608 6458
rect 37556 6394 37608 6400
rect 37476 5846 37504 6394
rect 37464 5840 37516 5846
rect 37464 5782 37516 5788
rect 37188 5636 37240 5642
rect 37188 5578 37240 5584
rect 37188 4072 37240 4078
rect 37188 4014 37240 4020
rect 37200 3738 37228 4014
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 37188 3732 37240 3738
rect 37188 3674 37240 3680
rect 37200 3534 37228 3674
rect 37752 3670 37780 6990
rect 37832 6860 37884 6866
rect 37832 6802 37884 6808
rect 37844 5710 37872 6802
rect 38384 6724 38436 6730
rect 38384 6666 38436 6672
rect 38396 6458 38424 6666
rect 38384 6452 38436 6458
rect 38384 6394 38436 6400
rect 38488 6322 38516 7278
rect 38476 6316 38528 6322
rect 38476 6258 38528 6264
rect 38660 6316 38712 6322
rect 38660 6258 38712 6264
rect 38488 6202 38516 6258
rect 38016 6180 38068 6186
rect 38488 6174 38608 6202
rect 38016 6122 38068 6128
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 38028 5642 38056 6122
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 38580 5574 38608 6174
rect 38672 5914 38700 6258
rect 38660 5908 38712 5914
rect 38660 5850 38712 5856
rect 38568 5568 38620 5574
rect 38568 5510 38620 5516
rect 38580 5234 38608 5510
rect 38568 5228 38620 5234
rect 38568 5170 38620 5176
rect 38580 4622 38608 5170
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 37372 3664 37424 3670
rect 37372 3606 37424 3612
rect 37740 3664 37792 3670
rect 37740 3606 37792 3612
rect 37384 3534 37412 3606
rect 34336 3528 34388 3534
rect 34336 3470 34388 3476
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 37924 3392 37976 3398
rect 37924 3334 37976 3340
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 25976 2746 26096 2774
rect 25976 2582 26004 2746
rect 25964 2576 26016 2582
rect 25964 2518 26016 2524
rect 33796 2514 33824 3334
rect 37936 3126 37964 3334
rect 37924 3120 37976 3126
rect 37924 3062 37976 3068
rect 38856 2854 38884 12406
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 39132 11082 39160 11698
rect 39224 11558 39252 12174
rect 39500 11898 39528 13262
rect 39868 12782 39896 13466
rect 39856 12776 39908 12782
rect 39856 12718 39908 12724
rect 39960 12442 39988 15200
rect 40316 13320 40368 13326
rect 40316 13262 40368 13268
rect 40132 13184 40184 13190
rect 40132 13126 40184 13132
rect 39948 12436 40000 12442
rect 39948 12378 40000 12384
rect 39856 12164 39908 12170
rect 39856 12106 39908 12112
rect 39304 11892 39356 11898
rect 39304 11834 39356 11840
rect 39488 11892 39540 11898
rect 39488 11834 39540 11840
rect 39316 11626 39344 11834
rect 39304 11620 39356 11626
rect 39304 11562 39356 11568
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39120 11076 39172 11082
rect 39120 11018 39172 11024
rect 39396 10464 39448 10470
rect 39396 10406 39448 10412
rect 39408 10266 39436 10406
rect 39396 10260 39448 10266
rect 39396 10202 39448 10208
rect 39396 9920 39448 9926
rect 39396 9862 39448 9868
rect 39408 9654 39436 9862
rect 39396 9648 39448 9654
rect 39396 9590 39448 9596
rect 39396 9172 39448 9178
rect 39396 9114 39448 9120
rect 39408 8566 39436 9114
rect 39762 8936 39818 8945
rect 39762 8871 39818 8880
rect 39776 8838 39804 8871
rect 39764 8832 39816 8838
rect 39764 8774 39816 8780
rect 38936 8560 38988 8566
rect 38936 8502 38988 8508
rect 39396 8560 39448 8566
rect 39396 8502 39448 8508
rect 38948 8022 38976 8502
rect 39304 8288 39356 8294
rect 39304 8230 39356 8236
rect 38936 8016 38988 8022
rect 38936 7958 38988 7964
rect 39120 8016 39172 8022
rect 39120 7958 39172 7964
rect 39132 7818 39160 7958
rect 39316 7886 39344 8230
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39120 7812 39172 7818
rect 39120 7754 39172 7760
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39868 2802 39896 12106
rect 40040 11824 40092 11830
rect 40040 11766 40092 11772
rect 40144 11778 40172 13126
rect 40224 12844 40276 12850
rect 40224 12786 40276 12792
rect 40236 12345 40264 12786
rect 40222 12336 40278 12345
rect 40222 12271 40278 12280
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 40236 11898 40264 12174
rect 40328 12170 40356 13262
rect 40394 13084 40702 13093
rect 40394 13082 40400 13084
rect 40456 13082 40480 13084
rect 40536 13082 40560 13084
rect 40616 13082 40640 13084
rect 40696 13082 40702 13084
rect 40456 13030 40458 13082
rect 40638 13030 40640 13082
rect 40394 13028 40400 13030
rect 40456 13028 40480 13030
rect 40536 13028 40560 13030
rect 40616 13028 40640 13030
rect 40696 13028 40702 13030
rect 40394 13019 40702 13028
rect 40316 12164 40368 12170
rect 40316 12106 40368 12112
rect 40224 11892 40276 11898
rect 40224 11834 40276 11840
rect 40052 11506 40080 11766
rect 40144 11750 40264 11778
rect 39960 11478 40080 11506
rect 39960 9364 39988 11478
rect 40040 11348 40092 11354
rect 40040 11290 40092 11296
rect 40052 10810 40080 11290
rect 40236 11150 40264 11750
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 40132 11076 40184 11082
rect 40132 11018 40184 11024
rect 40040 10804 40092 10810
rect 40040 10746 40092 10752
rect 40040 10532 40092 10538
rect 40040 10474 40092 10480
rect 40052 9518 40080 10474
rect 40144 10470 40172 11018
rect 40224 10668 40276 10674
rect 40224 10610 40276 10616
rect 40132 10464 40184 10470
rect 40132 10406 40184 10412
rect 40236 9654 40264 10610
rect 40224 9648 40276 9654
rect 40224 9590 40276 9596
rect 40040 9512 40092 9518
rect 40040 9454 40092 9460
rect 40224 9376 40276 9382
rect 39960 9336 40080 9364
rect 40052 8838 40080 9336
rect 40224 9318 40276 9324
rect 40236 9110 40264 9318
rect 40224 9104 40276 9110
rect 40224 9046 40276 9052
rect 40040 8832 40092 8838
rect 40040 8774 40092 8780
rect 40328 7546 40356 12106
rect 40394 11996 40702 12005
rect 40394 11994 40400 11996
rect 40456 11994 40480 11996
rect 40536 11994 40560 11996
rect 40616 11994 40640 11996
rect 40696 11994 40702 11996
rect 40456 11942 40458 11994
rect 40638 11942 40640 11994
rect 40394 11940 40400 11942
rect 40456 11940 40480 11942
rect 40536 11940 40560 11942
rect 40616 11940 40640 11942
rect 40696 11940 40702 11942
rect 40394 11931 40702 11940
rect 40788 11354 40816 15286
rect 41050 15200 41106 16000
rect 41602 15200 41658 16000
rect 42154 15314 42210 16000
rect 42706 15314 42762 16000
rect 41800 15286 42210 15314
rect 41064 13394 41092 15200
rect 41328 13796 41380 13802
rect 41328 13738 41380 13744
rect 41420 13796 41472 13802
rect 41420 13738 41472 13744
rect 41052 13388 41104 13394
rect 41052 13330 41104 13336
rect 41340 13326 41368 13738
rect 41144 13320 41196 13326
rect 41144 13262 41196 13268
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 41156 12434 41184 13262
rect 41156 12406 41276 12434
rect 40866 12336 40922 12345
rect 41248 12306 41276 12406
rect 40866 12271 40922 12280
rect 41236 12300 41288 12306
rect 40776 11348 40828 11354
rect 40776 11290 40828 11296
rect 40776 11008 40828 11014
rect 40776 10950 40828 10956
rect 40394 10908 40702 10917
rect 40394 10906 40400 10908
rect 40456 10906 40480 10908
rect 40536 10906 40560 10908
rect 40616 10906 40640 10908
rect 40696 10906 40702 10908
rect 40456 10854 40458 10906
rect 40638 10854 40640 10906
rect 40394 10852 40400 10854
rect 40456 10852 40480 10854
rect 40536 10852 40560 10854
rect 40616 10852 40640 10854
rect 40696 10852 40702 10854
rect 40394 10843 40702 10852
rect 40408 10804 40460 10810
rect 40408 10746 40460 10752
rect 40420 10266 40448 10746
rect 40788 10266 40816 10950
rect 40408 10260 40460 10266
rect 40408 10202 40460 10208
rect 40776 10260 40828 10266
rect 40776 10202 40828 10208
rect 40394 9820 40702 9829
rect 40394 9818 40400 9820
rect 40456 9818 40480 9820
rect 40536 9818 40560 9820
rect 40616 9818 40640 9820
rect 40696 9818 40702 9820
rect 40456 9766 40458 9818
rect 40638 9766 40640 9818
rect 40394 9764 40400 9766
rect 40456 9764 40480 9766
rect 40536 9764 40560 9766
rect 40616 9764 40640 9766
rect 40696 9764 40702 9766
rect 40394 9755 40702 9764
rect 40394 8732 40702 8741
rect 40394 8730 40400 8732
rect 40456 8730 40480 8732
rect 40536 8730 40560 8732
rect 40616 8730 40640 8732
rect 40696 8730 40702 8732
rect 40456 8678 40458 8730
rect 40638 8678 40640 8730
rect 40394 8676 40400 8678
rect 40456 8676 40480 8678
rect 40536 8676 40560 8678
rect 40616 8676 40640 8678
rect 40696 8676 40702 8678
rect 40394 8667 40702 8676
rect 40788 8362 40816 10202
rect 40776 8356 40828 8362
rect 40776 8298 40828 8304
rect 40776 7880 40828 7886
rect 40776 7822 40828 7828
rect 40394 7644 40702 7653
rect 40394 7642 40400 7644
rect 40456 7642 40480 7644
rect 40536 7642 40560 7644
rect 40616 7642 40640 7644
rect 40696 7642 40702 7644
rect 40456 7590 40458 7642
rect 40638 7590 40640 7642
rect 40394 7588 40400 7590
rect 40456 7588 40480 7590
rect 40536 7588 40560 7590
rect 40616 7588 40640 7590
rect 40696 7588 40702 7590
rect 40394 7579 40702 7588
rect 40316 7540 40368 7546
rect 40316 7482 40368 7488
rect 40788 7410 40816 7822
rect 40776 7404 40828 7410
rect 40776 7346 40828 7352
rect 40224 6996 40276 7002
rect 40224 6938 40276 6944
rect 40236 6322 40264 6938
rect 40394 6556 40702 6565
rect 40394 6554 40400 6556
rect 40456 6554 40480 6556
rect 40536 6554 40560 6556
rect 40616 6554 40640 6556
rect 40696 6554 40702 6556
rect 40456 6502 40458 6554
rect 40638 6502 40640 6554
rect 40394 6500 40400 6502
rect 40456 6500 40480 6502
rect 40536 6500 40560 6502
rect 40616 6500 40640 6502
rect 40696 6500 40702 6502
rect 40394 6491 40702 6500
rect 40880 6390 40908 12271
rect 41236 12242 41288 12248
rect 41248 11218 41276 12242
rect 41432 12238 41460 13738
rect 41512 13320 41564 13326
rect 41512 13262 41564 13268
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 41524 11762 41552 13262
rect 41616 12986 41644 15200
rect 41604 12980 41656 12986
rect 41604 12922 41656 12928
rect 41696 12912 41748 12918
rect 41696 12854 41748 12860
rect 41708 12753 41736 12854
rect 41694 12744 41750 12753
rect 41616 12702 41694 12730
rect 41512 11756 41564 11762
rect 41512 11698 41564 11704
rect 41328 11620 41380 11626
rect 41328 11562 41380 11568
rect 41340 11218 41368 11562
rect 41236 11212 41288 11218
rect 41236 11154 41288 11160
rect 41328 11212 41380 11218
rect 41328 11154 41380 11160
rect 41420 11144 41472 11150
rect 41420 11086 41472 11092
rect 41144 10668 41196 10674
rect 41144 10610 41196 10616
rect 41328 10668 41380 10674
rect 41328 10610 41380 10616
rect 40960 10464 41012 10470
rect 40960 10406 41012 10412
rect 40972 9654 41000 10406
rect 41052 10260 41104 10266
rect 41052 10202 41104 10208
rect 41064 10062 41092 10202
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 40960 9648 41012 9654
rect 40960 9590 41012 9596
rect 41052 8968 41104 8974
rect 41052 8910 41104 8916
rect 40960 8900 41012 8906
rect 40960 8842 41012 8848
rect 40868 6384 40920 6390
rect 40868 6326 40920 6332
rect 40224 6316 40276 6322
rect 40224 6258 40276 6264
rect 40972 6254 41000 8842
rect 41064 8838 41092 8910
rect 41052 8832 41104 8838
rect 41052 8774 41104 8780
rect 41052 8628 41104 8634
rect 41052 8570 41104 8576
rect 41064 8537 41092 8570
rect 41050 8528 41106 8537
rect 41156 8498 41184 10610
rect 41236 10532 41288 10538
rect 41236 10474 41288 10480
rect 41248 10198 41276 10474
rect 41236 10192 41288 10198
rect 41236 10134 41288 10140
rect 41234 9072 41290 9081
rect 41234 9007 41290 9016
rect 41050 8463 41106 8472
rect 41144 8492 41196 8498
rect 41144 8434 41196 8440
rect 41248 8362 41276 9007
rect 41236 8356 41288 8362
rect 41236 8298 41288 8304
rect 41236 7404 41288 7410
rect 41236 7346 41288 7352
rect 41248 6458 41276 7346
rect 41236 6452 41288 6458
rect 41236 6394 41288 6400
rect 40960 6248 41012 6254
rect 40960 6190 41012 6196
rect 41236 6180 41288 6186
rect 41236 6122 41288 6128
rect 41248 5710 41276 6122
rect 41236 5704 41288 5710
rect 41236 5646 41288 5652
rect 40394 5468 40702 5477
rect 40394 5466 40400 5468
rect 40456 5466 40480 5468
rect 40536 5466 40560 5468
rect 40616 5466 40640 5468
rect 40696 5466 40702 5468
rect 40456 5414 40458 5466
rect 40638 5414 40640 5466
rect 40394 5412 40400 5414
rect 40456 5412 40480 5414
rect 40536 5412 40560 5414
rect 40616 5412 40640 5414
rect 40696 5412 40702 5414
rect 40394 5403 40702 5412
rect 40394 4380 40702 4389
rect 40394 4378 40400 4380
rect 40456 4378 40480 4380
rect 40536 4378 40560 4380
rect 40616 4378 40640 4380
rect 40696 4378 40702 4380
rect 40456 4326 40458 4378
rect 40638 4326 40640 4378
rect 40394 4324 40400 4326
rect 40456 4324 40480 4326
rect 40536 4324 40560 4326
rect 40616 4324 40640 4326
rect 40696 4324 40702 4326
rect 40394 4315 40702 4324
rect 40394 3292 40702 3301
rect 40394 3290 40400 3292
rect 40456 3290 40480 3292
rect 40536 3290 40560 3292
rect 40616 3290 40640 3292
rect 40696 3290 40702 3292
rect 40456 3238 40458 3290
rect 40638 3238 40640 3290
rect 40394 3236 40400 3238
rect 40456 3236 40480 3238
rect 40536 3236 40560 3238
rect 40616 3236 40640 3238
rect 40696 3236 40702 3238
rect 40394 3227 40702 3236
rect 40316 2848 40368 2854
rect 39868 2796 40316 2802
rect 39868 2790 40368 2796
rect 39868 2774 40356 2790
rect 41340 2650 41368 10610
rect 41432 10266 41460 11086
rect 41512 11008 41564 11014
rect 41512 10950 41564 10956
rect 41524 10810 41552 10950
rect 41512 10804 41564 10810
rect 41512 10746 41564 10752
rect 41420 10260 41472 10266
rect 41420 10202 41472 10208
rect 41512 9580 41564 9586
rect 41512 9522 41564 9528
rect 41524 8906 41552 9522
rect 41616 8945 41644 12702
rect 41694 12679 41750 12688
rect 41800 12646 41828 15286
rect 42154 15200 42210 15286
rect 42444 15286 42762 15314
rect 42340 13728 42392 13734
rect 42340 13670 42392 13676
rect 41880 13320 41932 13326
rect 41880 13262 41932 13268
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41696 12436 41748 12442
rect 41696 12378 41748 12384
rect 41708 11898 41736 12378
rect 41696 11892 41748 11898
rect 41696 11834 41748 11840
rect 41708 10470 41736 11834
rect 41788 11144 41840 11150
rect 41788 11086 41840 11092
rect 41800 10606 41828 11086
rect 41788 10600 41840 10606
rect 41788 10542 41840 10548
rect 41696 10464 41748 10470
rect 41696 10406 41748 10412
rect 41708 8974 41736 10406
rect 41788 9920 41840 9926
rect 41788 9862 41840 9868
rect 41800 9586 41828 9862
rect 41788 9580 41840 9586
rect 41788 9522 41840 9528
rect 41892 9450 41920 13262
rect 42248 12912 42300 12918
rect 42248 12854 42300 12860
rect 42156 12368 42208 12374
rect 42154 12336 42156 12345
rect 42208 12336 42210 12345
rect 42154 12271 42210 12280
rect 42064 12232 42116 12238
rect 42064 12174 42116 12180
rect 41972 11756 42024 11762
rect 41972 11698 42024 11704
rect 41984 9602 42012 11698
rect 42076 11393 42104 12174
rect 42156 12096 42208 12102
rect 42156 12038 42208 12044
rect 42168 11762 42196 12038
rect 42156 11756 42208 11762
rect 42156 11698 42208 11704
rect 42062 11384 42118 11393
rect 42062 11319 42118 11328
rect 42260 11286 42288 12854
rect 42248 11280 42300 11286
rect 42248 11222 42300 11228
rect 41984 9574 42104 9602
rect 41880 9444 41932 9450
rect 41880 9386 41932 9392
rect 41696 8968 41748 8974
rect 41602 8936 41658 8945
rect 41512 8900 41564 8906
rect 41696 8910 41748 8916
rect 41602 8871 41658 8880
rect 41512 8842 41564 8848
rect 41708 8090 41736 8910
rect 41892 8906 41920 9386
rect 41972 9376 42024 9382
rect 42076 9353 42104 9574
rect 41972 9318 42024 9324
rect 42062 9344 42118 9353
rect 41880 8900 41932 8906
rect 41880 8842 41932 8848
rect 41788 8628 41840 8634
rect 41788 8570 41840 8576
rect 41800 8294 41828 8570
rect 41788 8288 41840 8294
rect 41788 8230 41840 8236
rect 41696 8084 41748 8090
rect 41696 8026 41748 8032
rect 41984 4078 42012 9318
rect 42062 9279 42118 9288
rect 42076 8362 42104 9279
rect 42064 8356 42116 8362
rect 42064 8298 42116 8304
rect 42076 7546 42104 8298
rect 42352 8294 42380 13670
rect 42444 13258 42472 15286
rect 42706 15200 42762 15286
rect 43258 15200 43314 16000
rect 43810 15314 43866 16000
rect 43364 15286 43866 15314
rect 42524 13796 42576 13802
rect 42524 13738 42576 13744
rect 43168 13796 43220 13802
rect 43168 13738 43220 13744
rect 42432 13252 42484 13258
rect 42432 13194 42484 13200
rect 42432 11552 42484 11558
rect 42432 11494 42484 11500
rect 42340 8288 42392 8294
rect 42340 8230 42392 8236
rect 42064 7540 42116 7546
rect 42064 7482 42116 7488
rect 42444 7410 42472 11494
rect 42536 11218 42564 13738
rect 42984 13524 43036 13530
rect 42984 13466 43036 13472
rect 42708 13320 42760 13326
rect 42708 13262 42760 13268
rect 42720 12850 42748 13262
rect 42800 13184 42852 13190
rect 42800 13126 42852 13132
rect 42708 12844 42760 12850
rect 42708 12786 42760 12792
rect 42708 12096 42760 12102
rect 42708 12038 42760 12044
rect 42616 11688 42668 11694
rect 42616 11630 42668 11636
rect 42628 11529 42656 11630
rect 42614 11520 42670 11529
rect 42614 11455 42670 11464
rect 42720 11286 42748 12038
rect 42812 11914 42840 13126
rect 42892 12640 42944 12646
rect 42892 12582 42944 12588
rect 42904 12102 42932 12582
rect 42892 12096 42944 12102
rect 42892 12038 42944 12044
rect 42812 11886 42932 11914
rect 42800 11756 42852 11762
rect 42800 11698 42852 11704
rect 42708 11280 42760 11286
rect 42708 11222 42760 11228
rect 42524 11212 42576 11218
rect 42524 11154 42576 11160
rect 42616 11008 42668 11014
rect 42616 10950 42668 10956
rect 42628 10810 42656 10950
rect 42616 10804 42668 10810
rect 42616 10746 42668 10752
rect 42616 10464 42668 10470
rect 42616 10406 42668 10412
rect 42628 7886 42656 10406
rect 42720 10062 42748 11222
rect 42708 10056 42760 10062
rect 42708 9998 42760 10004
rect 42812 8090 42840 11698
rect 42904 9654 42932 11886
rect 42892 9648 42944 9654
rect 42892 9590 42944 9596
rect 42996 8090 43024 13466
rect 43076 13456 43128 13462
rect 43076 13398 43128 13404
rect 43088 12866 43116 13398
rect 43180 13258 43208 13738
rect 43168 13252 43220 13258
rect 43168 13194 43220 13200
rect 43088 12838 43208 12866
rect 43074 11520 43130 11529
rect 43074 11455 43130 11464
rect 43088 9586 43116 11455
rect 43180 10146 43208 12838
rect 43272 11898 43300 15200
rect 43260 11892 43312 11898
rect 43260 11834 43312 11840
rect 43364 11370 43392 15286
rect 43810 15200 43866 15286
rect 44362 15200 44418 16000
rect 44914 15200 44970 16000
rect 45466 15314 45522 16000
rect 45112 15286 45522 15314
rect 43904 13932 43956 13938
rect 43904 13874 43956 13880
rect 43720 13252 43772 13258
rect 43720 13194 43772 13200
rect 43812 13252 43864 13258
rect 43812 13194 43864 13200
rect 43628 13184 43680 13190
rect 43628 13126 43680 13132
rect 43536 12368 43588 12374
rect 43536 12310 43588 12316
rect 43272 11354 43392 11370
rect 43260 11348 43392 11354
rect 43312 11342 43392 11348
rect 43260 11290 43312 11296
rect 43352 11076 43404 11082
rect 43352 11018 43404 11024
rect 43180 10118 43300 10146
rect 43168 10056 43220 10062
rect 43168 9998 43220 10004
rect 43076 9580 43128 9586
rect 43076 9522 43128 9528
rect 43180 9518 43208 9998
rect 43168 9512 43220 9518
rect 43168 9454 43220 9460
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 42984 8084 43036 8090
rect 42984 8026 43036 8032
rect 42616 7880 42668 7886
rect 42616 7822 42668 7828
rect 42892 7812 42944 7818
rect 42892 7754 42944 7760
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 42904 7274 42932 7754
rect 42892 7268 42944 7274
rect 42892 7210 42944 7216
rect 43088 4282 43116 9318
rect 43180 8974 43208 9454
rect 43168 8968 43220 8974
rect 43168 8910 43220 8916
rect 43180 7546 43208 8910
rect 43168 7540 43220 7546
rect 43168 7482 43220 7488
rect 43272 5914 43300 10118
rect 43260 5908 43312 5914
rect 43260 5850 43312 5856
rect 43364 5370 43392 11018
rect 43548 10062 43576 12310
rect 43640 11830 43668 13126
rect 43732 12918 43760 13194
rect 43824 12986 43852 13194
rect 43812 12980 43864 12986
rect 43812 12922 43864 12928
rect 43720 12912 43772 12918
rect 43720 12854 43772 12860
rect 43916 12374 43944 13874
rect 43994 13424 44050 13433
rect 43994 13359 44050 13368
rect 44008 12986 44036 13359
rect 43996 12980 44048 12986
rect 43996 12922 44048 12928
rect 43904 12368 43956 12374
rect 43904 12310 43956 12316
rect 44008 12306 44036 12922
rect 44272 12776 44324 12782
rect 44272 12718 44324 12724
rect 44284 12442 44312 12718
rect 44272 12436 44324 12442
rect 44272 12378 44324 12384
rect 43996 12300 44048 12306
rect 43996 12242 44048 12248
rect 44088 12096 44140 12102
rect 44088 12038 44140 12044
rect 43628 11824 43680 11830
rect 43628 11766 43680 11772
rect 43904 11824 43956 11830
rect 43904 11766 43956 11772
rect 43536 10056 43588 10062
rect 43536 9998 43588 10004
rect 43916 9382 43944 11766
rect 43904 9376 43956 9382
rect 43904 9318 43956 9324
rect 43996 8968 44048 8974
rect 43996 8910 44048 8916
rect 44008 8430 44036 8910
rect 44100 8480 44128 12038
rect 44180 11756 44232 11762
rect 44180 11698 44232 11704
rect 44192 8838 44220 11698
rect 44376 11694 44404 15200
rect 44364 11688 44416 11694
rect 44364 11630 44416 11636
rect 44928 10810 44956 15200
rect 45112 13802 45140 15286
rect 45466 15200 45522 15286
rect 46018 15200 46074 16000
rect 46570 15200 46626 16000
rect 47122 15200 47178 16000
rect 47674 15200 47730 16000
rect 48226 15200 48282 16000
rect 48778 15200 48834 16000
rect 49330 15200 49386 16000
rect 49882 15314 49938 16000
rect 49712 15286 49938 15314
rect 45100 13796 45152 13802
rect 45100 13738 45152 13744
rect 45560 13728 45612 13734
rect 45560 13670 45612 13676
rect 45572 13462 45600 13670
rect 45560 13456 45612 13462
rect 45560 13398 45612 13404
rect 45928 13320 45980 13326
rect 45928 13262 45980 13268
rect 45560 13184 45612 13190
rect 45560 13126 45612 13132
rect 45572 12782 45600 13126
rect 45560 12776 45612 12782
rect 45560 12718 45612 12724
rect 45558 12472 45614 12481
rect 45558 12407 45560 12416
rect 45612 12407 45614 12416
rect 45560 12378 45612 12384
rect 45940 12238 45968 13262
rect 45008 12232 45060 12238
rect 45468 12232 45520 12238
rect 45008 12174 45060 12180
rect 45466 12200 45468 12209
rect 45928 12232 45980 12238
rect 45520 12200 45522 12209
rect 44824 10804 44876 10810
rect 44824 10746 44876 10752
rect 44916 10804 44968 10810
rect 44916 10746 44968 10752
rect 44836 10690 44864 10746
rect 45020 10690 45048 12174
rect 45928 12174 45980 12180
rect 45466 12135 45522 12144
rect 45652 11756 45704 11762
rect 45652 11698 45704 11704
rect 45374 11384 45430 11393
rect 45374 11319 45430 11328
rect 45388 11286 45416 11319
rect 45664 11286 45692 11698
rect 45376 11280 45428 11286
rect 45376 11222 45428 11228
rect 45652 11280 45704 11286
rect 45652 11222 45704 11228
rect 45652 11144 45704 11150
rect 45652 11086 45704 11092
rect 45744 11144 45796 11150
rect 45744 11086 45796 11092
rect 45468 11076 45520 11082
rect 45468 11018 45520 11024
rect 44836 10662 45048 10690
rect 44916 10600 44968 10606
rect 44916 10542 44968 10548
rect 44456 10260 44508 10266
rect 44456 10202 44508 10208
rect 44180 8832 44232 8838
rect 44180 8774 44232 8780
rect 44180 8492 44232 8498
rect 44100 8452 44180 8480
rect 44180 8434 44232 8440
rect 43996 8424 44048 8430
rect 43996 8366 44048 8372
rect 44088 8356 44140 8362
rect 44088 8298 44140 8304
rect 43536 6792 43588 6798
rect 43536 6734 43588 6740
rect 43548 6662 43576 6734
rect 43536 6656 43588 6662
rect 43536 6598 43588 6604
rect 43548 6322 43576 6598
rect 43536 6316 43588 6322
rect 43536 6258 43588 6264
rect 43628 5840 43680 5846
rect 43628 5782 43680 5788
rect 43640 5574 43668 5782
rect 43628 5568 43680 5574
rect 43628 5510 43680 5516
rect 43352 5364 43404 5370
rect 43352 5306 43404 5312
rect 44100 4570 44128 8298
rect 44364 7200 44416 7206
rect 44364 7142 44416 7148
rect 44180 6792 44232 6798
rect 44180 6734 44232 6740
rect 44192 4758 44220 6734
rect 44376 6662 44404 7142
rect 44364 6656 44416 6662
rect 44364 6598 44416 6604
rect 44468 5914 44496 10202
rect 44928 10062 44956 10542
rect 44640 10056 44692 10062
rect 44640 9998 44692 10004
rect 44916 10056 44968 10062
rect 44916 9998 44968 10004
rect 44652 7886 44680 9998
rect 44732 9444 44784 9450
rect 44732 9386 44784 9392
rect 44744 9178 44772 9386
rect 44732 9172 44784 9178
rect 44732 9114 44784 9120
rect 44730 8528 44786 8537
rect 44730 8463 44732 8472
rect 44784 8463 44786 8472
rect 44732 8434 44784 8440
rect 44640 7880 44692 7886
rect 44640 7822 44692 7828
rect 44652 6440 44680 7822
rect 45020 6866 45048 10662
rect 45376 10668 45428 10674
rect 45112 10628 45376 10656
rect 45008 6860 45060 6866
rect 45008 6802 45060 6808
rect 45112 6798 45140 10628
rect 45376 10610 45428 10616
rect 45192 10464 45244 10470
rect 45192 10406 45244 10412
rect 45204 9722 45232 10406
rect 45192 9716 45244 9722
rect 45192 9658 45244 9664
rect 45192 9376 45244 9382
rect 45192 9318 45244 9324
rect 45100 6792 45152 6798
rect 45100 6734 45152 6740
rect 44732 6452 44784 6458
rect 44652 6412 44732 6440
rect 44456 5908 44508 5914
rect 44456 5850 44508 5856
rect 44652 5778 44680 6412
rect 44732 6394 44784 6400
rect 44640 5772 44692 5778
rect 44640 5714 44692 5720
rect 44180 4752 44232 4758
rect 44180 4694 44232 4700
rect 44008 4554 44128 4570
rect 43996 4548 44128 4554
rect 44048 4542 44128 4548
rect 43996 4490 44048 4496
rect 43076 4276 43128 4282
rect 43076 4218 43128 4224
rect 44652 4146 44680 5714
rect 45204 4978 45232 9318
rect 45480 9178 45508 11018
rect 45560 9920 45612 9926
rect 45560 9862 45612 9868
rect 45468 9172 45520 9178
rect 45468 9114 45520 9120
rect 45572 9042 45600 9862
rect 45560 9036 45612 9042
rect 45560 8978 45612 8984
rect 45376 8968 45428 8974
rect 45376 8910 45428 8916
rect 45388 8430 45416 8910
rect 45468 8900 45520 8906
rect 45468 8842 45520 8848
rect 45560 8900 45612 8906
rect 45560 8842 45612 8848
rect 45480 8634 45508 8842
rect 45468 8628 45520 8634
rect 45468 8570 45520 8576
rect 45376 8424 45428 8430
rect 45376 8366 45428 8372
rect 45388 8090 45416 8366
rect 45376 8084 45428 8090
rect 45376 8026 45428 8032
rect 45468 8084 45520 8090
rect 45468 8026 45520 8032
rect 45388 7546 45416 8026
rect 45480 7954 45508 8026
rect 45468 7948 45520 7954
rect 45468 7890 45520 7896
rect 45376 7540 45428 7546
rect 45376 7482 45428 7488
rect 45572 7478 45600 8842
rect 45664 8634 45692 11086
rect 45756 9382 45784 11086
rect 45940 10742 45968 12174
rect 46032 11558 46060 15200
rect 46112 13728 46164 13734
rect 46112 13670 46164 13676
rect 46020 11552 46072 11558
rect 46020 11494 46072 11500
rect 46124 10810 46152 13670
rect 46294 12744 46350 12753
rect 46294 12679 46350 12688
rect 46308 11150 46336 12679
rect 46388 11824 46440 11830
rect 46388 11766 46440 11772
rect 46400 11558 46428 11766
rect 46388 11552 46440 11558
rect 46388 11494 46440 11500
rect 46204 11144 46256 11150
rect 46204 11086 46256 11092
rect 46296 11144 46348 11150
rect 46296 11086 46348 11092
rect 46112 10804 46164 10810
rect 46112 10746 46164 10752
rect 45928 10736 45980 10742
rect 45928 10678 45980 10684
rect 46020 10736 46072 10742
rect 46020 10678 46072 10684
rect 46032 10266 46060 10678
rect 46020 10260 46072 10266
rect 46020 10202 46072 10208
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 45744 9376 45796 9382
rect 45744 9318 45796 9324
rect 45652 8628 45704 8634
rect 45652 8570 45704 8576
rect 45560 7472 45612 7478
rect 45560 7414 45612 7420
rect 45756 7206 45784 9318
rect 45928 8628 45980 8634
rect 45928 8570 45980 8576
rect 45836 7880 45888 7886
rect 45836 7822 45888 7828
rect 45848 7478 45876 7822
rect 45836 7472 45888 7478
rect 45836 7414 45888 7420
rect 45848 7342 45876 7414
rect 45836 7336 45888 7342
rect 45836 7278 45888 7284
rect 45744 7200 45796 7206
rect 45744 7142 45796 7148
rect 45468 6724 45520 6730
rect 45468 6666 45520 6672
rect 45376 5296 45428 5302
rect 45376 5238 45428 5244
rect 45204 4950 45324 4978
rect 45192 4820 45244 4826
rect 45192 4762 45244 4768
rect 42892 4140 42944 4146
rect 42892 4082 42944 4088
rect 44180 4140 44232 4146
rect 44180 4082 44232 4088
rect 44640 4140 44692 4146
rect 44640 4082 44692 4088
rect 41972 4072 42024 4078
rect 41972 4014 42024 4020
rect 42904 2990 42932 4082
rect 44192 3058 44220 4082
rect 45204 3670 45232 4762
rect 45296 4146 45324 4950
rect 45284 4140 45336 4146
rect 45284 4082 45336 4088
rect 45192 3664 45244 3670
rect 45192 3606 45244 3612
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 42892 2984 42944 2990
rect 42892 2926 42944 2932
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 45388 2378 45416 5238
rect 45480 4622 45508 6666
rect 45848 5778 45876 7278
rect 45940 6322 45968 8570
rect 46020 8288 46072 8294
rect 46020 8230 46072 8236
rect 46032 7886 46060 8230
rect 46020 7880 46072 7886
rect 46020 7822 46072 7828
rect 46020 6452 46072 6458
rect 46020 6394 46072 6400
rect 45928 6316 45980 6322
rect 45928 6258 45980 6264
rect 46032 6254 46060 6394
rect 46020 6248 46072 6254
rect 46020 6190 46072 6196
rect 46032 5778 46060 6190
rect 45836 5772 45888 5778
rect 45836 5714 45888 5720
rect 46020 5772 46072 5778
rect 46020 5714 46072 5720
rect 45848 5302 45876 5714
rect 45836 5296 45888 5302
rect 45836 5238 45888 5244
rect 46124 4826 46152 9998
rect 46216 8090 46244 11086
rect 46584 10266 46612 15200
rect 47136 13938 47164 15200
rect 47124 13932 47176 13938
rect 47124 13874 47176 13880
rect 46664 13796 46716 13802
rect 46664 13738 46716 13744
rect 46940 13796 46992 13802
rect 46940 13738 46992 13744
rect 46676 13462 46704 13738
rect 46664 13456 46716 13462
rect 46664 13398 46716 13404
rect 46952 12714 46980 13738
rect 47216 13320 47268 13326
rect 47216 13262 47268 13268
rect 47228 12782 47256 13262
rect 47216 12776 47268 12782
rect 47216 12718 47268 12724
rect 46940 12708 46992 12714
rect 46940 12650 46992 12656
rect 46938 12472 46994 12481
rect 47032 12436 47084 12442
rect 46994 12416 47032 12434
rect 46938 12407 47032 12416
rect 46952 12406 47032 12407
rect 47032 12378 47084 12384
rect 46754 12336 46810 12345
rect 46754 12271 46810 12280
rect 46664 12096 46716 12102
rect 46664 12038 46716 12044
rect 46676 11694 46704 12038
rect 46664 11688 46716 11694
rect 46664 11630 46716 11636
rect 46768 11626 46796 12271
rect 46940 11892 46992 11898
rect 46940 11834 46992 11840
rect 46756 11620 46808 11626
rect 46756 11562 46808 11568
rect 46848 11076 46900 11082
rect 46848 11018 46900 11024
rect 46572 10260 46624 10266
rect 46572 10202 46624 10208
rect 46756 9580 46808 9586
rect 46756 9522 46808 9528
rect 46768 9382 46796 9522
rect 46296 9376 46348 9382
rect 46294 9344 46296 9353
rect 46756 9376 46808 9382
rect 46348 9344 46350 9353
rect 46756 9318 46808 9324
rect 46294 9279 46350 9288
rect 46664 8968 46716 8974
rect 46664 8910 46716 8916
rect 46388 8832 46440 8838
rect 46388 8774 46440 8780
rect 46400 8566 46428 8774
rect 46388 8560 46440 8566
rect 46388 8502 46440 8508
rect 46676 8430 46704 8910
rect 46664 8424 46716 8430
rect 46664 8366 46716 8372
rect 46768 8294 46796 9318
rect 46756 8288 46808 8294
rect 46756 8230 46808 8236
rect 46204 8084 46256 8090
rect 46204 8026 46256 8032
rect 46664 7744 46716 7750
rect 46664 7686 46716 7692
rect 46204 6792 46256 6798
rect 46204 6734 46256 6740
rect 46216 6118 46244 6734
rect 46572 6724 46624 6730
rect 46572 6666 46624 6672
rect 46584 6458 46612 6666
rect 46572 6452 46624 6458
rect 46572 6394 46624 6400
rect 46676 6322 46704 7686
rect 46664 6316 46716 6322
rect 46664 6258 46716 6264
rect 46204 6112 46256 6118
rect 46204 6054 46256 6060
rect 46112 4820 46164 4826
rect 46112 4762 46164 4768
rect 45468 4616 45520 4622
rect 45468 4558 45520 4564
rect 45468 4004 45520 4010
rect 45468 3946 45520 3952
rect 45480 3738 45508 3946
rect 45468 3732 45520 3738
rect 45468 3674 45520 3680
rect 46572 3528 46624 3534
rect 46572 3470 46624 3476
rect 46584 3058 46612 3470
rect 46860 3398 46888 11018
rect 46952 10062 46980 11834
rect 47228 10674 47256 12718
rect 47308 12096 47360 12102
rect 47308 12038 47360 12044
rect 47320 11218 47348 12038
rect 47688 11762 47716 15200
rect 48136 13728 48188 13734
rect 48136 13670 48188 13676
rect 47860 12844 47912 12850
rect 47780 12804 47860 12832
rect 47780 12102 47808 12804
rect 47860 12786 47912 12792
rect 48044 12844 48096 12850
rect 48044 12786 48096 12792
rect 48056 12434 48084 12786
rect 47964 12406 48084 12434
rect 47768 12096 47820 12102
rect 47768 12038 47820 12044
rect 47676 11756 47728 11762
rect 47676 11698 47728 11704
rect 47584 11552 47636 11558
rect 47584 11494 47636 11500
rect 47676 11552 47728 11558
rect 47676 11494 47728 11500
rect 47308 11212 47360 11218
rect 47308 11154 47360 11160
rect 47216 10668 47268 10674
rect 47216 10610 47268 10616
rect 47492 10260 47544 10266
rect 47492 10202 47544 10208
rect 47504 10062 47532 10202
rect 46940 10056 46992 10062
rect 46940 9998 46992 10004
rect 47308 10056 47360 10062
rect 47308 9998 47360 10004
rect 47492 10056 47544 10062
rect 47492 9998 47544 10004
rect 47124 9716 47176 9722
rect 47124 9658 47176 9664
rect 47032 9580 47084 9586
rect 47032 9522 47084 9528
rect 47044 9110 47072 9522
rect 47032 9104 47084 9110
rect 47032 9046 47084 9052
rect 47032 8288 47084 8294
rect 47032 8230 47084 8236
rect 47044 7954 47072 8230
rect 47032 7948 47084 7954
rect 47032 7890 47084 7896
rect 47044 7206 47072 7890
rect 47032 7200 47084 7206
rect 47032 7142 47084 7148
rect 47044 6730 47072 7142
rect 47032 6724 47084 6730
rect 47032 6666 47084 6672
rect 47136 5846 47164 9658
rect 47320 9382 47348 9998
rect 47308 9376 47360 9382
rect 47308 9318 47360 9324
rect 47216 8832 47268 8838
rect 47216 8774 47268 8780
rect 47124 5840 47176 5846
rect 47124 5782 47176 5788
rect 47228 5574 47256 8774
rect 47308 5840 47360 5846
rect 47308 5782 47360 5788
rect 47320 5574 47348 5782
rect 47216 5568 47268 5574
rect 47216 5510 47268 5516
rect 47308 5568 47360 5574
rect 47308 5510 47360 5516
rect 47216 4548 47268 4554
rect 47216 4490 47268 4496
rect 46848 3392 46900 3398
rect 46848 3334 46900 3340
rect 47228 3126 47256 4490
rect 47216 3120 47268 3126
rect 47216 3062 47268 3068
rect 46572 3052 46624 3058
rect 46572 2994 46624 3000
rect 47320 2514 47348 5510
rect 47596 3942 47624 11494
rect 47688 9586 47716 11494
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47780 9722 47808 10610
rect 47860 10464 47912 10470
rect 47860 10406 47912 10412
rect 47872 9994 47900 10406
rect 47860 9988 47912 9994
rect 47860 9930 47912 9936
rect 47768 9716 47820 9722
rect 47768 9658 47820 9664
rect 47676 9580 47728 9586
rect 47676 9522 47728 9528
rect 47688 9353 47716 9522
rect 47674 9344 47730 9353
rect 47674 9279 47730 9288
rect 47688 9042 47716 9279
rect 47964 9081 47992 12406
rect 48148 11898 48176 13670
rect 48136 11892 48188 11898
rect 48136 11834 48188 11840
rect 48240 11830 48268 15200
rect 48320 13252 48372 13258
rect 48320 13194 48372 13200
rect 48228 11824 48280 11830
rect 48228 11766 48280 11772
rect 48332 11286 48360 13194
rect 48792 12442 48820 15200
rect 48964 12980 49016 12986
rect 48964 12922 49016 12928
rect 48780 12436 48832 12442
rect 48780 12378 48832 12384
rect 48780 12164 48832 12170
rect 48780 12106 48832 12112
rect 48792 11937 48820 12106
rect 48778 11928 48834 11937
rect 48778 11863 48834 11872
rect 48780 11620 48832 11626
rect 48780 11562 48832 11568
rect 48320 11280 48372 11286
rect 48320 11222 48372 11228
rect 48504 11280 48556 11286
rect 48504 11222 48556 11228
rect 48596 11280 48648 11286
rect 48596 11222 48648 11228
rect 48412 11008 48464 11014
rect 48412 10950 48464 10956
rect 48424 10674 48452 10950
rect 48516 10810 48544 11222
rect 48608 11150 48636 11222
rect 48596 11144 48648 11150
rect 48596 11086 48648 11092
rect 48688 11144 48740 11150
rect 48688 11086 48740 11092
rect 48596 11008 48648 11014
rect 48596 10950 48648 10956
rect 48504 10804 48556 10810
rect 48504 10746 48556 10752
rect 48608 10742 48636 10950
rect 48596 10736 48648 10742
rect 48596 10678 48648 10684
rect 48412 10668 48464 10674
rect 48412 10610 48464 10616
rect 48044 10464 48096 10470
rect 48044 10406 48096 10412
rect 47950 9072 48006 9081
rect 47676 9036 47728 9042
rect 47950 9007 48006 9016
rect 47676 8978 47728 8984
rect 47952 7744 48004 7750
rect 47952 7686 48004 7692
rect 47964 4146 47992 7686
rect 47952 4140 48004 4146
rect 47952 4082 48004 4088
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 48056 3058 48084 10406
rect 48228 10124 48280 10130
rect 48228 10066 48280 10072
rect 48240 9722 48268 10066
rect 48412 9920 48464 9926
rect 48412 9862 48464 9868
rect 48228 9716 48280 9722
rect 48228 9658 48280 9664
rect 48136 9648 48188 9654
rect 48136 9590 48188 9596
rect 48148 8090 48176 9590
rect 48320 9104 48372 9110
rect 48320 9046 48372 9052
rect 48136 8084 48188 8090
rect 48136 8026 48188 8032
rect 48332 5302 48360 9046
rect 48424 8974 48452 9862
rect 48608 9586 48636 10678
rect 48700 10266 48728 11086
rect 48792 11082 48820 11562
rect 48780 11076 48832 11082
rect 48780 11018 48832 11024
rect 48778 10432 48834 10441
rect 48778 10367 48834 10376
rect 48688 10260 48740 10266
rect 48688 10202 48740 10208
rect 48792 10198 48820 10367
rect 48780 10192 48832 10198
rect 48780 10134 48832 10140
rect 48596 9580 48648 9586
rect 48596 9522 48648 9528
rect 48872 9580 48924 9586
rect 48872 9522 48924 9528
rect 48688 9376 48740 9382
rect 48688 9318 48740 9324
rect 48412 8968 48464 8974
rect 48412 8910 48464 8916
rect 48424 8242 48452 8910
rect 48424 8214 48544 8242
rect 48516 5914 48544 8214
rect 48596 6248 48648 6254
rect 48596 6190 48648 6196
rect 48608 5914 48636 6190
rect 48504 5908 48556 5914
rect 48504 5850 48556 5856
rect 48596 5908 48648 5914
rect 48596 5850 48648 5856
rect 48320 5296 48372 5302
rect 48320 5238 48372 5244
rect 48700 5234 48728 9318
rect 48884 8537 48912 9522
rect 48870 8528 48926 8537
rect 48870 8463 48872 8472
rect 48924 8463 48926 8472
rect 48872 8434 48924 8440
rect 48884 8403 48912 8434
rect 48688 5228 48740 5234
rect 48688 5170 48740 5176
rect 48976 3942 49004 12922
rect 49148 12640 49200 12646
rect 49148 12582 49200 12588
rect 49160 11762 49188 12582
rect 49344 12434 49372 15200
rect 49712 13410 49740 15286
rect 49882 15200 49938 15286
rect 50434 15200 50490 16000
rect 50986 15200 51042 16000
rect 51538 15314 51594 16000
rect 51276 15286 51594 15314
rect 49792 13456 49844 13462
rect 49620 13382 49740 13410
rect 49790 13424 49792 13433
rect 49844 13424 49846 13433
rect 49620 12714 49648 13382
rect 49790 13359 49846 13368
rect 49700 13320 49752 13326
rect 49700 13262 49752 13268
rect 49884 13320 49936 13326
rect 49884 13262 49936 13268
rect 49608 12708 49660 12714
rect 49608 12650 49660 12656
rect 49252 12406 49372 12434
rect 49148 11756 49200 11762
rect 49148 11698 49200 11704
rect 49252 11694 49280 12406
rect 49712 12238 49740 13262
rect 49792 13184 49844 13190
rect 49792 13126 49844 13132
rect 49804 12238 49832 13126
rect 49700 12232 49752 12238
rect 49700 12174 49752 12180
rect 49792 12232 49844 12238
rect 49792 12174 49844 12180
rect 49516 11824 49568 11830
rect 49516 11766 49568 11772
rect 49332 11756 49384 11762
rect 49332 11698 49384 11704
rect 49240 11688 49292 11694
rect 49240 11630 49292 11636
rect 49056 11552 49108 11558
rect 49056 11494 49108 11500
rect 49068 5846 49096 11494
rect 49148 11144 49200 11150
rect 49148 11086 49200 11092
rect 49160 10985 49188 11086
rect 49240 11076 49292 11082
rect 49240 11018 49292 11024
rect 49146 10976 49202 10985
rect 49146 10911 49202 10920
rect 49146 10296 49202 10305
rect 49146 10231 49202 10240
rect 49160 9994 49188 10231
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 49252 9450 49280 11018
rect 49240 9444 49292 9450
rect 49240 9386 49292 9392
rect 49240 8832 49292 8838
rect 49240 8774 49292 8780
rect 49148 8492 49200 8498
rect 49148 8434 49200 8440
rect 49160 8090 49188 8434
rect 49148 8084 49200 8090
rect 49148 8026 49200 8032
rect 49056 5840 49108 5846
rect 49056 5782 49108 5788
rect 49252 4826 49280 8774
rect 49344 8022 49372 11698
rect 49528 11218 49556 11766
rect 49516 11212 49568 11218
rect 49516 11154 49568 11160
rect 49424 10804 49476 10810
rect 49424 10746 49476 10752
rect 49436 10606 49464 10746
rect 49424 10600 49476 10606
rect 49424 10542 49476 10548
rect 49516 10532 49568 10538
rect 49516 10474 49568 10480
rect 49528 9994 49556 10474
rect 49712 10062 49740 12174
rect 49792 11688 49844 11694
rect 49896 11676 49924 13262
rect 50448 12434 50476 15200
rect 50712 13932 50764 13938
rect 50712 13874 50764 13880
rect 50620 13796 50672 13802
rect 50620 13738 50672 13744
rect 50528 12844 50580 12850
rect 50528 12786 50580 12792
rect 50356 12406 50476 12434
rect 50252 12232 50304 12238
rect 50252 12174 50304 12180
rect 50160 12164 50212 12170
rect 50160 12106 50212 12112
rect 50068 11756 50120 11762
rect 50068 11698 50120 11704
rect 49844 11648 49924 11676
rect 49792 11630 49844 11636
rect 49804 11218 49832 11630
rect 49792 11212 49844 11218
rect 49792 11154 49844 11160
rect 49884 10668 49936 10674
rect 49884 10610 49936 10616
rect 49700 10056 49752 10062
rect 49620 10016 49700 10044
rect 49516 9988 49568 9994
rect 49516 9930 49568 9936
rect 49516 9444 49568 9450
rect 49516 9386 49568 9392
rect 49528 9110 49556 9386
rect 49620 9178 49648 10016
rect 49700 9998 49752 10004
rect 49896 9722 49924 10610
rect 49976 10056 50028 10062
rect 49976 9998 50028 10004
rect 49884 9716 49936 9722
rect 49884 9658 49936 9664
rect 49700 9648 49752 9654
rect 49700 9590 49752 9596
rect 49712 9178 49740 9590
rect 49792 9580 49844 9586
rect 49792 9522 49844 9528
rect 49608 9172 49660 9178
rect 49608 9114 49660 9120
rect 49700 9172 49752 9178
rect 49700 9114 49752 9120
rect 49424 9104 49476 9110
rect 49424 9046 49476 9052
rect 49516 9104 49568 9110
rect 49516 9046 49568 9052
rect 49436 8634 49464 9046
rect 49424 8628 49476 8634
rect 49424 8570 49476 8576
rect 49528 8090 49556 9046
rect 49516 8084 49568 8090
rect 49516 8026 49568 8032
rect 49332 8016 49384 8022
rect 49332 7958 49384 7964
rect 49528 7818 49556 8026
rect 49516 7812 49568 7818
rect 49516 7754 49568 7760
rect 49528 7478 49556 7754
rect 49620 7546 49648 9114
rect 49804 9058 49832 9522
rect 49884 9104 49936 9110
rect 49804 9052 49884 9058
rect 49804 9046 49936 9052
rect 49804 9030 49924 9046
rect 49804 8430 49832 9030
rect 49988 8838 50016 9998
rect 50080 8838 50108 11698
rect 50172 10849 50200 12106
rect 50158 10840 50214 10849
rect 50158 10775 50214 10784
rect 49976 8832 50028 8838
rect 49976 8774 50028 8780
rect 50068 8832 50120 8838
rect 50068 8774 50120 8780
rect 49792 8424 49844 8430
rect 49792 8366 49844 8372
rect 49700 8084 49752 8090
rect 49700 8026 49752 8032
rect 49608 7540 49660 7546
rect 49608 7482 49660 7488
rect 49516 7472 49568 7478
rect 49516 7414 49568 7420
rect 49712 7410 49740 8026
rect 49804 7750 49832 8366
rect 49792 7744 49844 7750
rect 49792 7686 49844 7692
rect 49804 7546 49832 7686
rect 49792 7540 49844 7546
rect 49792 7482 49844 7488
rect 49700 7404 49752 7410
rect 49700 7346 49752 7352
rect 50264 6186 50292 12174
rect 50356 10266 50384 12406
rect 50436 11008 50488 11014
rect 50436 10950 50488 10956
rect 50448 10674 50476 10950
rect 50436 10668 50488 10674
rect 50436 10610 50488 10616
rect 50436 10532 50488 10538
rect 50436 10474 50488 10480
rect 50344 10260 50396 10266
rect 50344 10202 50396 10208
rect 50344 9036 50396 9042
rect 50344 8978 50396 8984
rect 50356 7954 50384 8978
rect 50448 8566 50476 10474
rect 50436 8560 50488 8566
rect 50436 8502 50488 8508
rect 50344 7948 50396 7954
rect 50344 7890 50396 7896
rect 50540 6934 50568 12786
rect 50632 9926 50660 13738
rect 50724 13734 50752 13874
rect 50712 13728 50764 13734
rect 50712 13670 50764 13676
rect 50896 13524 50948 13530
rect 50896 13466 50948 13472
rect 50712 13184 50764 13190
rect 50712 13126 50764 13132
rect 50804 13184 50856 13190
rect 50804 13126 50856 13132
rect 50724 12889 50752 13126
rect 50710 12880 50766 12889
rect 50710 12815 50766 12824
rect 50816 12782 50844 13126
rect 50908 13025 50936 13466
rect 50894 13016 50950 13025
rect 50894 12951 50950 12960
rect 50804 12776 50856 12782
rect 50804 12718 50856 12724
rect 50896 12640 50948 12646
rect 50896 12582 50948 12588
rect 50908 12345 50936 12582
rect 50894 12336 50950 12345
rect 50894 12271 50950 12280
rect 51000 11898 51028 15200
rect 51080 14068 51132 14074
rect 51080 14010 51132 14016
rect 51092 12306 51120 14010
rect 51170 13016 51226 13025
rect 51170 12951 51226 12960
rect 51184 12850 51212 12951
rect 51172 12844 51224 12850
rect 51172 12786 51224 12792
rect 51080 12300 51132 12306
rect 51080 12242 51132 12248
rect 50988 11892 51040 11898
rect 50988 11834 51040 11840
rect 51080 11688 51132 11694
rect 51080 11630 51132 11636
rect 50710 11520 50766 11529
rect 50710 11455 50766 11464
rect 50620 9920 50672 9926
rect 50620 9862 50672 9868
rect 50620 9648 50672 9654
rect 50620 9590 50672 9596
rect 50632 7818 50660 9590
rect 50620 7812 50672 7818
rect 50620 7754 50672 7760
rect 50528 6928 50580 6934
rect 50528 6870 50580 6876
rect 50436 6860 50488 6866
rect 50436 6802 50488 6808
rect 50252 6180 50304 6186
rect 50252 6122 50304 6128
rect 49240 4820 49292 4826
rect 49240 4762 49292 4768
rect 50448 4758 50476 6802
rect 50724 6730 50752 11455
rect 50896 11144 50948 11150
rect 50816 11092 50896 11098
rect 50816 11086 50948 11092
rect 50816 11070 50936 11086
rect 51092 11082 51120 11630
rect 51080 11076 51132 11082
rect 50816 9654 50844 11070
rect 51080 11018 51132 11024
rect 51170 10976 51226 10985
rect 51170 10911 51226 10920
rect 50896 10668 50948 10674
rect 50896 10610 50948 10616
rect 50804 9648 50856 9654
rect 50804 9590 50856 9596
rect 50804 8832 50856 8838
rect 50804 8774 50856 8780
rect 50816 7274 50844 8774
rect 50804 7268 50856 7274
rect 50804 7210 50856 7216
rect 50712 6724 50764 6730
rect 50712 6666 50764 6672
rect 50724 6390 50752 6666
rect 50712 6384 50764 6390
rect 50712 6326 50764 6332
rect 50804 6316 50856 6322
rect 50804 6258 50856 6264
rect 50816 6118 50844 6258
rect 50804 6112 50856 6118
rect 50804 6054 50856 6060
rect 50436 4752 50488 4758
rect 50436 4694 50488 4700
rect 49792 4072 49844 4078
rect 49792 4014 49844 4020
rect 48964 3936 49016 3942
rect 48964 3878 49016 3884
rect 49700 3460 49752 3466
rect 49700 3402 49752 3408
rect 49608 3392 49660 3398
rect 49606 3360 49608 3369
rect 49660 3360 49662 3369
rect 49606 3295 49662 3304
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 49712 2922 49740 3402
rect 49804 3058 49832 4014
rect 50816 3194 50844 6054
rect 50908 3738 50936 10610
rect 51184 10606 51212 10911
rect 51172 10600 51224 10606
rect 51092 10560 51172 10588
rect 51092 8430 51120 10560
rect 51172 10542 51224 10548
rect 51276 10266 51304 15286
rect 51538 15200 51594 15286
rect 52090 15200 52146 16000
rect 52642 15200 52698 16000
rect 53194 15314 53250 16000
rect 53194 15286 53420 15314
rect 53194 15200 53250 15286
rect 51632 12640 51684 12646
rect 51632 12582 51684 12588
rect 51448 12368 51500 12374
rect 51448 12310 51500 12316
rect 51264 10260 51316 10266
rect 51264 10202 51316 10208
rect 51460 10062 51488 12310
rect 51644 12238 51672 12582
rect 51632 12232 51684 12238
rect 51632 12174 51684 12180
rect 51724 12232 51776 12238
rect 51724 12174 51776 12180
rect 51540 11688 51592 11694
rect 51540 11630 51592 11636
rect 51552 10169 51580 11630
rect 51632 11348 51684 11354
rect 51632 11290 51684 11296
rect 51644 11257 51672 11290
rect 51630 11248 51686 11257
rect 51736 11218 51764 12174
rect 52000 12164 52052 12170
rect 52000 12106 52052 12112
rect 51908 11756 51960 11762
rect 51828 11716 51908 11744
rect 51630 11183 51686 11192
rect 51724 11212 51776 11218
rect 51724 11154 51776 11160
rect 51538 10160 51594 10169
rect 51538 10095 51594 10104
rect 51172 10056 51224 10062
rect 51172 9998 51224 10004
rect 51448 10056 51500 10062
rect 51448 9998 51500 10004
rect 51184 9382 51212 9998
rect 51460 9654 51488 9998
rect 51448 9648 51500 9654
rect 51448 9590 51500 9596
rect 51172 9376 51224 9382
rect 51172 9318 51224 9324
rect 51460 8634 51488 9590
rect 51448 8628 51500 8634
rect 51448 8570 51500 8576
rect 51080 8424 51132 8430
rect 51080 8366 51132 8372
rect 51356 8424 51408 8430
rect 51356 8366 51408 8372
rect 50988 8356 51040 8362
rect 50988 8298 51040 8304
rect 51000 4214 51028 8298
rect 51092 5166 51120 8366
rect 51368 7954 51396 8366
rect 51828 7970 51856 11716
rect 51908 11698 51960 11704
rect 51908 10668 51960 10674
rect 51908 10610 51960 10616
rect 51920 8294 51948 10610
rect 52012 10062 52040 12106
rect 52104 11694 52132 15200
rect 52368 12776 52420 12782
rect 52368 12718 52420 12724
rect 52380 12442 52408 12718
rect 52368 12436 52420 12442
rect 52368 12378 52420 12384
rect 52368 11892 52420 11898
rect 52368 11834 52420 11840
rect 52092 11688 52144 11694
rect 52092 11630 52144 11636
rect 52182 10160 52238 10169
rect 52182 10095 52238 10104
rect 52000 10056 52052 10062
rect 52000 9998 52052 10004
rect 52196 9382 52224 10095
rect 52184 9376 52236 9382
rect 52184 9318 52236 9324
rect 52196 8650 52224 9318
rect 52104 8622 52316 8650
rect 52104 8430 52132 8622
rect 52288 8498 52316 8622
rect 52184 8492 52236 8498
rect 52184 8434 52236 8440
rect 52276 8492 52328 8498
rect 52276 8434 52328 8440
rect 52092 8424 52144 8430
rect 52092 8366 52144 8372
rect 51908 8288 51960 8294
rect 51908 8230 51960 8236
rect 51356 7948 51408 7954
rect 51356 7890 51408 7896
rect 51736 7942 51856 7970
rect 51080 5160 51132 5166
rect 51080 5102 51132 5108
rect 50988 4208 51040 4214
rect 50988 4150 51040 4156
rect 50896 3732 50948 3738
rect 50896 3674 50948 3680
rect 51092 3398 51120 5102
rect 51080 3392 51132 3398
rect 51080 3334 51132 3340
rect 50804 3188 50856 3194
rect 50804 3130 50856 3136
rect 51092 3058 51120 3334
rect 49792 3052 49844 3058
rect 49792 2994 49844 3000
rect 51080 3052 51132 3058
rect 51080 2994 51132 3000
rect 49700 2916 49752 2922
rect 49700 2858 49752 2864
rect 49804 2774 49832 2994
rect 51736 2854 51764 7942
rect 51816 7880 51868 7886
rect 51816 7822 51868 7828
rect 51828 6390 51856 7822
rect 51920 7750 51948 8230
rect 51908 7744 51960 7750
rect 51908 7686 51960 7692
rect 52104 6866 52132 8366
rect 52092 6860 52144 6866
rect 52092 6802 52144 6808
rect 52196 6730 52224 8434
rect 52380 7868 52408 11834
rect 52460 11756 52512 11762
rect 52460 11698 52512 11704
rect 52472 10266 52500 11698
rect 52552 11552 52604 11558
rect 52550 11520 52552 11529
rect 52604 11520 52606 11529
rect 52550 11455 52606 11464
rect 52552 11076 52604 11082
rect 52552 11018 52604 11024
rect 52564 10713 52592 11018
rect 52656 10810 52684 15200
rect 52920 13388 52972 13394
rect 52920 13330 52972 13336
rect 52826 11928 52882 11937
rect 52826 11863 52828 11872
rect 52880 11863 52882 11872
rect 52828 11834 52880 11840
rect 52644 10804 52696 10810
rect 52644 10746 52696 10752
rect 52550 10704 52606 10713
rect 52550 10639 52606 10648
rect 52644 10668 52696 10674
rect 52644 10610 52696 10616
rect 52460 10260 52512 10266
rect 52460 10202 52512 10208
rect 52656 10146 52684 10610
rect 52472 10130 52684 10146
rect 52460 10124 52696 10130
rect 52512 10118 52644 10124
rect 52460 10066 52512 10072
rect 52644 10066 52696 10072
rect 52932 9466 52960 13330
rect 53012 13184 53064 13190
rect 53012 13126 53064 13132
rect 53024 12714 53052 13126
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 53012 12708 53064 12714
rect 53012 12650 53064 12656
rect 53208 12434 53236 12786
rect 53208 12406 53328 12434
rect 53012 12164 53064 12170
rect 53012 12106 53064 12112
rect 53024 11694 53052 12106
rect 53012 11688 53064 11694
rect 53012 11630 53064 11636
rect 53102 10704 53158 10713
rect 53102 10639 53158 10648
rect 53012 10600 53064 10606
rect 53012 10542 53064 10548
rect 53024 9586 53052 10542
rect 53012 9580 53064 9586
rect 53012 9522 53064 9528
rect 52840 9450 52960 9466
rect 52828 9444 52960 9450
rect 52880 9438 52960 9444
rect 52828 9386 52880 9392
rect 52736 8832 52788 8838
rect 52736 8774 52788 8780
rect 52552 8492 52604 8498
rect 52552 8434 52604 8440
rect 52564 7954 52592 8434
rect 52748 8430 52776 8774
rect 52736 8424 52788 8430
rect 52736 8366 52788 8372
rect 52552 7948 52604 7954
rect 52552 7890 52604 7896
rect 52460 7880 52512 7886
rect 52380 7840 52460 7868
rect 52460 7822 52512 7828
rect 52276 7812 52328 7818
rect 52276 7754 52328 7760
rect 52288 6798 52316 7754
rect 53116 7410 53144 10639
rect 53300 9994 53328 12406
rect 53196 9988 53248 9994
rect 53196 9930 53248 9936
rect 53288 9988 53340 9994
rect 53288 9930 53340 9936
rect 53104 7404 53156 7410
rect 53104 7346 53156 7352
rect 52368 7336 52420 7342
rect 52368 7278 52420 7284
rect 52380 7002 52408 7278
rect 52368 6996 52420 7002
rect 52368 6938 52420 6944
rect 52276 6792 52328 6798
rect 52276 6734 52328 6740
rect 52184 6724 52236 6730
rect 52184 6666 52236 6672
rect 53208 6458 53236 9930
rect 53392 9178 53420 15286
rect 53746 15200 53802 16000
rect 54298 15200 54354 16000
rect 54850 15200 54906 16000
rect 55402 15314 55458 16000
rect 55232 15286 55458 15314
rect 53760 14074 53788 15200
rect 53748 14068 53800 14074
rect 53748 14010 53800 14016
rect 53564 13320 53616 13326
rect 53616 13280 53696 13308
rect 53564 13262 53616 13268
rect 53472 12912 53524 12918
rect 53472 12854 53524 12860
rect 53484 11354 53512 12854
rect 53668 12850 53696 13280
rect 54312 12986 54340 15200
rect 54300 12980 54352 12986
rect 54300 12922 54352 12928
rect 54392 12980 54444 12986
rect 54392 12922 54444 12928
rect 54404 12866 54432 12922
rect 54128 12850 54432 12866
rect 53656 12844 53708 12850
rect 53656 12786 53708 12792
rect 54116 12844 54432 12850
rect 54168 12838 54432 12844
rect 54760 12844 54812 12850
rect 54116 12786 54168 12792
rect 54760 12786 54812 12792
rect 54036 12714 54432 12730
rect 54024 12708 54432 12714
rect 54076 12702 54432 12708
rect 54024 12650 54076 12656
rect 54404 12646 54432 12702
rect 54300 12640 54352 12646
rect 54300 12582 54352 12588
rect 54392 12640 54444 12646
rect 54392 12582 54444 12588
rect 54312 12374 54340 12582
rect 54300 12368 54352 12374
rect 54300 12310 54352 12316
rect 54300 12232 54352 12238
rect 54300 12174 54352 12180
rect 54312 11898 54340 12174
rect 54576 12096 54628 12102
rect 54576 12038 54628 12044
rect 54300 11892 54352 11898
rect 54300 11834 54352 11840
rect 54392 11892 54444 11898
rect 54392 11834 54444 11840
rect 53564 11756 53616 11762
rect 53564 11698 53616 11704
rect 53472 11348 53524 11354
rect 53472 11290 53524 11296
rect 53576 10742 53604 11698
rect 54024 11688 54076 11694
rect 53930 11656 53986 11665
rect 54024 11630 54076 11636
rect 53930 11591 53986 11600
rect 53838 10840 53894 10849
rect 53838 10775 53894 10784
rect 53564 10736 53616 10742
rect 53564 10678 53616 10684
rect 53852 9654 53880 10775
rect 53840 9648 53892 9654
rect 53840 9590 53892 9596
rect 53472 9580 53524 9586
rect 53472 9522 53524 9528
rect 53380 9172 53432 9178
rect 53380 9114 53432 9120
rect 53380 8968 53432 8974
rect 53380 8910 53432 8916
rect 53392 8566 53420 8910
rect 53484 8838 53512 9522
rect 53840 8968 53892 8974
rect 53840 8910 53892 8916
rect 53472 8832 53524 8838
rect 53472 8774 53524 8780
rect 53380 8560 53432 8566
rect 53380 8502 53432 8508
rect 53748 7744 53800 7750
rect 53748 7686 53800 7692
rect 53380 6656 53432 6662
rect 53380 6598 53432 6604
rect 52368 6452 52420 6458
rect 52368 6394 52420 6400
rect 53196 6452 53248 6458
rect 53196 6394 53248 6400
rect 51816 6384 51868 6390
rect 51816 6326 51868 6332
rect 52276 5160 52328 5166
rect 52276 5102 52328 5108
rect 52288 4622 52316 5102
rect 52276 4616 52328 4622
rect 52276 4558 52328 4564
rect 52380 3602 52408 6394
rect 53392 6322 53420 6598
rect 53380 6316 53432 6322
rect 53380 6258 53432 6264
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 53760 3534 53788 7686
rect 53852 7410 53880 8910
rect 53944 8362 53972 11591
rect 54036 10198 54064 11630
rect 54404 11558 54432 11834
rect 54392 11552 54444 11558
rect 54392 11494 54444 11500
rect 54024 10192 54076 10198
rect 54024 10134 54076 10140
rect 54390 10160 54446 10169
rect 54036 9042 54064 10134
rect 54390 10095 54392 10104
rect 54444 10095 54446 10104
rect 54392 10066 54444 10072
rect 54206 10024 54262 10033
rect 54588 9994 54616 12038
rect 54772 10010 54800 12786
rect 54864 12238 54892 15200
rect 54852 12232 54904 12238
rect 54852 12174 54904 12180
rect 55126 12200 55182 12209
rect 55126 12135 55182 12144
rect 55036 10056 55088 10062
rect 54206 9959 54262 9968
rect 54576 9988 54628 9994
rect 54114 9888 54170 9897
rect 54114 9823 54170 9832
rect 54024 9036 54076 9042
rect 54024 8978 54076 8984
rect 54128 8974 54156 9823
rect 54220 9722 54248 9959
rect 54772 9982 54984 10010
rect 55036 9998 55088 10004
rect 54576 9930 54628 9936
rect 54956 9926 54984 9982
rect 54392 9920 54444 9926
rect 54392 9862 54444 9868
rect 54852 9920 54904 9926
rect 54852 9862 54904 9868
rect 54944 9920 54996 9926
rect 54944 9862 54996 9868
rect 54208 9716 54260 9722
rect 54208 9658 54260 9664
rect 54404 9674 54432 9862
rect 54404 9654 54524 9674
rect 54404 9648 54536 9654
rect 54404 9646 54484 9648
rect 54484 9590 54536 9596
rect 54300 9580 54352 9586
rect 54300 9522 54352 9528
rect 54208 9376 54260 9382
rect 54208 9318 54260 9324
rect 54220 9110 54248 9318
rect 54208 9104 54260 9110
rect 54208 9046 54260 9052
rect 54312 8974 54340 9522
rect 54116 8968 54168 8974
rect 54116 8910 54168 8916
rect 54300 8968 54352 8974
rect 54300 8910 54352 8916
rect 54116 8424 54168 8430
rect 54116 8366 54168 8372
rect 53932 8356 53984 8362
rect 53932 8298 53984 8304
rect 54128 7886 54156 8366
rect 54208 8288 54260 8294
rect 54208 8230 54260 8236
rect 54220 7886 54248 8230
rect 54116 7880 54168 7886
rect 54116 7822 54168 7828
rect 54208 7880 54260 7886
rect 54208 7822 54260 7828
rect 53840 7404 53892 7410
rect 53840 7346 53892 7352
rect 54128 6322 54156 7822
rect 54220 7002 54248 7822
rect 54312 7410 54340 8910
rect 54576 8832 54628 8838
rect 54576 8774 54628 8780
rect 54588 8294 54616 8774
rect 54576 8288 54628 8294
rect 54576 8230 54628 8236
rect 54760 7744 54812 7750
rect 54760 7686 54812 7692
rect 54772 7478 54800 7686
rect 54760 7472 54812 7478
rect 54760 7414 54812 7420
rect 54300 7404 54352 7410
rect 54300 7346 54352 7352
rect 54208 6996 54260 7002
rect 54208 6938 54260 6944
rect 54312 6798 54340 7346
rect 54300 6792 54352 6798
rect 54300 6734 54352 6740
rect 54116 6316 54168 6322
rect 54116 6258 54168 6264
rect 54208 6180 54260 6186
rect 54208 6122 54260 6128
rect 54220 5710 54248 6122
rect 54864 6118 54892 9862
rect 54944 8832 54996 8838
rect 54944 8774 54996 8780
rect 54956 7886 54984 8774
rect 54944 7880 54996 7886
rect 54944 7822 54996 7828
rect 54852 6112 54904 6118
rect 54852 6054 54904 6060
rect 54668 5772 54720 5778
rect 54668 5714 54720 5720
rect 54208 5704 54260 5710
rect 54208 5646 54260 5652
rect 54680 3942 54708 5714
rect 55048 5370 55076 9998
rect 55140 8548 55168 12135
rect 55232 11830 55260 15286
rect 55402 15200 55458 15286
rect 55954 15314 56010 16000
rect 55954 15286 56272 15314
rect 55954 15200 56010 15286
rect 55864 13456 55916 13462
rect 55864 13398 55916 13404
rect 55404 13320 55456 13326
rect 55404 13262 55456 13268
rect 55588 13320 55640 13326
rect 55588 13262 55640 13268
rect 55416 13161 55444 13262
rect 55402 13152 55458 13161
rect 55402 13087 55458 13096
rect 55600 12442 55628 13262
rect 55680 12912 55732 12918
rect 55680 12854 55732 12860
rect 55692 12782 55720 12854
rect 55680 12776 55732 12782
rect 55680 12718 55732 12724
rect 55588 12436 55640 12442
rect 55588 12378 55640 12384
rect 55312 12096 55364 12102
rect 55312 12038 55364 12044
rect 55496 12096 55548 12102
rect 55496 12038 55548 12044
rect 55324 11830 55352 12038
rect 55220 11824 55272 11830
rect 55220 11766 55272 11772
rect 55312 11824 55364 11830
rect 55312 11766 55364 11772
rect 55404 11280 55456 11286
rect 55404 11222 55456 11228
rect 55312 11144 55364 11150
rect 55312 11086 55364 11092
rect 55220 11076 55272 11082
rect 55220 11018 55272 11024
rect 55232 10742 55260 11018
rect 55220 10736 55272 10742
rect 55220 10678 55272 10684
rect 55324 10606 55352 11086
rect 55312 10600 55364 10606
rect 55312 10542 55364 10548
rect 55324 10470 55352 10542
rect 55312 10464 55364 10470
rect 55312 10406 55364 10412
rect 55416 8974 55444 11222
rect 55508 9586 55536 12038
rect 55600 11150 55628 12378
rect 55692 12322 55720 12718
rect 55692 12294 55812 12322
rect 55680 12232 55732 12238
rect 55680 12174 55732 12180
rect 55588 11144 55640 11150
rect 55588 11086 55640 11092
rect 55600 9674 55628 11086
rect 55692 11082 55720 12174
rect 55784 11694 55812 12294
rect 55772 11688 55824 11694
rect 55772 11630 55824 11636
rect 55680 11076 55732 11082
rect 55680 11018 55732 11024
rect 55692 10810 55720 11018
rect 55680 10804 55732 10810
rect 55680 10746 55732 10752
rect 55784 10606 55812 11630
rect 55772 10600 55824 10606
rect 55772 10542 55824 10548
rect 55600 9646 55720 9674
rect 55496 9580 55548 9586
rect 55496 9522 55548 9528
rect 55404 8968 55456 8974
rect 55404 8910 55456 8916
rect 55220 8560 55272 8566
rect 55140 8520 55220 8548
rect 55220 8502 55272 8508
rect 55692 8498 55720 9646
rect 55876 9178 55904 13398
rect 56048 13252 56100 13258
rect 56100 13212 56180 13240
rect 56048 13194 56100 13200
rect 56046 12880 56102 12889
rect 56046 12815 56048 12824
rect 56100 12815 56102 12824
rect 56048 12786 56100 12792
rect 56152 12442 56180 13212
rect 56140 12436 56192 12442
rect 56140 12378 56192 12384
rect 55954 12336 56010 12345
rect 55954 12271 56010 12280
rect 55968 12238 55996 12271
rect 55956 12232 56008 12238
rect 55956 12174 56008 12180
rect 56048 12232 56100 12238
rect 56048 12174 56100 12180
rect 55968 11014 55996 12174
rect 56060 11898 56088 12174
rect 56048 11892 56100 11898
rect 56048 11834 56100 11840
rect 56140 11688 56192 11694
rect 56140 11630 56192 11636
rect 56152 11082 56180 11630
rect 56140 11076 56192 11082
rect 56140 11018 56192 11024
rect 55956 11008 56008 11014
rect 55956 10950 56008 10956
rect 56048 10668 56100 10674
rect 56048 10610 56100 10616
rect 55956 10192 56008 10198
rect 55954 10160 55956 10169
rect 56008 10160 56010 10169
rect 55954 10095 56010 10104
rect 55864 9172 55916 9178
rect 55864 9114 55916 9120
rect 55680 8492 55732 8498
rect 55680 8434 55732 8440
rect 56060 8362 56088 10610
rect 56152 8634 56180 11018
rect 56244 10198 56272 15286
rect 56506 15200 56562 16000
rect 57058 15314 57114 16000
rect 57610 15314 57666 16000
rect 56612 15286 57114 15314
rect 56322 13288 56378 13297
rect 56322 13223 56378 13232
rect 56336 12238 56364 13223
rect 56324 12232 56376 12238
rect 56324 12174 56376 12180
rect 56416 11824 56468 11830
rect 56416 11766 56468 11772
rect 56324 10804 56376 10810
rect 56324 10746 56376 10752
rect 56232 10192 56284 10198
rect 56232 10134 56284 10140
rect 56230 9616 56286 9625
rect 56230 9551 56232 9560
rect 56284 9551 56286 9560
rect 56232 9522 56284 9528
rect 56140 8628 56192 8634
rect 56140 8570 56192 8576
rect 56048 8356 56100 8362
rect 56048 8298 56100 8304
rect 56152 8090 56180 8570
rect 56140 8084 56192 8090
rect 56140 8026 56192 8032
rect 55772 6928 55824 6934
rect 55772 6870 55824 6876
rect 55404 6316 55456 6322
rect 55404 6258 55456 6264
rect 55036 5364 55088 5370
rect 55036 5306 55088 5312
rect 55416 5166 55444 6258
rect 55404 5160 55456 5166
rect 55404 5102 55456 5108
rect 55784 4010 55812 6870
rect 56336 6866 56364 10746
rect 56428 9382 56456 11766
rect 56520 11098 56548 15200
rect 56612 12288 56640 15286
rect 57058 15200 57114 15286
rect 57256 15286 57666 15314
rect 56692 13320 56744 13326
rect 56690 13288 56692 13297
rect 56744 13288 56746 13297
rect 56690 13223 56746 13232
rect 56968 12912 57020 12918
rect 56968 12854 57020 12860
rect 56876 12844 56928 12850
rect 56876 12786 56928 12792
rect 56784 12436 56836 12442
rect 56784 12378 56836 12384
rect 56692 12300 56744 12306
rect 56612 12260 56692 12288
rect 56692 12242 56744 12248
rect 56796 12102 56824 12378
rect 56784 12096 56836 12102
rect 56784 12038 56836 12044
rect 56520 11070 56640 11098
rect 56508 10736 56560 10742
rect 56508 10678 56560 10684
rect 56520 10441 56548 10678
rect 56506 10432 56562 10441
rect 56506 10367 56562 10376
rect 56612 9722 56640 11070
rect 56692 11008 56744 11014
rect 56692 10950 56744 10956
rect 56704 10062 56732 10950
rect 56888 10282 56916 12786
rect 56796 10254 56916 10282
rect 56692 10056 56744 10062
rect 56692 9998 56744 10004
rect 56796 9908 56824 10254
rect 56876 10056 56928 10062
rect 56876 9998 56928 10004
rect 56704 9880 56824 9908
rect 56600 9716 56652 9722
rect 56600 9658 56652 9664
rect 56704 9602 56732 9880
rect 56888 9636 56916 9998
rect 56612 9574 56732 9602
rect 56796 9608 56916 9636
rect 56612 9450 56640 9574
rect 56692 9512 56744 9518
rect 56692 9454 56744 9460
rect 56600 9444 56652 9450
rect 56600 9386 56652 9392
rect 56416 9376 56468 9382
rect 56416 9318 56468 9324
rect 56416 8832 56468 8838
rect 56416 8774 56468 8780
rect 56324 6860 56376 6866
rect 56324 6802 56376 6808
rect 55772 4004 55824 4010
rect 55772 3946 55824 3952
rect 54668 3936 54720 3942
rect 54668 3878 54720 3884
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 53564 3392 53616 3398
rect 53562 3360 53564 3369
rect 53616 3360 53618 3369
rect 53562 3295 53618 3304
rect 56428 3126 56456 8774
rect 56416 3120 56468 3126
rect 56416 3062 56468 3068
rect 51724 2848 51776 2854
rect 51724 2790 51776 2796
rect 56704 2774 56732 9454
rect 56796 8090 56824 9608
rect 56876 9512 56928 9518
rect 56876 9454 56928 9460
rect 56888 9178 56916 9454
rect 56980 9178 57008 12854
rect 57256 12374 57284 15286
rect 57610 15200 57666 15286
rect 58162 15314 58218 16000
rect 58162 15286 58480 15314
rect 58162 15200 58218 15286
rect 57520 13184 57572 13190
rect 57520 13126 57572 13132
rect 57428 12980 57480 12986
rect 57428 12922 57480 12928
rect 57244 12368 57296 12374
rect 57150 12336 57206 12345
rect 57244 12310 57296 12316
rect 57150 12271 57152 12280
rect 57204 12271 57206 12280
rect 57152 12242 57204 12248
rect 57060 12232 57112 12238
rect 57060 12174 57112 12180
rect 57244 12232 57296 12238
rect 57244 12174 57296 12180
rect 57336 12232 57388 12238
rect 57336 12174 57388 12180
rect 57072 10198 57100 12174
rect 57256 11898 57284 12174
rect 57244 11892 57296 11898
rect 57244 11834 57296 11840
rect 57348 11762 57376 12174
rect 57336 11756 57388 11762
rect 57336 11698 57388 11704
rect 57440 10538 57468 12922
rect 57428 10532 57480 10538
rect 57428 10474 57480 10480
rect 57532 10305 57560 13126
rect 58256 12844 58308 12850
rect 58256 12786 58308 12792
rect 57980 12640 58032 12646
rect 58164 12640 58216 12646
rect 57980 12582 58032 12588
rect 58084 12600 58164 12628
rect 57888 12436 57940 12442
rect 57888 12378 57940 12384
rect 57900 11762 57928 12378
rect 57888 11756 57940 11762
rect 57888 11698 57940 11704
rect 57704 11144 57756 11150
rect 57704 11086 57756 11092
rect 57716 10810 57744 11086
rect 57704 10804 57756 10810
rect 57704 10746 57756 10752
rect 57518 10296 57574 10305
rect 57518 10231 57574 10240
rect 57900 10198 57928 11698
rect 57060 10192 57112 10198
rect 57060 10134 57112 10140
rect 57612 10192 57664 10198
rect 57612 10134 57664 10140
rect 57888 10192 57940 10198
rect 57888 10134 57940 10140
rect 57072 10033 57100 10134
rect 57058 10024 57114 10033
rect 57058 9959 57114 9968
rect 57624 9926 57652 10134
rect 57704 9988 57756 9994
rect 57704 9930 57756 9936
rect 57796 9988 57848 9994
rect 57796 9930 57848 9936
rect 57060 9920 57112 9926
rect 57060 9862 57112 9868
rect 57520 9920 57572 9926
rect 57520 9862 57572 9868
rect 57612 9920 57664 9926
rect 57612 9862 57664 9868
rect 57072 9722 57100 9862
rect 57060 9716 57112 9722
rect 57060 9658 57112 9664
rect 57152 9648 57204 9654
rect 57150 9616 57152 9625
rect 57204 9616 57206 9625
rect 57532 9586 57560 9862
rect 57716 9586 57744 9930
rect 57808 9897 57836 9930
rect 57794 9888 57850 9897
rect 57794 9823 57850 9832
rect 57150 9551 57206 9560
rect 57520 9580 57572 9586
rect 57520 9522 57572 9528
rect 57704 9580 57756 9586
rect 57704 9522 57756 9528
rect 56876 9172 56928 9178
rect 56876 9114 56928 9120
rect 56968 9172 57020 9178
rect 56968 9114 57020 9120
rect 57716 9110 57744 9522
rect 57704 9104 57756 9110
rect 57704 9046 57756 9052
rect 57992 8974 58020 12582
rect 58084 10742 58112 12600
rect 58164 12582 58216 12588
rect 58268 12442 58296 12786
rect 58256 12436 58308 12442
rect 58256 12378 58308 12384
rect 58164 11144 58216 11150
rect 58164 11086 58216 11092
rect 58072 10736 58124 10742
rect 58072 10678 58124 10684
rect 58072 10464 58124 10470
rect 58072 10406 58124 10412
rect 58084 9654 58112 10406
rect 58072 9648 58124 9654
rect 58072 9590 58124 9596
rect 58072 9376 58124 9382
rect 58072 9318 58124 9324
rect 57704 8968 57756 8974
rect 57704 8910 57756 8916
rect 57796 8968 57848 8974
rect 57796 8910 57848 8916
rect 57980 8968 58032 8974
rect 57980 8910 58032 8916
rect 57336 8832 57388 8838
rect 57336 8774 57388 8780
rect 57520 8832 57572 8838
rect 57520 8774 57572 8780
rect 57348 8498 57376 8774
rect 57336 8492 57388 8498
rect 57336 8434 57388 8440
rect 57532 8430 57560 8774
rect 57520 8424 57572 8430
rect 57520 8366 57572 8372
rect 56784 8084 56836 8090
rect 56784 8026 56836 8032
rect 57532 6798 57560 8366
rect 57716 7546 57744 8910
rect 57808 7546 57836 8910
rect 58084 8566 58112 9318
rect 58176 8906 58204 11086
rect 58346 10840 58402 10849
rect 58256 10804 58308 10810
rect 58346 10775 58402 10784
rect 58256 10746 58308 10752
rect 58164 8900 58216 8906
rect 58164 8842 58216 8848
rect 58268 8838 58296 10746
rect 58360 10674 58388 10775
rect 58348 10668 58400 10674
rect 58348 10610 58400 10616
rect 58452 9450 58480 15286
rect 58714 15200 58770 16000
rect 59266 15200 59322 16000
rect 59818 15200 59874 16000
rect 60370 15314 60426 16000
rect 60370 15286 60504 15314
rect 60370 15200 60426 15286
rect 58624 13320 58676 13326
rect 58624 13262 58676 13268
rect 58636 13025 58664 13262
rect 58622 13016 58678 13025
rect 58622 12951 58678 12960
rect 58636 11898 58664 12951
rect 58624 11892 58676 11898
rect 58624 11834 58676 11840
rect 58622 11248 58678 11257
rect 58622 11183 58678 11192
rect 58636 11150 58664 11183
rect 58624 11144 58676 11150
rect 58544 11104 58624 11132
rect 58440 9444 58492 9450
rect 58440 9386 58492 9392
rect 58256 8832 58308 8838
rect 58256 8774 58308 8780
rect 58072 8560 58124 8566
rect 58072 8502 58124 8508
rect 58544 7546 58572 11104
rect 58624 11086 58676 11092
rect 58624 10532 58676 10538
rect 58624 10474 58676 10480
rect 58636 8106 58664 10474
rect 58728 10198 58756 15200
rect 58808 13184 58860 13190
rect 58808 13126 58860 13132
rect 58820 12782 58848 13126
rect 58808 12776 58860 12782
rect 58808 12718 58860 12724
rect 59176 12776 59228 12782
rect 59176 12718 59228 12724
rect 58820 12345 58848 12718
rect 58806 12336 58862 12345
rect 58806 12271 58862 12280
rect 59084 11892 59136 11898
rect 59084 11834 59136 11840
rect 58808 11280 58860 11286
rect 58808 11222 58860 11228
rect 58716 10192 58768 10198
rect 58716 10134 58768 10140
rect 58820 10062 58848 11222
rect 58992 11144 59044 11150
rect 58992 11086 59044 11092
rect 59004 10169 59032 11086
rect 59096 10674 59124 11834
rect 59188 10810 59216 12718
rect 59280 11354 59308 15200
rect 59450 13424 59506 13433
rect 59450 13359 59506 13368
rect 59464 11898 59492 13359
rect 59544 12776 59596 12782
rect 59544 12718 59596 12724
rect 59556 12238 59584 12718
rect 59544 12232 59596 12238
rect 59544 12174 59596 12180
rect 59452 11892 59504 11898
rect 59452 11834 59504 11840
rect 59544 11756 59596 11762
rect 59544 11698 59596 11704
rect 59268 11348 59320 11354
rect 59268 11290 59320 11296
rect 59176 10804 59228 10810
rect 59176 10746 59228 10752
rect 59084 10668 59136 10674
rect 59084 10610 59136 10616
rect 58990 10160 59046 10169
rect 58990 10095 59046 10104
rect 58808 10056 58860 10062
rect 58808 9998 58860 10004
rect 58636 8078 58848 8106
rect 58820 8022 58848 8078
rect 58808 8016 58860 8022
rect 58808 7958 58860 7964
rect 57704 7540 57756 7546
rect 57704 7482 57756 7488
rect 57796 7540 57848 7546
rect 57796 7482 57848 7488
rect 58532 7540 58584 7546
rect 58532 7482 58584 7488
rect 57520 6792 57572 6798
rect 57520 6734 57572 6740
rect 57152 6724 57204 6730
rect 57152 6666 57204 6672
rect 56784 5024 56836 5030
rect 56784 4966 56836 4972
rect 56796 4282 56824 4966
rect 56784 4276 56836 4282
rect 56784 4218 56836 4224
rect 57164 3398 57192 6666
rect 58624 6656 58676 6662
rect 58624 6598 58676 6604
rect 58636 5710 58664 6598
rect 58624 5704 58676 5710
rect 58624 5646 58676 5652
rect 58440 5568 58492 5574
rect 58440 5510 58492 5516
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57152 3392 57204 3398
rect 57152 3334 57204 3340
rect 57256 2922 57284 3538
rect 58452 3534 58480 5510
rect 58820 5234 58848 7958
rect 59004 6866 59032 10095
rect 59096 8294 59124 10610
rect 59188 10606 59216 10746
rect 59176 10600 59228 10606
rect 59176 10542 59228 10548
rect 59084 8288 59136 8294
rect 59084 8230 59136 8236
rect 59096 7886 59124 8230
rect 59556 8090 59584 11698
rect 59832 10198 59860 15200
rect 60117 13628 60425 13637
rect 60117 13626 60123 13628
rect 60179 13626 60203 13628
rect 60259 13626 60283 13628
rect 60339 13626 60363 13628
rect 60419 13626 60425 13628
rect 60179 13574 60181 13626
rect 60361 13574 60363 13626
rect 60117 13572 60123 13574
rect 60179 13572 60203 13574
rect 60259 13572 60283 13574
rect 60339 13572 60363 13574
rect 60419 13572 60425 13574
rect 60117 13563 60425 13572
rect 60370 13288 60426 13297
rect 60370 13223 60372 13232
rect 60424 13223 60426 13232
rect 60372 13194 60424 13200
rect 60117 12540 60425 12549
rect 60117 12538 60123 12540
rect 60179 12538 60203 12540
rect 60259 12538 60283 12540
rect 60339 12538 60363 12540
rect 60419 12538 60425 12540
rect 60179 12486 60181 12538
rect 60361 12486 60363 12538
rect 60117 12484 60123 12486
rect 60179 12484 60203 12486
rect 60259 12484 60283 12486
rect 60339 12484 60363 12486
rect 60419 12484 60425 12486
rect 60117 12475 60425 12484
rect 60476 12434 60504 15286
rect 60922 15200 60978 16000
rect 61474 15200 61530 16000
rect 62026 15200 62082 16000
rect 62578 15200 62634 16000
rect 63130 15314 63186 16000
rect 63682 15314 63738 16000
rect 64234 15314 64290 16000
rect 63130 15286 63264 15314
rect 63130 15200 63186 15286
rect 60556 13796 60608 13802
rect 60556 13738 60608 13744
rect 60568 12850 60596 13738
rect 60648 13456 60700 13462
rect 60648 13398 60700 13404
rect 60660 13326 60688 13398
rect 60648 13320 60700 13326
rect 60648 13262 60700 13268
rect 60740 13320 60792 13326
rect 60740 13262 60792 13268
rect 60832 13320 60884 13326
rect 60832 13262 60884 13268
rect 60648 13184 60700 13190
rect 60646 13152 60648 13161
rect 60700 13152 60702 13161
rect 60646 13087 60702 13096
rect 60556 12844 60608 12850
rect 60556 12786 60608 12792
rect 60384 12406 60504 12434
rect 60004 11892 60056 11898
rect 60004 11834 60056 11840
rect 60016 11354 60044 11834
rect 60096 11824 60148 11830
rect 60096 11766 60148 11772
rect 60108 11558 60136 11766
rect 60384 11626 60412 12406
rect 60648 11756 60700 11762
rect 60752 11744 60780 13262
rect 60844 13025 60872 13262
rect 60830 13016 60886 13025
rect 60830 12951 60886 12960
rect 60844 12850 60872 12951
rect 60832 12844 60884 12850
rect 60832 12786 60884 12792
rect 60936 11898 60964 15200
rect 61384 13796 61436 13802
rect 61384 13738 61436 13744
rect 61108 13252 61160 13258
rect 61108 13194 61160 13200
rect 61016 12776 61068 12782
rect 61016 12718 61068 12724
rect 61028 12374 61056 12718
rect 61016 12368 61068 12374
rect 61016 12310 61068 12316
rect 61028 12238 61056 12310
rect 61016 12232 61068 12238
rect 61016 12174 61068 12180
rect 61028 11898 61056 12174
rect 60924 11892 60976 11898
rect 60924 11834 60976 11840
rect 61016 11892 61068 11898
rect 61016 11834 61068 11840
rect 60752 11716 60964 11744
rect 60648 11698 60700 11704
rect 60660 11642 60688 11698
rect 60372 11620 60424 11626
rect 60660 11614 60780 11642
rect 60372 11562 60424 11568
rect 60096 11552 60148 11558
rect 60096 11494 60148 11500
rect 60556 11552 60608 11558
rect 60556 11494 60608 11500
rect 60117 11452 60425 11461
rect 60117 11450 60123 11452
rect 60179 11450 60203 11452
rect 60259 11450 60283 11452
rect 60339 11450 60363 11452
rect 60419 11450 60425 11452
rect 60179 11398 60181 11450
rect 60361 11398 60363 11450
rect 60117 11396 60123 11398
rect 60179 11396 60203 11398
rect 60259 11396 60283 11398
rect 60339 11396 60363 11398
rect 60419 11396 60425 11398
rect 60117 11387 60425 11396
rect 60004 11348 60056 11354
rect 60004 11290 60056 11296
rect 60004 10668 60056 10674
rect 60004 10610 60056 10616
rect 59820 10192 59872 10198
rect 60016 10169 60044 10610
rect 60117 10364 60425 10373
rect 60117 10362 60123 10364
rect 60179 10362 60203 10364
rect 60259 10362 60283 10364
rect 60339 10362 60363 10364
rect 60419 10362 60425 10364
rect 60179 10310 60181 10362
rect 60361 10310 60363 10362
rect 60117 10308 60123 10310
rect 60179 10308 60203 10310
rect 60259 10308 60283 10310
rect 60339 10308 60363 10310
rect 60419 10308 60425 10310
rect 60117 10299 60425 10308
rect 59820 10134 59872 10140
rect 60002 10160 60058 10169
rect 60002 10095 60058 10104
rect 60464 9920 60516 9926
rect 60464 9862 60516 9868
rect 60476 9761 60504 9862
rect 60462 9752 60518 9761
rect 60462 9687 60518 9696
rect 60004 9580 60056 9586
rect 60004 9522 60056 9528
rect 59820 9172 59872 9178
rect 59820 9114 59872 9120
rect 59728 8832 59780 8838
rect 59728 8774 59780 8780
rect 59740 8430 59768 8774
rect 59832 8498 59860 9114
rect 60016 8634 60044 9522
rect 60117 9276 60425 9285
rect 60117 9274 60123 9276
rect 60179 9274 60203 9276
rect 60259 9274 60283 9276
rect 60339 9274 60363 9276
rect 60419 9274 60425 9276
rect 60179 9222 60181 9274
rect 60361 9222 60363 9274
rect 60117 9220 60123 9222
rect 60179 9220 60203 9222
rect 60259 9220 60283 9222
rect 60339 9220 60363 9222
rect 60419 9220 60425 9222
rect 60117 9211 60425 9220
rect 60004 8628 60056 8634
rect 60004 8570 60056 8576
rect 59820 8492 59872 8498
rect 59820 8434 59872 8440
rect 59728 8424 59780 8430
rect 59728 8366 59780 8372
rect 59544 8084 59596 8090
rect 59544 8026 59596 8032
rect 59556 7954 59584 8026
rect 59544 7948 59596 7954
rect 59544 7890 59596 7896
rect 59084 7880 59136 7886
rect 59084 7822 59136 7828
rect 59268 7812 59320 7818
rect 59268 7754 59320 7760
rect 59176 7540 59228 7546
rect 59176 7482 59228 7488
rect 58992 6860 59044 6866
rect 58992 6802 59044 6808
rect 58808 5228 58860 5234
rect 58808 5170 58860 5176
rect 58532 4072 58584 4078
rect 58532 4014 58584 4020
rect 58544 3602 58572 4014
rect 59188 3670 59216 7482
rect 59176 3664 59228 3670
rect 59176 3606 59228 3612
rect 58532 3596 58584 3602
rect 58532 3538 58584 3544
rect 58716 3596 58768 3602
rect 58716 3538 58768 3544
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 57612 3392 57664 3398
rect 57612 3334 57664 3340
rect 57244 2916 57296 2922
rect 57244 2858 57296 2864
rect 57624 2854 57652 3334
rect 57612 2848 57664 2854
rect 57612 2790 57664 2796
rect 49712 2746 49832 2774
rect 56612 2746 56732 2774
rect 49712 2650 49740 2746
rect 49700 2644 49752 2650
rect 49700 2586 49752 2592
rect 47308 2508 47360 2514
rect 47308 2450 47360 2456
rect 56612 2446 56640 2746
rect 58728 2514 58756 3538
rect 58716 2508 58768 2514
rect 58716 2450 58768 2456
rect 59280 2446 59308 7754
rect 59740 7546 59768 8366
rect 59728 7540 59780 7546
rect 59728 7482 59780 7488
rect 59728 6792 59780 6798
rect 59728 6734 59780 6740
rect 59740 6458 59768 6734
rect 59728 6452 59780 6458
rect 59728 6394 59780 6400
rect 59832 2650 59860 8434
rect 60016 8378 60044 8570
rect 59924 8350 60044 8378
rect 59924 5914 59952 8350
rect 60004 8288 60056 8294
rect 60004 8230 60056 8236
rect 60016 7410 60044 8230
rect 60117 8188 60425 8197
rect 60117 8186 60123 8188
rect 60179 8186 60203 8188
rect 60259 8186 60283 8188
rect 60339 8186 60363 8188
rect 60419 8186 60425 8188
rect 60179 8134 60181 8186
rect 60361 8134 60363 8186
rect 60117 8132 60123 8134
rect 60179 8132 60203 8134
rect 60259 8132 60283 8134
rect 60339 8132 60363 8134
rect 60419 8132 60425 8134
rect 60117 8123 60425 8132
rect 60568 7410 60596 11494
rect 60752 10742 60780 11614
rect 60740 10736 60792 10742
rect 60740 10678 60792 10684
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 60660 10130 60688 10610
rect 60830 10160 60886 10169
rect 60648 10124 60700 10130
rect 60700 10084 60780 10112
rect 60830 10095 60886 10104
rect 60648 10066 60700 10072
rect 60648 9920 60700 9926
rect 60648 9862 60700 9868
rect 60660 9110 60688 9862
rect 60752 9586 60780 10084
rect 60740 9580 60792 9586
rect 60740 9522 60792 9528
rect 60648 9104 60700 9110
rect 60648 9046 60700 9052
rect 60660 8498 60688 9046
rect 60844 8906 60872 10095
rect 60832 8900 60884 8906
rect 60832 8842 60884 8848
rect 60832 8560 60884 8566
rect 60832 8502 60884 8508
rect 60648 8492 60700 8498
rect 60648 8434 60700 8440
rect 60844 7750 60872 8502
rect 60936 7818 60964 11716
rect 61016 11688 61068 11694
rect 61016 11630 61068 11636
rect 61028 11014 61056 11630
rect 61016 11008 61068 11014
rect 61016 10950 61068 10956
rect 61028 9926 61056 10950
rect 61120 10282 61148 13194
rect 61396 12850 61424 13738
rect 61488 12986 61516 15200
rect 61476 12980 61528 12986
rect 61476 12922 61528 12928
rect 61384 12844 61436 12850
rect 61384 12786 61436 12792
rect 61936 12640 61988 12646
rect 61936 12582 61988 12588
rect 61660 12164 61712 12170
rect 61660 12106 61712 12112
rect 61292 11892 61344 11898
rect 61292 11834 61344 11840
rect 61304 11694 61332 11834
rect 61566 11792 61622 11801
rect 61566 11727 61568 11736
rect 61620 11727 61622 11736
rect 61568 11698 61620 11704
rect 61292 11688 61344 11694
rect 61292 11630 61344 11636
rect 61120 10254 61332 10282
rect 61016 9920 61068 9926
rect 61016 9862 61068 9868
rect 61200 9716 61252 9722
rect 61200 9658 61252 9664
rect 61212 8022 61240 9658
rect 61304 8838 61332 10254
rect 61672 9382 61700 12106
rect 61948 11762 61976 12582
rect 61936 11756 61988 11762
rect 61936 11698 61988 11704
rect 62040 11354 62068 15200
rect 62396 12232 62448 12238
rect 62396 12174 62448 12180
rect 62488 12232 62540 12238
rect 62488 12174 62540 12180
rect 62304 11892 62356 11898
rect 62304 11834 62356 11840
rect 62316 11694 62344 11834
rect 62304 11688 62356 11694
rect 62304 11630 62356 11636
rect 62028 11348 62080 11354
rect 62028 11290 62080 11296
rect 62028 11212 62080 11218
rect 62028 11154 62080 11160
rect 62040 11014 62068 11154
rect 62120 11144 62172 11150
rect 62120 11086 62172 11092
rect 62028 11008 62080 11014
rect 62028 10950 62080 10956
rect 62028 10464 62080 10470
rect 62028 10406 62080 10412
rect 62040 10198 62068 10406
rect 62028 10192 62080 10198
rect 62028 10134 62080 10140
rect 62132 9654 62160 11086
rect 62212 10600 62264 10606
rect 62212 10542 62264 10548
rect 62120 9648 62172 9654
rect 62120 9590 62172 9596
rect 61660 9376 61712 9382
rect 61660 9318 61712 9324
rect 61672 8974 61700 9318
rect 62132 9042 62160 9590
rect 62120 9036 62172 9042
rect 62120 8978 62172 8984
rect 61660 8968 61712 8974
rect 61660 8910 61712 8916
rect 61752 8900 61804 8906
rect 61752 8842 61804 8848
rect 61292 8832 61344 8838
rect 61292 8774 61344 8780
rect 61660 8832 61712 8838
rect 61660 8774 61712 8780
rect 61200 8016 61252 8022
rect 61200 7958 61252 7964
rect 61568 7948 61620 7954
rect 61568 7890 61620 7896
rect 60924 7812 60976 7818
rect 60924 7754 60976 7760
rect 60832 7744 60884 7750
rect 60832 7686 60884 7692
rect 60004 7404 60056 7410
rect 60004 7346 60056 7352
rect 60556 7404 60608 7410
rect 60556 7346 60608 7352
rect 60844 7274 60872 7686
rect 61580 7410 61608 7890
rect 61568 7404 61620 7410
rect 61568 7346 61620 7352
rect 60832 7268 60884 7274
rect 60832 7210 60884 7216
rect 61108 7200 61160 7206
rect 61108 7142 61160 7148
rect 60117 7100 60425 7109
rect 60117 7098 60123 7100
rect 60179 7098 60203 7100
rect 60259 7098 60283 7100
rect 60339 7098 60363 7100
rect 60419 7098 60425 7100
rect 60179 7046 60181 7098
rect 60361 7046 60363 7098
rect 60117 7044 60123 7046
rect 60179 7044 60203 7046
rect 60259 7044 60283 7046
rect 60339 7044 60363 7046
rect 60419 7044 60425 7046
rect 60117 7035 60425 7044
rect 60464 6724 60516 6730
rect 60464 6666 60516 6672
rect 60117 6012 60425 6021
rect 60117 6010 60123 6012
rect 60179 6010 60203 6012
rect 60259 6010 60283 6012
rect 60339 6010 60363 6012
rect 60419 6010 60425 6012
rect 60179 5958 60181 6010
rect 60361 5958 60363 6010
rect 60117 5956 60123 5958
rect 60179 5956 60203 5958
rect 60259 5956 60283 5958
rect 60339 5956 60363 5958
rect 60419 5956 60425 5958
rect 60117 5947 60425 5956
rect 59912 5908 59964 5914
rect 59912 5850 59964 5856
rect 60117 4924 60425 4933
rect 60117 4922 60123 4924
rect 60179 4922 60203 4924
rect 60259 4922 60283 4924
rect 60339 4922 60363 4924
rect 60419 4922 60425 4924
rect 60179 4870 60181 4922
rect 60361 4870 60363 4922
rect 60117 4868 60123 4870
rect 60179 4868 60203 4870
rect 60259 4868 60283 4870
rect 60339 4868 60363 4870
rect 60419 4868 60425 4870
rect 60117 4859 60425 4868
rect 60476 3942 60504 6666
rect 61120 5234 61148 7142
rect 61672 6934 61700 8774
rect 61660 6928 61712 6934
rect 61660 6870 61712 6876
rect 61764 5234 61792 8842
rect 62224 8634 62252 10542
rect 62408 10130 62436 12174
rect 62500 10538 62528 12174
rect 62592 11898 62620 15200
rect 62764 12640 62816 12646
rect 62764 12582 62816 12588
rect 62580 11892 62632 11898
rect 62580 11834 62632 11840
rect 62776 11150 62804 12582
rect 63236 12442 63264 15286
rect 63682 15286 63816 15314
rect 63682 15200 63738 15286
rect 63408 13320 63460 13326
rect 63408 13262 63460 13268
rect 63592 13320 63644 13326
rect 63592 13262 63644 13268
rect 63682 13288 63738 13297
rect 63420 12918 63448 13262
rect 63408 12912 63460 12918
rect 63408 12854 63460 12860
rect 63224 12436 63276 12442
rect 63224 12378 63276 12384
rect 62764 11144 62816 11150
rect 62764 11086 62816 11092
rect 63224 11076 63276 11082
rect 63224 11018 63276 11024
rect 62488 10532 62540 10538
rect 62488 10474 62540 10480
rect 62396 10124 62448 10130
rect 62396 10066 62448 10072
rect 62212 8628 62264 8634
rect 62212 8570 62264 8576
rect 62028 5636 62080 5642
rect 62028 5578 62080 5584
rect 61108 5228 61160 5234
rect 61108 5170 61160 5176
rect 61752 5228 61804 5234
rect 61752 5170 61804 5176
rect 60464 3936 60516 3942
rect 60464 3878 60516 3884
rect 60117 3836 60425 3845
rect 60117 3834 60123 3836
rect 60179 3834 60203 3836
rect 60259 3834 60283 3836
rect 60339 3834 60363 3836
rect 60419 3834 60425 3836
rect 60179 3782 60181 3834
rect 60361 3782 60363 3834
rect 60117 3780 60123 3782
rect 60179 3780 60203 3782
rect 60259 3780 60283 3782
rect 60339 3780 60363 3782
rect 60419 3780 60425 3782
rect 60117 3771 60425 3780
rect 62040 3466 62068 5578
rect 62408 5370 62436 10066
rect 63040 10056 63092 10062
rect 63040 9998 63092 10004
rect 62580 9920 62632 9926
rect 62580 9862 62632 9868
rect 62592 9761 62620 9862
rect 62578 9752 62634 9761
rect 63052 9722 63080 9998
rect 62578 9687 62634 9696
rect 63040 9716 63092 9722
rect 63040 9658 63092 9664
rect 62670 8936 62726 8945
rect 62670 8871 62672 8880
rect 62724 8871 62726 8880
rect 62672 8842 62724 8848
rect 62684 8634 62712 8842
rect 62672 8628 62724 8634
rect 62672 8570 62724 8576
rect 62672 7880 62724 7886
rect 62672 7822 62724 7828
rect 62684 7342 62712 7822
rect 63236 7546 63264 11018
rect 63420 11014 63448 12854
rect 63604 11558 63632 13262
rect 63682 13223 63738 13232
rect 63592 11552 63644 11558
rect 63592 11494 63644 11500
rect 63408 11008 63460 11014
rect 63408 10950 63460 10956
rect 63420 10606 63448 10950
rect 63408 10600 63460 10606
rect 63408 10542 63460 10548
rect 63408 9920 63460 9926
rect 63408 9862 63460 9868
rect 63224 7540 63276 7546
rect 63224 7482 63276 7488
rect 63420 7410 63448 9862
rect 63500 9580 63552 9586
rect 63500 9522 63552 9528
rect 63512 9110 63540 9522
rect 63696 9518 63724 13223
rect 63788 12442 63816 15286
rect 63880 15286 64290 15314
rect 63880 12986 63908 15286
rect 64234 15200 64290 15286
rect 64786 15200 64842 16000
rect 65338 15314 65394 16000
rect 65890 15314 65946 16000
rect 65338 15286 65472 15314
rect 65338 15200 65394 15286
rect 64144 13184 64196 13190
rect 64144 13126 64196 13132
rect 63868 12980 63920 12986
rect 63868 12922 63920 12928
rect 64052 12708 64104 12714
rect 64052 12650 64104 12656
rect 63776 12436 63828 12442
rect 63776 12378 63828 12384
rect 63868 11008 63920 11014
rect 63868 10950 63920 10956
rect 63880 10849 63908 10950
rect 63866 10840 63922 10849
rect 63866 10775 63922 10784
rect 63866 10704 63922 10713
rect 63866 10639 63868 10648
rect 63920 10639 63922 10648
rect 63868 10610 63920 10616
rect 63960 9988 64012 9994
rect 63960 9930 64012 9936
rect 63684 9512 63736 9518
rect 63684 9454 63736 9460
rect 63500 9104 63552 9110
rect 63500 9046 63552 9052
rect 63408 7404 63460 7410
rect 63408 7346 63460 7352
rect 62672 7336 62724 7342
rect 62672 7278 62724 7284
rect 63512 6458 63540 9046
rect 63592 8832 63644 8838
rect 63592 8774 63644 8780
rect 63500 6452 63552 6458
rect 63500 6394 63552 6400
rect 63512 6118 63540 6394
rect 63500 6112 63552 6118
rect 63500 6054 63552 6060
rect 63316 5772 63368 5778
rect 63316 5714 63368 5720
rect 63328 5370 63356 5714
rect 62396 5364 62448 5370
rect 62396 5306 62448 5312
rect 63316 5364 63368 5370
rect 63316 5306 63368 5312
rect 63328 4282 63356 5306
rect 63316 4276 63368 4282
rect 63316 4218 63368 4224
rect 62120 4140 62172 4146
rect 62120 4082 62172 4088
rect 62132 3738 62160 4082
rect 62120 3732 62172 3738
rect 62120 3674 62172 3680
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 62040 3058 62068 3402
rect 62028 3052 62080 3058
rect 62028 2994 62080 3000
rect 60117 2748 60425 2757
rect 60117 2746 60123 2748
rect 60179 2746 60203 2748
rect 60259 2746 60283 2748
rect 60339 2746 60363 2748
rect 60419 2746 60425 2748
rect 60179 2694 60181 2746
rect 60361 2694 60363 2746
rect 60117 2692 60123 2694
rect 60179 2692 60203 2694
rect 60259 2692 60283 2694
rect 60339 2692 60363 2694
rect 60419 2692 60425 2694
rect 60117 2683 60425 2692
rect 63328 2650 63356 4218
rect 63512 3738 63540 6054
rect 63604 5302 63632 8774
rect 63696 7002 63724 9454
rect 63776 9376 63828 9382
rect 63776 9318 63828 9324
rect 63684 6996 63736 7002
rect 63684 6938 63736 6944
rect 63788 5710 63816 9318
rect 63972 6186 64000 9930
rect 64064 6458 64092 12650
rect 64156 10674 64184 13126
rect 64420 12844 64472 12850
rect 64420 12786 64472 12792
rect 64236 10736 64288 10742
rect 64236 10678 64288 10684
rect 64144 10668 64196 10674
rect 64144 10610 64196 10616
rect 64248 10266 64276 10678
rect 64236 10260 64288 10266
rect 64236 10202 64288 10208
rect 64248 8566 64276 10202
rect 64432 9926 64460 12786
rect 64800 12442 64828 15200
rect 65156 13252 65208 13258
rect 65156 13194 65208 13200
rect 65168 12918 65196 13194
rect 65444 12986 65472 15286
rect 65890 15286 66116 15314
rect 65890 15200 65946 15286
rect 65524 13932 65576 13938
rect 65524 13874 65576 13880
rect 65536 13326 65564 13874
rect 65892 13796 65944 13802
rect 65892 13738 65944 13744
rect 65904 13462 65932 13738
rect 65892 13456 65944 13462
rect 65892 13398 65944 13404
rect 65524 13320 65576 13326
rect 65524 13262 65576 13268
rect 65616 13320 65668 13326
rect 65668 13280 66024 13308
rect 65616 13262 65668 13268
rect 65996 13190 66024 13280
rect 65892 13184 65944 13190
rect 65892 13126 65944 13132
rect 65984 13184 66036 13190
rect 65984 13126 66036 13132
rect 65432 12980 65484 12986
rect 65432 12922 65484 12928
rect 65156 12912 65208 12918
rect 65156 12854 65208 12860
rect 64788 12436 64840 12442
rect 64788 12378 64840 12384
rect 65800 12232 65852 12238
rect 65800 12174 65852 12180
rect 65708 11756 65760 11762
rect 65628 11716 65708 11744
rect 65628 11558 65656 11716
rect 65708 11698 65760 11704
rect 65064 11552 65116 11558
rect 65064 11494 65116 11500
rect 65616 11552 65668 11558
rect 65616 11494 65668 11500
rect 64512 11144 64564 11150
rect 64512 11086 64564 11092
rect 64420 9920 64472 9926
rect 64420 9862 64472 9868
rect 64236 8560 64288 8566
rect 64236 8502 64288 8508
rect 64248 7478 64276 8502
rect 64236 7472 64288 7478
rect 64236 7414 64288 7420
rect 64524 6798 64552 11086
rect 64788 11076 64840 11082
rect 64788 11018 64840 11024
rect 64604 10464 64656 10470
rect 64604 10406 64656 10412
rect 64696 10464 64748 10470
rect 64696 10406 64748 10412
rect 64616 7410 64644 10406
rect 64708 10062 64736 10406
rect 64696 10056 64748 10062
rect 64696 9998 64748 10004
rect 64800 7546 64828 11018
rect 64972 9716 65024 9722
rect 64972 9658 65024 9664
rect 64984 9586 65012 9658
rect 64880 9580 64932 9586
rect 64880 9522 64932 9528
rect 64972 9580 65024 9586
rect 64972 9522 65024 9528
rect 64892 9178 64920 9522
rect 64984 9178 65012 9522
rect 64880 9172 64932 9178
rect 64880 9114 64932 9120
rect 64972 9172 65024 9178
rect 64972 9114 65024 9120
rect 64984 8022 65012 9114
rect 65076 8838 65104 11494
rect 65248 11212 65300 11218
rect 65248 11154 65300 11160
rect 65260 10130 65288 11154
rect 65812 10538 65840 12174
rect 65904 11642 65932 13126
rect 66088 12986 66116 15286
rect 66442 15200 66498 16000
rect 66994 15200 67050 16000
rect 67546 15200 67602 16000
rect 68098 15200 68154 16000
rect 68650 15200 68706 16000
rect 69202 15200 69258 16000
rect 69754 15200 69810 16000
rect 70306 15314 70362 16000
rect 69952 15286 70362 15314
rect 66456 13530 66484 15200
rect 66628 13728 66680 13734
rect 66628 13670 66680 13676
rect 66640 13530 66668 13670
rect 66444 13524 66496 13530
rect 66444 13466 66496 13472
rect 66628 13524 66680 13530
rect 66628 13466 66680 13472
rect 66904 13252 66956 13258
rect 66904 13194 66956 13200
rect 66076 12980 66128 12986
rect 66076 12922 66128 12928
rect 66916 12918 66944 13194
rect 67008 12986 67036 15200
rect 67560 12986 67588 15200
rect 68112 13530 68140 15200
rect 68100 13524 68152 13530
rect 68100 13466 68152 13472
rect 66996 12980 67048 12986
rect 66996 12922 67048 12928
rect 67548 12980 67600 12986
rect 67548 12922 67600 12928
rect 66904 12912 66956 12918
rect 66904 12854 66956 12860
rect 66260 12844 66312 12850
rect 66812 12844 66864 12850
rect 66312 12804 66484 12832
rect 66260 12786 66312 12792
rect 66166 12744 66222 12753
rect 66456 12714 66484 12804
rect 66812 12786 66864 12792
rect 66166 12679 66222 12688
rect 66444 12708 66496 12714
rect 66180 12374 66208 12679
rect 66444 12650 66496 12656
rect 66168 12368 66220 12374
rect 66168 12310 66220 12316
rect 66824 12102 66852 12786
rect 66916 12782 66944 12854
rect 66904 12776 66956 12782
rect 66904 12718 66956 12724
rect 66168 12096 66220 12102
rect 66168 12038 66220 12044
rect 66812 12096 66864 12102
rect 66812 12038 66864 12044
rect 65904 11614 66024 11642
rect 65892 11552 65944 11558
rect 65892 11494 65944 11500
rect 65800 10532 65852 10538
rect 65800 10474 65852 10480
rect 65248 10124 65300 10130
rect 65248 10066 65300 10072
rect 65260 9722 65288 10066
rect 65248 9716 65300 9722
rect 65248 9658 65300 9664
rect 65260 9058 65288 9658
rect 65800 9376 65852 9382
rect 65800 9318 65852 9324
rect 65168 9030 65288 9058
rect 65064 8832 65116 8838
rect 65064 8774 65116 8780
rect 65168 8634 65196 9030
rect 65812 8974 65840 9318
rect 65904 8974 65932 11494
rect 65248 8968 65300 8974
rect 65248 8910 65300 8916
rect 65800 8968 65852 8974
rect 65800 8910 65852 8916
rect 65892 8968 65944 8974
rect 65892 8910 65944 8916
rect 65156 8628 65208 8634
rect 65156 8570 65208 8576
rect 65260 8294 65288 8910
rect 65892 8356 65944 8362
rect 65892 8298 65944 8304
rect 65248 8288 65300 8294
rect 65248 8230 65300 8236
rect 64972 8016 65024 8022
rect 64972 7958 65024 7964
rect 65260 7886 65288 8230
rect 65904 8022 65932 8298
rect 65892 8016 65944 8022
rect 65892 7958 65944 7964
rect 65248 7880 65300 7886
rect 65248 7822 65300 7828
rect 65260 7546 65288 7822
rect 64788 7540 64840 7546
rect 64788 7482 64840 7488
rect 65248 7540 65300 7546
rect 65248 7482 65300 7488
rect 64604 7404 64656 7410
rect 64604 7346 64656 7352
rect 64420 6792 64472 6798
rect 64420 6734 64472 6740
rect 64512 6792 64564 6798
rect 64512 6734 64564 6740
rect 64432 6458 64460 6734
rect 65996 6474 66024 11614
rect 66076 9920 66128 9926
rect 66076 9862 66128 9868
rect 65904 6458 66024 6474
rect 66088 6458 66116 9862
rect 64052 6452 64104 6458
rect 64052 6394 64104 6400
rect 64420 6452 64472 6458
rect 64420 6394 64472 6400
rect 65892 6452 66024 6458
rect 65944 6446 66024 6452
rect 65892 6394 65944 6400
rect 63960 6180 64012 6186
rect 63960 6122 64012 6128
rect 65996 5794 66024 6446
rect 66076 6452 66128 6458
rect 66076 6394 66128 6400
rect 65904 5778 66024 5794
rect 65892 5772 66024 5778
rect 65944 5766 66024 5772
rect 65892 5714 65944 5720
rect 63776 5704 63828 5710
rect 63776 5646 63828 5652
rect 65800 5568 65852 5574
rect 65800 5510 65852 5516
rect 63592 5296 63644 5302
rect 63592 5238 63644 5244
rect 64880 4072 64932 4078
rect 64880 4014 64932 4020
rect 64892 3738 64920 4014
rect 63500 3732 63552 3738
rect 63500 3674 63552 3680
rect 64604 3732 64656 3738
rect 64604 3674 64656 3680
rect 64880 3732 64932 3738
rect 64880 3674 64932 3680
rect 64616 3058 64644 3674
rect 65812 3534 65840 5510
rect 65904 5370 65932 5714
rect 66088 5710 66116 6394
rect 66076 5704 66128 5710
rect 66076 5646 66128 5652
rect 65892 5364 65944 5370
rect 65892 5306 65944 5312
rect 65800 3528 65852 3534
rect 65800 3470 65852 3476
rect 64604 3052 64656 3058
rect 64604 2994 64656 3000
rect 66088 2774 66116 5646
rect 66180 3398 66208 12038
rect 66720 11280 66772 11286
rect 66720 11222 66772 11228
rect 66732 11082 66760 11222
rect 66720 11076 66772 11082
rect 66720 11018 66772 11024
rect 66260 10464 66312 10470
rect 66260 10406 66312 10412
rect 66272 9450 66300 10406
rect 66732 9994 66760 11018
rect 66720 9988 66772 9994
rect 66720 9930 66772 9936
rect 66916 9654 66944 12718
rect 67640 12640 67692 12646
rect 67640 12582 67692 12588
rect 67180 11824 67232 11830
rect 67180 11766 67232 11772
rect 66996 11212 67048 11218
rect 66996 11154 67048 11160
rect 66904 9648 66956 9654
rect 66904 9590 66956 9596
rect 66260 9444 66312 9450
rect 66260 9386 66312 9392
rect 66720 9376 66772 9382
rect 66720 9318 66772 9324
rect 66732 8090 66760 9318
rect 66720 8084 66772 8090
rect 66720 8026 66772 8032
rect 66916 7886 66944 9590
rect 66904 7880 66956 7886
rect 66904 7822 66956 7828
rect 67008 7410 67036 11154
rect 67192 10606 67220 11766
rect 67180 10600 67232 10606
rect 67180 10542 67232 10548
rect 67192 10130 67220 10542
rect 67180 10124 67232 10130
rect 67180 10066 67232 10072
rect 67652 10033 67680 12582
rect 68664 12442 68692 15200
rect 69216 13530 69244 15200
rect 69204 13524 69256 13530
rect 69204 13466 69256 13472
rect 68836 13320 68888 13326
rect 68836 13262 68888 13268
rect 69664 13320 69716 13326
rect 69664 13262 69716 13268
rect 68652 12436 68704 12442
rect 68652 12378 68704 12384
rect 67916 12300 67968 12306
rect 67916 12242 67968 12248
rect 67730 10976 67786 10985
rect 67730 10911 67786 10920
rect 67638 10024 67694 10033
rect 67638 9959 67694 9968
rect 67744 9926 67772 10911
rect 67824 10464 67876 10470
rect 67824 10406 67876 10412
rect 67836 9926 67864 10406
rect 67732 9920 67784 9926
rect 67732 9862 67784 9868
rect 67824 9920 67876 9926
rect 67824 9862 67876 9868
rect 67638 9752 67694 9761
rect 67638 9687 67694 9696
rect 67456 9580 67508 9586
rect 67456 9522 67508 9528
rect 67468 8634 67496 9522
rect 67456 8628 67508 8634
rect 67456 8570 67508 8576
rect 67652 8498 67680 9687
rect 67640 8492 67692 8498
rect 67640 8434 67692 8440
rect 67088 7812 67140 7818
rect 67088 7754 67140 7760
rect 67100 7546 67128 7754
rect 67088 7540 67140 7546
rect 67088 7482 67140 7488
rect 66996 7404 67048 7410
rect 66996 7346 67048 7352
rect 66536 6792 66588 6798
rect 66536 6734 66588 6740
rect 66260 6656 66312 6662
rect 66260 6598 66312 6604
rect 66272 5710 66300 6598
rect 66548 6458 66576 6734
rect 66628 6724 66680 6730
rect 66628 6666 66680 6672
rect 66536 6452 66588 6458
rect 66536 6394 66588 6400
rect 66640 5914 66668 6666
rect 66628 5908 66680 5914
rect 66628 5850 66680 5856
rect 67652 5846 67680 8434
rect 67836 8430 67864 9862
rect 67824 8424 67876 8430
rect 67824 8366 67876 8372
rect 67928 6662 67956 12242
rect 68848 12170 68876 13262
rect 69676 13161 69704 13262
rect 69662 13152 69718 13161
rect 69662 13087 69718 13096
rect 69480 12844 69532 12850
rect 69480 12786 69532 12792
rect 69112 12368 69164 12374
rect 69112 12310 69164 12316
rect 68836 12164 68888 12170
rect 68836 12106 68888 12112
rect 68744 12096 68796 12102
rect 68744 12038 68796 12044
rect 68560 11756 68612 11762
rect 68560 11698 68612 11704
rect 68376 11552 68428 11558
rect 68376 11494 68428 11500
rect 68388 11150 68416 11494
rect 68572 11150 68600 11698
rect 68756 11558 68784 12038
rect 68744 11552 68796 11558
rect 68744 11494 68796 11500
rect 68376 11144 68428 11150
rect 68376 11086 68428 11092
rect 68560 11144 68612 11150
rect 68560 11086 68612 11092
rect 68756 10470 68784 11494
rect 68376 10464 68428 10470
rect 68376 10406 68428 10412
rect 68744 10464 68796 10470
rect 68744 10406 68796 10412
rect 68388 8838 68416 10406
rect 68848 10198 68876 12106
rect 68928 11688 68980 11694
rect 68928 11630 68980 11636
rect 68940 11014 68968 11630
rect 68928 11008 68980 11014
rect 68928 10950 68980 10956
rect 68928 10668 68980 10674
rect 68928 10610 68980 10616
rect 68836 10192 68888 10198
rect 68836 10134 68888 10140
rect 68376 8832 68428 8838
rect 68376 8774 68428 8780
rect 68388 8430 68416 8774
rect 68376 8424 68428 8430
rect 68376 8366 68428 8372
rect 68388 7206 68416 8366
rect 68940 8090 68968 10610
rect 69020 10124 69072 10130
rect 69020 10066 69072 10072
rect 69032 9178 69060 10066
rect 69020 9172 69072 9178
rect 69020 9114 69072 9120
rect 68928 8084 68980 8090
rect 68928 8026 68980 8032
rect 68376 7200 68428 7206
rect 68376 7142 68428 7148
rect 67916 6656 67968 6662
rect 67916 6598 67968 6604
rect 68388 6322 68416 7142
rect 69124 6866 69152 12310
rect 69296 11076 69348 11082
rect 69296 11018 69348 11024
rect 69308 10742 69336 11018
rect 69296 10736 69348 10742
rect 69296 10678 69348 10684
rect 69112 6860 69164 6866
rect 69112 6802 69164 6808
rect 69124 6458 69152 6802
rect 69112 6452 69164 6458
rect 69112 6394 69164 6400
rect 68928 6384 68980 6390
rect 68928 6326 68980 6332
rect 68376 6316 68428 6322
rect 68376 6258 68428 6264
rect 68940 5914 68968 6326
rect 68928 5908 68980 5914
rect 68928 5850 68980 5856
rect 69124 5846 69152 6394
rect 69308 5914 69336 10678
rect 69492 10130 69520 12786
rect 69768 12442 69796 15200
rect 69952 13530 69980 15286
rect 70306 15200 70362 15286
rect 70858 15200 70914 16000
rect 71410 15314 71466 16000
rect 71332 15286 71466 15314
rect 70872 13530 70900 15200
rect 71332 13530 71360 15286
rect 71410 15200 71466 15286
rect 71962 15314 72018 16000
rect 71962 15286 72096 15314
rect 71962 15200 72018 15286
rect 72068 13530 72096 15286
rect 72514 15200 72570 16000
rect 73066 15314 73122 16000
rect 72804 15286 73122 15314
rect 69940 13524 69992 13530
rect 69940 13466 69992 13472
rect 70860 13524 70912 13530
rect 70860 13466 70912 13472
rect 71320 13524 71372 13530
rect 71320 13466 71372 13472
rect 72056 13524 72108 13530
rect 72056 13466 72108 13472
rect 71136 13320 71188 13326
rect 71136 13262 71188 13268
rect 71688 13320 71740 13326
rect 71688 13262 71740 13268
rect 70952 13252 71004 13258
rect 70952 13194 71004 13200
rect 69940 12776 69992 12782
rect 69940 12718 69992 12724
rect 69756 12436 69808 12442
rect 69756 12378 69808 12384
rect 69952 12374 69980 12718
rect 70964 12434 70992 13194
rect 70964 12406 71084 12434
rect 69940 12368 69992 12374
rect 69940 12310 69992 12316
rect 70952 11892 71004 11898
rect 70952 11834 71004 11840
rect 70964 11694 70992 11834
rect 70952 11688 71004 11694
rect 70952 11630 71004 11636
rect 70216 11620 70268 11626
rect 70216 11562 70268 11568
rect 70228 11354 70256 11562
rect 70308 11552 70360 11558
rect 70308 11494 70360 11500
rect 70584 11552 70636 11558
rect 70584 11494 70636 11500
rect 70216 11348 70268 11354
rect 70216 11290 70268 11296
rect 70320 11218 70348 11494
rect 70596 11354 70624 11494
rect 70584 11348 70636 11354
rect 70584 11290 70636 11296
rect 70308 11212 70360 11218
rect 70308 11154 70360 11160
rect 70032 11144 70084 11150
rect 70032 11086 70084 11092
rect 70044 11014 70072 11086
rect 70032 11008 70084 11014
rect 70032 10950 70084 10956
rect 69480 10124 69532 10130
rect 69480 10066 69532 10072
rect 70044 9926 70072 10950
rect 70492 10668 70544 10674
rect 70492 10610 70544 10616
rect 70504 10169 70532 10610
rect 70490 10160 70546 10169
rect 70490 10095 70546 10104
rect 70032 9920 70084 9926
rect 70032 9862 70084 9868
rect 69756 9104 69808 9110
rect 69756 9046 69808 9052
rect 69768 8634 69796 9046
rect 69848 8900 69900 8906
rect 69848 8842 69900 8848
rect 69860 8634 69888 8842
rect 69756 8628 69808 8634
rect 69756 8570 69808 8576
rect 69848 8628 69900 8634
rect 69848 8570 69900 8576
rect 70216 8492 70268 8498
rect 70216 8434 70268 8440
rect 70228 8401 70256 8434
rect 70214 8392 70270 8401
rect 70214 8327 70270 8336
rect 69296 5908 69348 5914
rect 69296 5850 69348 5856
rect 67640 5840 67692 5846
rect 67640 5782 67692 5788
rect 69112 5840 69164 5846
rect 69112 5782 69164 5788
rect 66260 5704 66312 5710
rect 66260 5646 66312 5652
rect 69124 5642 69152 5782
rect 69112 5636 69164 5642
rect 69112 5578 69164 5584
rect 66260 3936 66312 3942
rect 66260 3878 66312 3884
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 66272 3194 66300 3878
rect 67548 3460 67600 3466
rect 67548 3402 67600 3408
rect 66260 3188 66312 3194
rect 66260 3130 66312 3136
rect 67560 3058 67588 3402
rect 69124 3194 69152 5578
rect 69204 3392 69256 3398
rect 69204 3334 69256 3340
rect 69216 3194 69244 3334
rect 69112 3188 69164 3194
rect 69112 3130 69164 3136
rect 69204 3188 69256 3194
rect 69204 3130 69256 3136
rect 67548 3052 67600 3058
rect 67548 2994 67600 3000
rect 69124 2990 69152 3130
rect 69112 2984 69164 2990
rect 69112 2926 69164 2932
rect 65996 2746 66116 2774
rect 59820 2644 59872 2650
rect 59820 2586 59872 2592
rect 63316 2644 63368 2650
rect 63316 2586 63368 2592
rect 65996 2582 66024 2746
rect 71056 2650 71084 12406
rect 71148 12102 71176 13262
rect 71700 12102 71728 13262
rect 72528 12986 72556 15200
rect 72804 13530 72832 15286
rect 73066 15200 73122 15286
rect 73618 15200 73674 16000
rect 74170 15314 74226 16000
rect 74722 15314 74778 16000
rect 73908 15286 74226 15314
rect 72792 13524 72844 13530
rect 72792 13466 72844 13472
rect 73632 12986 73660 15200
rect 73908 13530 73936 15286
rect 74170 15200 74226 15286
rect 74644 15286 74778 15314
rect 73988 13728 74040 13734
rect 73988 13670 74040 13676
rect 73896 13524 73948 13530
rect 73896 13466 73948 13472
rect 74000 13394 74028 13670
rect 74644 13530 74672 15286
rect 74722 15200 74778 15286
rect 75274 15200 75330 16000
rect 75826 15314 75882 16000
rect 75472 15286 75882 15314
rect 74632 13524 74684 13530
rect 74632 13466 74684 13472
rect 73988 13388 74040 13394
rect 73988 13330 74040 13336
rect 73896 13320 73948 13326
rect 73896 13262 73948 13268
rect 75092 13320 75144 13326
rect 75092 13262 75144 13268
rect 71780 12980 71832 12986
rect 71780 12922 71832 12928
rect 72516 12980 72568 12986
rect 72516 12922 72568 12928
rect 73620 12980 73672 12986
rect 73620 12922 73672 12928
rect 71792 12442 71820 12922
rect 72332 12844 72384 12850
rect 72332 12786 72384 12792
rect 73068 12844 73120 12850
rect 73068 12786 73120 12792
rect 71780 12436 71832 12442
rect 71780 12378 71832 12384
rect 72344 12374 72372 12786
rect 73080 12442 73108 12786
rect 73344 12708 73396 12714
rect 73344 12650 73396 12656
rect 73068 12436 73120 12442
rect 73068 12378 73120 12384
rect 72332 12368 72384 12374
rect 72332 12310 72384 12316
rect 71136 12096 71188 12102
rect 71136 12038 71188 12044
rect 71688 12096 71740 12102
rect 71688 12038 71740 12044
rect 71148 9042 71176 12038
rect 71226 10160 71282 10169
rect 71226 10095 71282 10104
rect 71240 10062 71268 10095
rect 71228 10056 71280 10062
rect 71228 9998 71280 10004
rect 71136 9036 71188 9042
rect 71136 8978 71188 8984
rect 71700 8906 71728 12038
rect 72344 11830 72372 12310
rect 73160 12232 73212 12238
rect 73160 12174 73212 12180
rect 72332 11824 72384 11830
rect 72332 11766 72384 11772
rect 72608 11824 72660 11830
rect 72608 11766 72660 11772
rect 72620 11626 72648 11766
rect 72700 11688 72752 11694
rect 72700 11630 72752 11636
rect 72608 11620 72660 11626
rect 72608 11562 72660 11568
rect 71872 11552 71924 11558
rect 71872 11494 71924 11500
rect 71884 11218 71912 11494
rect 71872 11212 71924 11218
rect 71872 11154 71924 11160
rect 72332 11076 72384 11082
rect 72332 11018 72384 11024
rect 71780 10600 71832 10606
rect 71780 10542 71832 10548
rect 71792 10470 71820 10542
rect 71780 10464 71832 10470
rect 71780 10406 71832 10412
rect 71792 9926 71820 10406
rect 71780 9920 71832 9926
rect 71780 9862 71832 9868
rect 71792 9654 71820 9862
rect 71780 9648 71832 9654
rect 71780 9590 71832 9596
rect 71688 8900 71740 8906
rect 71688 8842 71740 8848
rect 72344 8498 72372 11018
rect 72608 10668 72660 10674
rect 72608 10610 72660 10616
rect 72620 9926 72648 10610
rect 72608 9920 72660 9926
rect 72608 9862 72660 9868
rect 72620 9722 72648 9862
rect 72608 9716 72660 9722
rect 72608 9658 72660 9664
rect 72332 8492 72384 8498
rect 72332 8434 72384 8440
rect 72344 6662 72372 8434
rect 72332 6656 72384 6662
rect 72332 6598 72384 6604
rect 72712 5846 72740 11630
rect 72976 11552 73028 11558
rect 72976 11494 73028 11500
rect 72988 11150 73016 11494
rect 72976 11144 73028 11150
rect 72974 11112 72976 11121
rect 73028 11112 73030 11121
rect 72974 11047 73030 11056
rect 72988 11021 73016 11047
rect 73172 9926 73200 12174
rect 73160 9920 73212 9926
rect 73160 9862 73212 9868
rect 73252 8832 73304 8838
rect 73252 8774 73304 8780
rect 73160 8356 73212 8362
rect 73160 8298 73212 8304
rect 72882 7440 72938 7449
rect 72882 7375 72884 7384
rect 72936 7375 72938 7384
rect 72884 7346 72936 7352
rect 72896 6458 72924 7346
rect 73172 7342 73200 8298
rect 73264 7886 73292 8774
rect 73356 8430 73384 12650
rect 73620 11212 73672 11218
rect 73620 11154 73672 11160
rect 73436 9988 73488 9994
rect 73436 9930 73488 9936
rect 73448 9654 73476 9930
rect 73436 9648 73488 9654
rect 73436 9590 73488 9596
rect 73632 9602 73660 11154
rect 73712 10192 73764 10198
rect 73712 10134 73764 10140
rect 73724 9722 73752 10134
rect 73712 9716 73764 9722
rect 73712 9658 73764 9664
rect 73632 9586 73752 9602
rect 73632 9580 73764 9586
rect 73632 9574 73712 9580
rect 73712 9522 73764 9528
rect 73528 9376 73580 9382
rect 73528 9318 73580 9324
rect 73344 8424 73396 8430
rect 73344 8366 73396 8372
rect 73252 7880 73304 7886
rect 73252 7822 73304 7828
rect 73160 7336 73212 7342
rect 73160 7278 73212 7284
rect 73172 6798 73200 7278
rect 73160 6792 73212 6798
rect 73160 6734 73212 6740
rect 73344 6724 73396 6730
rect 73344 6666 73396 6672
rect 72884 6452 72936 6458
rect 72884 6394 72936 6400
rect 72700 5840 72752 5846
rect 72700 5782 72752 5788
rect 73160 5704 73212 5710
rect 73160 5646 73212 5652
rect 73172 5370 73200 5646
rect 73160 5364 73212 5370
rect 73160 5306 73212 5312
rect 73356 4826 73384 6666
rect 73160 4820 73212 4826
rect 73160 4762 73212 4768
rect 73344 4820 73396 4826
rect 73344 4762 73396 4768
rect 73172 3738 73200 4762
rect 73540 4622 73568 9318
rect 73620 8016 73672 8022
rect 73620 7958 73672 7964
rect 73632 7546 73660 7958
rect 73620 7540 73672 7546
rect 73620 7482 73672 7488
rect 73724 6118 73752 9522
rect 73804 6792 73856 6798
rect 73804 6734 73856 6740
rect 73816 6458 73844 6734
rect 73804 6452 73856 6458
rect 73804 6394 73856 6400
rect 73908 6322 73936 13262
rect 74632 12844 74684 12850
rect 74632 12786 74684 12792
rect 74816 12844 74868 12850
rect 74816 12786 74868 12792
rect 74172 12776 74224 12782
rect 74172 12718 74224 12724
rect 73896 6316 73948 6322
rect 73896 6258 73948 6264
rect 73712 6112 73764 6118
rect 73712 6054 73764 6060
rect 74184 5710 74212 12718
rect 74644 12714 74672 12786
rect 74632 12708 74684 12714
rect 74632 12650 74684 12656
rect 74264 12640 74316 12646
rect 74828 12617 74856 12786
rect 75000 12776 75052 12782
rect 75000 12718 75052 12724
rect 74264 12582 74316 12588
rect 74814 12608 74870 12617
rect 74276 12434 74304 12582
rect 74814 12543 74870 12552
rect 74276 12406 74396 12434
rect 74368 11014 74396 12406
rect 74724 11824 74776 11830
rect 74724 11766 74776 11772
rect 74736 11558 74764 11766
rect 74724 11552 74776 11558
rect 74724 11494 74776 11500
rect 74632 11076 74684 11082
rect 74632 11018 74684 11024
rect 74356 11008 74408 11014
rect 74644 10985 74672 11018
rect 74356 10950 74408 10956
rect 74630 10976 74686 10985
rect 74368 10606 74396 10950
rect 74630 10911 74686 10920
rect 74448 10736 74500 10742
rect 74448 10678 74500 10684
rect 74356 10600 74408 10606
rect 74356 10542 74408 10548
rect 74368 8294 74396 10542
rect 74460 9518 74488 10678
rect 74644 10674 74672 10911
rect 74632 10668 74684 10674
rect 74632 10610 74684 10616
rect 74724 10532 74776 10538
rect 74724 10474 74776 10480
rect 74736 10198 74764 10474
rect 74816 10464 74868 10470
rect 74816 10406 74868 10412
rect 74828 10266 74856 10406
rect 74816 10260 74868 10266
rect 74816 10202 74868 10208
rect 74724 10192 74776 10198
rect 74724 10134 74776 10140
rect 74722 10024 74778 10033
rect 74722 9959 74724 9968
rect 74776 9959 74778 9968
rect 74724 9930 74776 9936
rect 74736 9654 74764 9930
rect 74724 9648 74776 9654
rect 74724 9590 74776 9596
rect 74448 9512 74500 9518
rect 74448 9454 74500 9460
rect 74356 8288 74408 8294
rect 74356 8230 74408 8236
rect 74368 7886 74396 8230
rect 74356 7880 74408 7886
rect 74356 7822 74408 7828
rect 74632 7880 74684 7886
rect 74632 7822 74684 7828
rect 74172 5704 74224 5710
rect 74172 5646 74224 5652
rect 74368 5370 74396 7822
rect 74644 6662 74672 7822
rect 74736 7546 74764 9590
rect 74724 7540 74776 7546
rect 74724 7482 74776 7488
rect 74632 6656 74684 6662
rect 74632 6598 74684 6604
rect 75012 6458 75040 12718
rect 75104 8294 75132 13262
rect 75288 12986 75316 15200
rect 75472 13530 75500 15286
rect 75826 15200 75882 15286
rect 76378 15200 76434 16000
rect 76930 15200 76986 16000
rect 77482 15314 77538 16000
rect 77482 15286 77800 15314
rect 77482 15200 77538 15286
rect 75460 13524 75512 13530
rect 75460 13466 75512 13472
rect 75368 13320 75420 13326
rect 75368 13262 75420 13268
rect 75276 12980 75328 12986
rect 75276 12922 75328 12928
rect 75380 12442 75408 13262
rect 75736 13252 75788 13258
rect 75736 13194 75788 13200
rect 75828 13252 75880 13258
rect 75828 13194 75880 13200
rect 75748 12714 75776 13194
rect 75736 12708 75788 12714
rect 75736 12650 75788 12656
rect 75644 12640 75696 12646
rect 75644 12582 75696 12588
rect 75368 12436 75420 12442
rect 75368 12378 75420 12384
rect 75276 12096 75328 12102
rect 75276 12038 75328 12044
rect 75552 12096 75604 12102
rect 75552 12038 75604 12044
rect 75288 11558 75316 12038
rect 75276 11552 75328 11558
rect 75276 11494 75328 11500
rect 75276 11144 75328 11150
rect 75276 11086 75328 11092
rect 75184 9920 75236 9926
rect 75184 9862 75236 9868
rect 75196 8974 75224 9862
rect 75184 8968 75236 8974
rect 75184 8910 75236 8916
rect 75092 8288 75144 8294
rect 75092 8230 75144 8236
rect 75288 8090 75316 11086
rect 75460 11008 75512 11014
rect 75460 10950 75512 10956
rect 75472 9042 75500 10950
rect 75460 9036 75512 9042
rect 75460 8978 75512 8984
rect 75368 8968 75420 8974
rect 75368 8910 75420 8916
rect 75276 8084 75328 8090
rect 75276 8026 75328 8032
rect 75380 6746 75408 8910
rect 75564 7886 75592 12038
rect 75656 11286 75684 12582
rect 75644 11280 75696 11286
rect 75644 11222 75696 11228
rect 75840 10198 75868 13194
rect 76392 12986 76420 15200
rect 76944 13530 76972 15200
rect 77482 13560 77538 13569
rect 76932 13524 76984 13530
rect 77482 13495 77538 13504
rect 76932 13466 76984 13472
rect 77116 13320 77168 13326
rect 77116 13262 77168 13268
rect 77208 13320 77260 13326
rect 77208 13262 77260 13268
rect 76838 13152 76894 13161
rect 76838 13087 76894 13096
rect 76380 12980 76432 12986
rect 76380 12922 76432 12928
rect 76656 12980 76708 12986
rect 76656 12922 76708 12928
rect 76668 12782 76696 12922
rect 76852 12850 76880 13087
rect 76840 12844 76892 12850
rect 76840 12786 76892 12792
rect 76656 12776 76708 12782
rect 76656 12718 76708 12724
rect 76196 12436 76248 12442
rect 76196 12378 76248 12384
rect 75920 12300 75972 12306
rect 75920 12242 75972 12248
rect 75932 11762 75960 12242
rect 76208 11762 76236 12378
rect 76748 12300 76800 12306
rect 76748 12242 76800 12248
rect 75920 11756 75972 11762
rect 75920 11698 75972 11704
rect 76196 11756 76248 11762
rect 76196 11698 76248 11704
rect 75920 11620 75972 11626
rect 75920 11562 75972 11568
rect 75828 10192 75880 10198
rect 75828 10134 75880 10140
rect 75932 9654 75960 11562
rect 76208 10674 76236 11698
rect 76760 11150 76788 12242
rect 76748 11144 76800 11150
rect 76748 11086 76800 11092
rect 76760 10674 76788 11086
rect 77128 11014 77156 13262
rect 77220 12986 77248 13262
rect 77390 13016 77446 13025
rect 77208 12980 77260 12986
rect 77390 12951 77392 12960
rect 77208 12922 77260 12928
rect 77444 12951 77446 12960
rect 77392 12922 77444 12928
rect 77392 12844 77444 12850
rect 77392 12786 77444 12792
rect 77300 12776 77352 12782
rect 77300 12718 77352 12724
rect 77312 12481 77340 12718
rect 77298 12472 77354 12481
rect 77298 12407 77354 12416
rect 77404 12306 77432 12786
rect 77496 12646 77524 13495
rect 77576 13184 77628 13190
rect 77576 13126 77628 13132
rect 77588 12918 77616 13126
rect 77772 12986 77800 15286
rect 78034 15200 78090 16000
rect 78586 15314 78642 16000
rect 78586 15286 78812 15314
rect 78586 15200 78642 15286
rect 78048 13530 78076 15200
rect 78036 13524 78088 13530
rect 78036 13466 78088 13472
rect 78784 12986 78812 15286
rect 79138 15200 79194 16000
rect 79690 15314 79746 16000
rect 79690 15286 79824 15314
rect 79690 15200 79746 15286
rect 79152 13530 79180 15200
rect 79796 13530 79824 15286
rect 80242 15200 80298 16000
rect 80794 15200 80850 16000
rect 81346 15200 81402 16000
rect 81898 15200 81954 16000
rect 82450 15200 82506 16000
rect 83002 15200 83058 16000
rect 83554 15200 83610 16000
rect 84106 15200 84162 16000
rect 84658 15200 84714 16000
rect 85210 15200 85266 16000
rect 85762 15200 85818 16000
rect 86314 15314 86370 16000
rect 86314 15286 86632 15314
rect 86314 15200 86370 15286
rect 80256 13530 80284 15200
rect 80612 13864 80664 13870
rect 80612 13806 80664 13812
rect 79140 13524 79192 13530
rect 79140 13466 79192 13472
rect 79784 13524 79836 13530
rect 79784 13466 79836 13472
rect 80244 13524 80296 13530
rect 80244 13466 80296 13472
rect 79968 13388 80020 13394
rect 79968 13330 80020 13336
rect 79140 13320 79192 13326
rect 79980 13297 80008 13330
rect 79140 13262 79192 13268
rect 79966 13288 80022 13297
rect 77760 12980 77812 12986
rect 77760 12922 77812 12928
rect 78772 12980 78824 12986
rect 78772 12922 78824 12928
rect 77576 12912 77628 12918
rect 77576 12854 77628 12860
rect 78956 12844 79008 12850
rect 78956 12786 79008 12792
rect 77484 12640 77536 12646
rect 77484 12582 77536 12588
rect 77484 12436 77536 12442
rect 77484 12378 77536 12384
rect 77760 12436 77812 12442
rect 77760 12378 77812 12384
rect 77392 12300 77444 12306
rect 77392 12242 77444 12248
rect 77298 12200 77354 12209
rect 77298 12135 77300 12144
rect 77352 12135 77354 12144
rect 77300 12106 77352 12112
rect 77312 11762 77340 12106
rect 77496 12102 77524 12378
rect 77772 12306 77800 12378
rect 78586 12336 78642 12345
rect 77760 12300 77812 12306
rect 78586 12271 78642 12280
rect 77760 12242 77812 12248
rect 78600 12238 78628 12271
rect 78588 12232 78640 12238
rect 78588 12174 78640 12180
rect 77484 12096 77536 12102
rect 77484 12038 77536 12044
rect 78968 11898 78996 12786
rect 79152 12102 79180 13262
rect 79966 13223 80022 13232
rect 80242 13152 80298 13161
rect 79839 13084 80147 13093
rect 80242 13087 80298 13096
rect 79839 13082 79845 13084
rect 79901 13082 79925 13084
rect 79981 13082 80005 13084
rect 80061 13082 80085 13084
rect 80141 13082 80147 13084
rect 79901 13030 79903 13082
rect 80083 13030 80085 13082
rect 79839 13028 79845 13030
rect 79901 13028 79925 13030
rect 79981 13028 80005 13030
rect 80061 13028 80085 13030
rect 80141 13028 80147 13030
rect 79506 13016 79562 13025
rect 79839 13019 80147 13028
rect 80256 12986 80284 13087
rect 79506 12951 79508 12960
rect 79560 12951 79562 12960
rect 80244 12980 80296 12986
rect 79508 12922 79560 12928
rect 80244 12922 80296 12928
rect 80520 12708 80572 12714
rect 80520 12650 80572 12656
rect 80244 12640 80296 12646
rect 80244 12582 80296 12588
rect 80256 12481 80284 12582
rect 80242 12472 80298 12481
rect 80242 12407 80298 12416
rect 79692 12368 79744 12374
rect 79692 12310 79744 12316
rect 79140 12096 79192 12102
rect 79140 12038 79192 12044
rect 78956 11892 79008 11898
rect 78956 11834 79008 11840
rect 78772 11824 78824 11830
rect 78772 11766 78824 11772
rect 77300 11756 77352 11762
rect 77300 11698 77352 11704
rect 78680 11688 78732 11694
rect 78784 11665 78812 11766
rect 78680 11630 78732 11636
rect 78770 11656 78826 11665
rect 77944 11552 77996 11558
rect 77944 11494 77996 11500
rect 77956 11218 77984 11494
rect 77944 11212 77996 11218
rect 77944 11154 77996 11160
rect 77300 11076 77352 11082
rect 77300 11018 77352 11024
rect 77116 11008 77168 11014
rect 77116 10950 77168 10956
rect 76196 10668 76248 10674
rect 76196 10610 76248 10616
rect 76472 10668 76524 10674
rect 76472 10610 76524 10616
rect 76748 10668 76800 10674
rect 76748 10610 76800 10616
rect 76380 10464 76432 10470
rect 76380 10406 76432 10412
rect 76392 10062 76420 10406
rect 76380 10056 76432 10062
rect 76380 9998 76432 10004
rect 75920 9648 75972 9654
rect 75920 9590 75972 9596
rect 75932 9178 75960 9590
rect 75920 9172 75972 9178
rect 75920 9114 75972 9120
rect 76024 8894 76420 8922
rect 76024 8838 76052 8894
rect 76392 8838 76420 8894
rect 76012 8832 76064 8838
rect 76012 8774 76064 8780
rect 76288 8832 76340 8838
rect 76288 8774 76340 8780
rect 76380 8832 76432 8838
rect 76380 8774 76432 8780
rect 76300 7886 76328 8774
rect 76484 8498 76512 10610
rect 76656 10056 76708 10062
rect 76656 9998 76708 10004
rect 76564 9920 76616 9926
rect 76564 9862 76616 9868
rect 76576 9518 76604 9862
rect 76668 9654 76696 9998
rect 76656 9648 76708 9654
rect 76656 9590 76708 9596
rect 76564 9512 76616 9518
rect 76564 9454 76616 9460
rect 76576 8498 76604 9454
rect 76668 8974 76696 9590
rect 77312 9450 77340 11018
rect 77852 10668 77904 10674
rect 77852 10610 77904 10616
rect 77864 9926 77892 10610
rect 77852 9920 77904 9926
rect 77852 9862 77904 9868
rect 77864 9625 77892 9862
rect 77850 9616 77906 9625
rect 77850 9551 77906 9560
rect 78692 9450 78720 11630
rect 78770 11591 78826 11600
rect 79140 11620 79192 11626
rect 79140 11562 79192 11568
rect 78864 11144 78916 11150
rect 78864 11086 78916 11092
rect 78876 10606 78904 11086
rect 79152 10742 79180 11562
rect 78956 10736 79008 10742
rect 78956 10678 79008 10684
rect 79140 10736 79192 10742
rect 79140 10678 79192 10684
rect 78864 10600 78916 10606
rect 78864 10542 78916 10548
rect 77300 9444 77352 9450
rect 77300 9386 77352 9392
rect 78680 9444 78732 9450
rect 78680 9386 78732 9392
rect 76656 8968 76708 8974
rect 76656 8910 76708 8916
rect 76472 8492 76524 8498
rect 76472 8434 76524 8440
rect 76564 8492 76616 8498
rect 76564 8434 76616 8440
rect 75552 7880 75604 7886
rect 75552 7822 75604 7828
rect 76288 7880 76340 7886
rect 76288 7822 76340 7828
rect 75552 7744 75604 7750
rect 75552 7686 75604 7692
rect 76012 7744 76064 7750
rect 76012 7686 76064 7692
rect 75196 6730 75408 6746
rect 75184 6724 75408 6730
rect 75236 6718 75408 6724
rect 75184 6666 75236 6672
rect 75092 6656 75144 6662
rect 75092 6598 75144 6604
rect 75000 6452 75052 6458
rect 75000 6394 75052 6400
rect 75104 6322 75132 6598
rect 75092 6316 75144 6322
rect 75092 6258 75144 6264
rect 74448 5636 74500 5642
rect 74448 5578 74500 5584
rect 74356 5364 74408 5370
rect 74356 5306 74408 5312
rect 73528 4616 73580 4622
rect 73528 4558 73580 4564
rect 73160 3732 73212 3738
rect 73160 3674 73212 3680
rect 74460 3466 74488 5578
rect 75380 5574 75408 6718
rect 75368 5568 75420 5574
rect 75368 5510 75420 5516
rect 74816 5228 74868 5234
rect 74816 5170 74868 5176
rect 74828 3942 74856 5170
rect 75564 5166 75592 7686
rect 75920 7336 75972 7342
rect 75920 7278 75972 7284
rect 75932 6798 75960 7278
rect 75920 6792 75972 6798
rect 75920 6734 75972 6740
rect 75932 6066 75960 6734
rect 76024 6730 76052 7686
rect 76012 6724 76064 6730
rect 76012 6666 76064 6672
rect 76484 6254 76512 8434
rect 76576 8090 76604 8434
rect 78864 8356 78916 8362
rect 78864 8298 78916 8304
rect 76564 8084 76616 8090
rect 76564 8026 76616 8032
rect 78876 6458 78904 8298
rect 78864 6452 78916 6458
rect 78864 6394 78916 6400
rect 76472 6248 76524 6254
rect 76472 6190 76524 6196
rect 77116 6248 77168 6254
rect 77116 6190 77168 6196
rect 75932 6038 76052 6066
rect 75920 5908 75972 5914
rect 75920 5850 75972 5856
rect 75932 5370 75960 5850
rect 76024 5778 76052 6038
rect 76748 5908 76800 5914
rect 76748 5850 76800 5856
rect 76012 5772 76064 5778
rect 76012 5714 76064 5720
rect 76024 5574 76052 5714
rect 76760 5710 76788 5850
rect 76748 5704 76800 5710
rect 76748 5646 76800 5652
rect 76012 5568 76064 5574
rect 76012 5510 76064 5516
rect 75920 5364 75972 5370
rect 75920 5306 75972 5312
rect 76024 5302 76052 5510
rect 76012 5296 76064 5302
rect 76012 5238 76064 5244
rect 75552 5160 75604 5166
rect 75552 5102 75604 5108
rect 74816 3936 74868 3942
rect 74816 3878 74868 3884
rect 74540 3528 74592 3534
rect 74828 3505 74856 3878
rect 74540 3470 74592 3476
rect 74814 3496 74870 3505
rect 74448 3460 74500 3466
rect 74448 3402 74500 3408
rect 74552 2990 74580 3470
rect 74814 3431 74870 3440
rect 74540 2984 74592 2990
rect 74540 2926 74592 2932
rect 71044 2644 71096 2650
rect 71044 2586 71096 2592
rect 65984 2576 66036 2582
rect 65984 2518 66036 2524
rect 74552 2446 74580 2926
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 59268 2440 59320 2446
rect 59268 2382 59320 2388
rect 74540 2440 74592 2446
rect 75564 2394 75592 5102
rect 76024 4078 76052 5238
rect 76378 4584 76434 4593
rect 76378 4519 76380 4528
rect 76432 4519 76434 4528
rect 76380 4490 76432 4496
rect 76392 4146 76420 4490
rect 76380 4140 76432 4146
rect 76380 4082 76432 4088
rect 76012 4072 76064 4078
rect 76012 4014 76064 4020
rect 77128 3738 77156 6190
rect 78876 5710 78904 6394
rect 78864 5704 78916 5710
rect 78864 5646 78916 5652
rect 77208 5636 77260 5642
rect 77208 5578 77260 5584
rect 77220 5098 77248 5578
rect 77208 5092 77260 5098
rect 77208 5034 77260 5040
rect 78968 4146 78996 10678
rect 79704 10606 79732 12310
rect 79839 11996 80147 12005
rect 79839 11994 79845 11996
rect 79901 11994 79925 11996
rect 79981 11994 80005 11996
rect 80061 11994 80085 11996
rect 80141 11994 80147 11996
rect 79901 11942 79903 11994
rect 80083 11942 80085 11994
rect 79839 11940 79845 11942
rect 79901 11940 79925 11942
rect 79981 11940 80005 11942
rect 80061 11940 80085 11942
rect 80141 11940 80147 11942
rect 79839 11931 80147 11940
rect 79839 10908 80147 10917
rect 79839 10906 79845 10908
rect 79901 10906 79925 10908
rect 79981 10906 80005 10908
rect 80061 10906 80085 10908
rect 80141 10906 80147 10908
rect 79901 10854 79903 10906
rect 80083 10854 80085 10906
rect 79839 10852 79845 10854
rect 79901 10852 79925 10854
rect 79981 10852 80005 10854
rect 80061 10852 80085 10854
rect 80141 10852 80147 10854
rect 79839 10843 80147 10852
rect 79876 10736 79928 10742
rect 79874 10704 79876 10713
rect 79928 10704 79930 10713
rect 79874 10639 79930 10648
rect 79692 10600 79744 10606
rect 79692 10542 79744 10548
rect 79600 9988 79652 9994
rect 79600 9930 79652 9936
rect 79612 9382 79640 9930
rect 79704 9586 79732 10542
rect 79839 9820 80147 9829
rect 79839 9818 79845 9820
rect 79901 9818 79925 9820
rect 79981 9818 80005 9820
rect 80061 9818 80085 9820
rect 80141 9818 80147 9820
rect 79901 9766 79903 9818
rect 80083 9766 80085 9818
rect 79839 9764 79845 9766
rect 79901 9764 79925 9766
rect 79981 9764 80005 9766
rect 80061 9764 80085 9766
rect 80141 9764 80147 9766
rect 79839 9755 80147 9764
rect 79876 9648 79928 9654
rect 79876 9590 79928 9596
rect 79692 9580 79744 9586
rect 79692 9522 79744 9528
rect 79600 9376 79652 9382
rect 79600 9318 79652 9324
rect 79888 9058 79916 9590
rect 79968 9444 80020 9450
rect 79968 9386 80020 9392
rect 79704 9042 79916 9058
rect 79692 9036 79916 9042
rect 79744 9030 79916 9036
rect 79692 8978 79744 8984
rect 79980 8906 80008 9386
rect 79968 8900 80020 8906
rect 79968 8842 80020 8848
rect 79839 8732 80147 8741
rect 79839 8730 79845 8732
rect 79901 8730 79925 8732
rect 79981 8730 80005 8732
rect 80061 8730 80085 8732
rect 80141 8730 80147 8732
rect 79901 8678 79903 8730
rect 80083 8678 80085 8730
rect 79839 8676 79845 8678
rect 79901 8676 79925 8678
rect 79981 8676 80005 8678
rect 80061 8676 80085 8678
rect 80141 8676 80147 8678
rect 79839 8667 80147 8676
rect 79839 7644 80147 7653
rect 79839 7642 79845 7644
rect 79901 7642 79925 7644
rect 79981 7642 80005 7644
rect 80061 7642 80085 7644
rect 80141 7642 80147 7644
rect 79901 7590 79903 7642
rect 80083 7590 80085 7642
rect 79839 7588 79845 7590
rect 79901 7588 79925 7590
rect 79981 7588 80005 7590
rect 80061 7588 80085 7590
rect 80141 7588 80147 7590
rect 79839 7579 80147 7588
rect 79048 7336 79100 7342
rect 79048 7278 79100 7284
rect 79060 6798 79088 7278
rect 79048 6792 79100 6798
rect 79048 6734 79100 6740
rect 79140 6792 79192 6798
rect 79140 6734 79192 6740
rect 79152 6186 79180 6734
rect 79324 6656 79376 6662
rect 79324 6598 79376 6604
rect 79336 6458 79364 6598
rect 79839 6556 80147 6565
rect 79839 6554 79845 6556
rect 79901 6554 79925 6556
rect 79981 6554 80005 6556
rect 80061 6554 80085 6556
rect 80141 6554 80147 6556
rect 79901 6502 79903 6554
rect 80083 6502 80085 6554
rect 79839 6500 79845 6502
rect 79901 6500 79925 6502
rect 79981 6500 80005 6502
rect 80061 6500 80085 6502
rect 80141 6500 80147 6502
rect 79839 6491 80147 6500
rect 79324 6452 79376 6458
rect 79324 6394 79376 6400
rect 79140 6180 79192 6186
rect 79140 6122 79192 6128
rect 79839 5468 80147 5477
rect 79839 5466 79845 5468
rect 79901 5466 79925 5468
rect 79981 5466 80005 5468
rect 80061 5466 80085 5468
rect 80141 5466 80147 5468
rect 79901 5414 79903 5466
rect 80083 5414 80085 5466
rect 79839 5412 79845 5414
rect 79901 5412 79925 5414
rect 79981 5412 80005 5414
rect 80061 5412 80085 5414
rect 80141 5412 80147 5414
rect 79839 5403 80147 5412
rect 79839 4380 80147 4389
rect 79839 4378 79845 4380
rect 79901 4378 79925 4380
rect 79981 4378 80005 4380
rect 80061 4378 80085 4380
rect 80141 4378 80147 4380
rect 79901 4326 79903 4378
rect 80083 4326 80085 4378
rect 79839 4324 79845 4326
rect 79901 4324 79925 4326
rect 79981 4324 80005 4326
rect 80061 4324 80085 4326
rect 80141 4324 80147 4326
rect 79839 4315 80147 4324
rect 78956 4140 79008 4146
rect 78956 4082 79008 4088
rect 77116 3732 77168 3738
rect 77116 3674 77168 3680
rect 80256 3670 80284 12407
rect 80532 12374 80560 12650
rect 80520 12368 80572 12374
rect 80520 12310 80572 12316
rect 80520 12232 80572 12238
rect 80520 12174 80572 12180
rect 80532 11762 80560 12174
rect 80520 11756 80572 11762
rect 80520 11698 80572 11704
rect 80336 8968 80388 8974
rect 80336 8910 80388 8916
rect 80348 8362 80376 8910
rect 80336 8356 80388 8362
rect 80336 8298 80388 8304
rect 80624 8090 80652 13806
rect 80808 13530 80836 15200
rect 80796 13524 80848 13530
rect 80796 13466 80848 13472
rect 81360 13462 81388 15200
rect 81912 13530 81940 15200
rect 82084 13728 82136 13734
rect 82084 13670 82136 13676
rect 82176 13728 82228 13734
rect 82176 13670 82228 13676
rect 81900 13524 81952 13530
rect 81900 13466 81952 13472
rect 81348 13456 81400 13462
rect 81348 13398 81400 13404
rect 81072 13320 81124 13326
rect 81072 13262 81124 13268
rect 81164 13320 81216 13326
rect 81164 13262 81216 13268
rect 81530 13288 81586 13297
rect 80704 12096 80756 12102
rect 80704 12038 80756 12044
rect 80612 8084 80664 8090
rect 80612 8026 80664 8032
rect 80428 7948 80480 7954
rect 80428 7890 80480 7896
rect 80440 7206 80468 7890
rect 80624 7886 80652 8026
rect 80612 7880 80664 7886
rect 80612 7822 80664 7828
rect 80428 7200 80480 7206
rect 80428 7142 80480 7148
rect 80612 6656 80664 6662
rect 80612 6598 80664 6604
rect 80624 6458 80652 6598
rect 80612 6452 80664 6458
rect 80612 6394 80664 6400
rect 80428 6248 80480 6254
rect 80428 6190 80480 6196
rect 80440 5778 80468 6190
rect 80716 6186 80744 12038
rect 81084 10810 81112 13262
rect 81072 10804 81124 10810
rect 81072 10746 81124 10752
rect 81072 7336 81124 7342
rect 81072 7278 81124 7284
rect 81084 6458 81112 7278
rect 81176 6866 81204 13262
rect 81530 13223 81586 13232
rect 81348 12844 81400 12850
rect 81348 12786 81400 12792
rect 81360 12481 81388 12786
rect 81346 12472 81402 12481
rect 81346 12407 81402 12416
rect 81348 11892 81400 11898
rect 81348 11834 81400 11840
rect 81360 11014 81388 11834
rect 81440 11824 81492 11830
rect 81440 11766 81492 11772
rect 81452 11354 81480 11766
rect 81544 11354 81572 13223
rect 82096 12782 82124 13670
rect 82188 13569 82216 13670
rect 82174 13560 82230 13569
rect 82174 13495 82230 13504
rect 82268 13320 82320 13326
rect 82268 13262 82320 13268
rect 82084 12776 82136 12782
rect 82084 12718 82136 12724
rect 81912 12406 82216 12434
rect 81912 12345 81940 12406
rect 82188 12374 82216 12406
rect 82176 12368 82228 12374
rect 81898 12336 81954 12345
rect 81898 12271 81954 12280
rect 82082 12336 82138 12345
rect 82176 12310 82228 12316
rect 82082 12271 82138 12280
rect 82096 12238 82124 12271
rect 81716 12232 81768 12238
rect 81716 12174 81768 12180
rect 82084 12232 82136 12238
rect 82084 12174 82136 12180
rect 81728 12102 81756 12174
rect 81624 12096 81676 12102
rect 81624 12038 81676 12044
rect 81716 12096 81768 12102
rect 81716 12038 81768 12044
rect 81636 11762 81664 12038
rect 81624 11756 81676 11762
rect 81624 11698 81676 11704
rect 81440 11348 81492 11354
rect 81440 11290 81492 11296
rect 81532 11348 81584 11354
rect 81532 11290 81584 11296
rect 81256 11008 81308 11014
rect 81254 10976 81256 10985
rect 81348 11008 81400 11014
rect 81308 10976 81310 10985
rect 81348 10950 81400 10956
rect 81254 10911 81310 10920
rect 81256 10056 81308 10062
rect 81256 9998 81308 10004
rect 81268 9897 81296 9998
rect 81254 9888 81310 9897
rect 81254 9823 81310 9832
rect 81440 9376 81492 9382
rect 81440 9318 81492 9324
rect 81452 7818 81480 9318
rect 81440 7812 81492 7818
rect 81440 7754 81492 7760
rect 81256 7744 81308 7750
rect 81256 7686 81308 7692
rect 81164 6860 81216 6866
rect 81164 6802 81216 6808
rect 81164 6724 81216 6730
rect 81164 6666 81216 6672
rect 81072 6452 81124 6458
rect 81072 6394 81124 6400
rect 81084 6254 81112 6394
rect 81072 6248 81124 6254
rect 81072 6190 81124 6196
rect 80704 6180 80756 6186
rect 80704 6122 80756 6128
rect 80428 5772 80480 5778
rect 80428 5714 80480 5720
rect 81072 5228 81124 5234
rect 81072 5170 81124 5176
rect 81084 4826 81112 5170
rect 81072 4820 81124 4826
rect 81072 4762 81124 4768
rect 80244 3664 80296 3670
rect 80244 3606 80296 3612
rect 76104 3392 76156 3398
rect 76104 3334 76156 3340
rect 76116 3194 76144 3334
rect 79839 3292 80147 3301
rect 79839 3290 79845 3292
rect 79901 3290 79925 3292
rect 79981 3290 80005 3292
rect 80061 3290 80085 3292
rect 80141 3290 80147 3292
rect 79901 3238 79903 3290
rect 80083 3238 80085 3290
rect 79839 3236 79845 3238
rect 79901 3236 79925 3238
rect 79981 3236 80005 3238
rect 80061 3236 80085 3238
rect 80141 3236 80147 3238
rect 79839 3227 80147 3236
rect 81176 3194 81204 6666
rect 81268 5710 81296 7686
rect 81256 5704 81308 5710
rect 81256 5646 81308 5652
rect 81268 5302 81296 5646
rect 81256 5296 81308 5302
rect 81256 5238 81308 5244
rect 76104 3188 76156 3194
rect 76104 3130 76156 3136
rect 81164 3188 81216 3194
rect 81164 3130 81216 3136
rect 81348 3188 81400 3194
rect 81348 3130 81400 3136
rect 81360 2446 81388 3130
rect 81728 2774 81756 12038
rect 81900 10464 81952 10470
rect 81900 10406 81952 10412
rect 81912 9994 81940 10406
rect 81900 9988 81952 9994
rect 81900 9930 81952 9936
rect 82280 9450 82308 13262
rect 82464 12986 82492 15200
rect 83016 13530 83044 15200
rect 83004 13524 83056 13530
rect 83004 13466 83056 13472
rect 83188 13456 83240 13462
rect 83188 13398 83240 13404
rect 82452 12980 82504 12986
rect 82452 12922 82504 12928
rect 83200 12850 83228 13398
rect 83568 12986 83596 15200
rect 84120 13530 84148 15200
rect 84672 13530 84700 15200
rect 84108 13524 84160 13530
rect 84108 13466 84160 13472
rect 84568 13524 84620 13530
rect 84568 13466 84620 13472
rect 84660 13524 84712 13530
rect 84660 13466 84712 13472
rect 84016 13320 84068 13326
rect 84016 13262 84068 13268
rect 84292 13320 84344 13326
rect 84292 13262 84344 13268
rect 84028 12986 84056 13262
rect 83556 12980 83608 12986
rect 83556 12922 83608 12928
rect 84016 12980 84068 12986
rect 84016 12922 84068 12928
rect 83188 12844 83240 12850
rect 83188 12786 83240 12792
rect 84108 12844 84160 12850
rect 84108 12786 84160 12792
rect 82452 12640 82504 12646
rect 82452 12582 82504 12588
rect 82464 12170 82492 12582
rect 83186 12472 83242 12481
rect 84120 12434 84148 12786
rect 83242 12416 83320 12434
rect 83186 12407 83320 12416
rect 83200 12406 83320 12407
rect 83096 12300 83148 12306
rect 83096 12242 83148 12248
rect 82452 12164 82504 12170
rect 82452 12106 82504 12112
rect 82636 12096 82688 12102
rect 82636 12038 82688 12044
rect 82648 11898 82676 12038
rect 82636 11892 82688 11898
rect 82636 11834 82688 11840
rect 82820 11552 82872 11558
rect 82820 11494 82872 11500
rect 82832 11082 82860 11494
rect 82820 11076 82872 11082
rect 82820 11018 82872 11024
rect 82544 10600 82596 10606
rect 82544 10542 82596 10548
rect 83004 10600 83056 10606
rect 83004 10542 83056 10548
rect 82556 10180 82584 10542
rect 82728 10192 82780 10198
rect 82556 10152 82728 10180
rect 82556 9518 82584 10152
rect 82728 10134 82780 10140
rect 82728 9716 82780 9722
rect 82728 9658 82780 9664
rect 82544 9512 82596 9518
rect 82544 9454 82596 9460
rect 82268 9444 82320 9450
rect 82268 9386 82320 9392
rect 82636 9376 82688 9382
rect 82636 9318 82688 9324
rect 82648 9178 82676 9318
rect 82740 9178 82768 9658
rect 83016 9518 83044 10542
rect 83108 10198 83136 12242
rect 83292 12102 83320 12406
rect 84028 12406 84148 12434
rect 83280 12096 83332 12102
rect 83280 12038 83332 12044
rect 83096 10192 83148 10198
rect 83096 10134 83148 10140
rect 83108 9926 83136 10134
rect 83096 9920 83148 9926
rect 83096 9862 83148 9868
rect 83004 9512 83056 9518
rect 83004 9454 83056 9460
rect 82636 9172 82688 9178
rect 82636 9114 82688 9120
rect 82728 9172 82780 9178
rect 82728 9114 82780 9120
rect 83108 8004 83136 9862
rect 83016 7976 83136 8004
rect 82636 7268 82688 7274
rect 82636 7210 82688 7216
rect 82452 7200 82504 7206
rect 82648 7154 82676 7210
rect 82504 7148 82676 7154
rect 82452 7142 82676 7148
rect 82464 7126 82676 7142
rect 83016 6934 83044 7976
rect 83096 7404 83148 7410
rect 83096 7346 83148 7352
rect 83108 7206 83136 7346
rect 83096 7200 83148 7206
rect 83096 7142 83148 7148
rect 83004 6928 83056 6934
rect 83004 6870 83056 6876
rect 82636 6792 82688 6798
rect 82636 6734 82688 6740
rect 82648 6458 82676 6734
rect 82636 6452 82688 6458
rect 82636 6394 82688 6400
rect 83016 5166 83044 6870
rect 83004 5160 83056 5166
rect 83004 5102 83056 5108
rect 81900 5024 81952 5030
rect 81900 4966 81952 4972
rect 81912 4690 81940 4966
rect 81900 4684 81952 4690
rect 81900 4626 81952 4632
rect 83108 3194 83136 7142
rect 83292 5710 83320 12038
rect 83924 11688 83976 11694
rect 83924 11630 83976 11636
rect 83832 11552 83884 11558
rect 83832 11494 83884 11500
rect 83556 11348 83608 11354
rect 83556 11290 83608 11296
rect 83568 11082 83596 11290
rect 83556 11076 83608 11082
rect 83556 11018 83608 11024
rect 83844 10742 83872 11494
rect 83936 11150 83964 11630
rect 83924 11144 83976 11150
rect 83924 11086 83976 11092
rect 83832 10736 83884 10742
rect 83832 10678 83884 10684
rect 83372 10600 83424 10606
rect 83372 10542 83424 10548
rect 83384 8537 83412 10542
rect 83832 10464 83884 10470
rect 83832 10406 83884 10412
rect 83464 9920 83516 9926
rect 83464 9862 83516 9868
rect 83370 8528 83426 8537
rect 83370 8463 83426 8472
rect 83476 7478 83504 9862
rect 83844 8498 83872 10406
rect 84028 10146 84056 12406
rect 84108 12300 84160 12306
rect 84108 12242 84160 12248
rect 84120 11694 84148 12242
rect 84304 12102 84332 13262
rect 84580 13190 84608 13466
rect 84568 13184 84620 13190
rect 84568 13126 84620 13132
rect 84476 12844 84528 12850
rect 84476 12786 84528 12792
rect 84488 12434 84516 12786
rect 84660 12640 84712 12646
rect 84660 12582 84712 12588
rect 84396 12406 84516 12434
rect 84292 12096 84344 12102
rect 84292 12038 84344 12044
rect 84200 11892 84252 11898
rect 84200 11834 84252 11840
rect 84108 11688 84160 11694
rect 84108 11630 84160 11636
rect 84212 11286 84240 11834
rect 84200 11280 84252 11286
rect 84200 11222 84252 11228
rect 84396 10282 84424 12406
rect 84476 12096 84528 12102
rect 84476 12038 84528 12044
rect 84120 10266 84424 10282
rect 84108 10260 84424 10266
rect 84160 10254 84424 10260
rect 84108 10202 84160 10208
rect 84488 10180 84516 12038
rect 84568 11008 84620 11014
rect 84568 10950 84620 10956
rect 84580 10470 84608 10950
rect 84568 10464 84620 10470
rect 84568 10406 84620 10412
rect 84568 10260 84620 10266
rect 84568 10202 84620 10208
rect 84212 10152 84516 10180
rect 84028 10118 84148 10146
rect 83924 9104 83976 9110
rect 83924 9046 83976 9052
rect 83936 8634 83964 9046
rect 84016 8832 84068 8838
rect 84016 8774 84068 8780
rect 84028 8634 84056 8774
rect 83924 8628 83976 8634
rect 83924 8570 83976 8576
rect 84016 8628 84068 8634
rect 84016 8570 84068 8576
rect 83648 8492 83700 8498
rect 83648 8434 83700 8440
rect 83832 8492 83884 8498
rect 83832 8434 83884 8440
rect 83464 7472 83516 7478
rect 83464 7414 83516 7420
rect 83660 7206 83688 8434
rect 84120 8294 84148 10118
rect 84212 9382 84240 10152
rect 84580 10062 84608 10202
rect 84568 10056 84620 10062
rect 84568 9998 84620 10004
rect 84200 9376 84252 9382
rect 84200 9318 84252 9324
rect 84292 9376 84344 9382
rect 84292 9318 84344 9324
rect 84476 9376 84528 9382
rect 84476 9318 84528 9324
rect 84304 8838 84332 9318
rect 84488 9042 84516 9318
rect 84476 9036 84528 9042
rect 84476 8978 84528 8984
rect 84292 8832 84344 8838
rect 84292 8774 84344 8780
rect 83924 8288 83976 8294
rect 83924 8230 83976 8236
rect 84108 8288 84160 8294
rect 84108 8230 84160 8236
rect 83936 8090 83964 8230
rect 83924 8084 83976 8090
rect 83924 8026 83976 8032
rect 84672 7410 84700 12582
rect 85224 12442 85252 15200
rect 85488 13184 85540 13190
rect 85488 13126 85540 13132
rect 85500 12782 85528 13126
rect 85396 12776 85448 12782
rect 85396 12718 85448 12724
rect 85488 12776 85540 12782
rect 85488 12718 85540 12724
rect 84752 12436 84804 12442
rect 84752 12378 84804 12384
rect 85212 12436 85264 12442
rect 85212 12378 85264 12384
rect 84764 12170 84792 12378
rect 85408 12306 85436 12718
rect 85500 12345 85528 12718
rect 85776 12442 85804 15200
rect 86604 12986 86632 15286
rect 86866 15200 86922 16000
rect 87418 15200 87474 16000
rect 87970 15200 88026 16000
rect 88522 15314 88578 16000
rect 88522 15286 88840 15314
rect 88522 15200 88578 15286
rect 86684 13184 86736 13190
rect 86684 13126 86736 13132
rect 86592 12980 86644 12986
rect 86592 12922 86644 12928
rect 85764 12436 85816 12442
rect 85764 12378 85816 12384
rect 85486 12336 85542 12345
rect 85396 12300 85448 12306
rect 85486 12271 85542 12280
rect 85396 12242 85448 12248
rect 86408 12232 86460 12238
rect 86408 12174 86460 12180
rect 84752 12164 84804 12170
rect 84752 12106 84804 12112
rect 86420 11898 86448 12174
rect 86408 11892 86460 11898
rect 86408 11834 86460 11840
rect 86224 11756 86276 11762
rect 86224 11698 86276 11704
rect 84844 11552 84896 11558
rect 84844 11494 84896 11500
rect 84856 11098 84884 11494
rect 86236 11393 86264 11698
rect 86696 11665 86724 13126
rect 86776 12640 86828 12646
rect 86776 12582 86828 12588
rect 86788 11778 86816 12582
rect 86880 11898 86908 15200
rect 87432 12918 87460 15200
rect 87880 13728 87932 13734
rect 87880 13670 87932 13676
rect 87328 12912 87380 12918
rect 87328 12854 87380 12860
rect 87420 12912 87472 12918
rect 87420 12854 87472 12860
rect 87340 12442 87368 12854
rect 87892 12850 87920 13670
rect 87880 12844 87932 12850
rect 87880 12786 87932 12792
rect 87984 12714 88012 15200
rect 88064 13728 88116 13734
rect 88064 13670 88116 13676
rect 88076 13258 88104 13670
rect 88812 13530 88840 15286
rect 89074 15200 89130 16000
rect 89626 15200 89682 16000
rect 90178 15200 90234 16000
rect 90730 15314 90786 16000
rect 90730 15286 91048 15314
rect 90730 15200 90786 15286
rect 88708 13524 88760 13530
rect 88708 13466 88760 13472
rect 88800 13524 88852 13530
rect 88800 13466 88852 13472
rect 88616 13456 88668 13462
rect 88616 13398 88668 13404
rect 88432 13320 88484 13326
rect 88432 13262 88484 13268
rect 88064 13252 88116 13258
rect 88064 13194 88116 13200
rect 88156 12844 88208 12850
rect 88156 12786 88208 12792
rect 87972 12708 88024 12714
rect 87972 12650 88024 12656
rect 87328 12436 87380 12442
rect 87328 12378 87380 12384
rect 87880 12436 87932 12442
rect 87880 12378 87932 12384
rect 86868 11892 86920 11898
rect 86868 11834 86920 11840
rect 87512 11824 87564 11830
rect 86788 11762 86908 11778
rect 87512 11766 87564 11772
rect 86788 11756 86920 11762
rect 86788 11750 86868 11756
rect 86682 11656 86738 11665
rect 86682 11591 86738 11600
rect 86222 11384 86278 11393
rect 86222 11319 86278 11328
rect 86684 11212 86736 11218
rect 86684 11154 86736 11160
rect 84856 11082 85068 11098
rect 84856 11076 85080 11082
rect 84856 11070 85028 11076
rect 84752 11008 84804 11014
rect 84752 10950 84804 10956
rect 84764 10198 84792 10950
rect 84856 10606 84884 11070
rect 85028 11018 85080 11024
rect 84936 11008 84988 11014
rect 84936 10950 84988 10956
rect 84948 10810 84976 10950
rect 86696 10810 86724 11154
rect 84936 10804 84988 10810
rect 84936 10746 84988 10752
rect 86684 10804 86736 10810
rect 86684 10746 86736 10752
rect 84844 10600 84896 10606
rect 84844 10542 84896 10548
rect 85304 10464 85356 10470
rect 85304 10406 85356 10412
rect 84752 10192 84804 10198
rect 84752 10134 84804 10140
rect 84764 10062 84792 10134
rect 84752 10056 84804 10062
rect 84752 9998 84804 10004
rect 84844 9988 84896 9994
rect 84844 9930 84896 9936
rect 84856 9897 84884 9930
rect 84842 9888 84898 9897
rect 84842 9823 84898 9832
rect 84844 9648 84896 9654
rect 85120 9648 85172 9654
rect 84896 9608 85120 9636
rect 84844 9590 84896 9596
rect 85120 9590 85172 9596
rect 85212 9444 85264 9450
rect 85212 9386 85264 9392
rect 85224 8566 85252 9386
rect 85212 8560 85264 8566
rect 85212 8502 85264 8508
rect 85316 7546 85344 10406
rect 86788 10198 86816 11750
rect 86868 11698 86920 11704
rect 86960 11756 87012 11762
rect 86960 11698 87012 11704
rect 86868 11620 86920 11626
rect 86868 11562 86920 11568
rect 86880 11286 86908 11562
rect 86868 11280 86920 11286
rect 86868 11222 86920 11228
rect 86866 10976 86922 10985
rect 86866 10911 86922 10920
rect 86880 10606 86908 10911
rect 86868 10600 86920 10606
rect 86868 10542 86920 10548
rect 86408 10192 86460 10198
rect 86408 10134 86460 10140
rect 86776 10192 86828 10198
rect 86776 10134 86828 10140
rect 85488 10056 85540 10062
rect 85488 9998 85540 10004
rect 85396 9580 85448 9586
rect 85396 9522 85448 9528
rect 85408 9110 85436 9522
rect 85396 9104 85448 9110
rect 85396 9046 85448 9052
rect 85304 7540 85356 7546
rect 85304 7482 85356 7488
rect 84660 7404 84712 7410
rect 84660 7346 84712 7352
rect 83648 7200 83700 7206
rect 83648 7142 83700 7148
rect 85500 6474 85528 9998
rect 86420 8974 86448 10134
rect 86972 10130 87000 11698
rect 87524 11354 87552 11766
rect 87788 11552 87840 11558
rect 87892 11540 87920 12378
rect 88168 12374 88196 12786
rect 88444 12782 88472 13262
rect 88628 13258 88656 13398
rect 88616 13252 88668 13258
rect 88616 13194 88668 13200
rect 88432 12776 88484 12782
rect 88432 12718 88484 12724
rect 88156 12368 88208 12374
rect 88156 12310 88208 12316
rect 88064 12164 88116 12170
rect 88064 12106 88116 12112
rect 87972 11688 88024 11694
rect 87972 11630 88024 11636
rect 87840 11512 87920 11540
rect 87788 11494 87840 11500
rect 87512 11348 87564 11354
rect 87512 11290 87564 11296
rect 87236 10736 87288 10742
rect 87236 10678 87288 10684
rect 87248 10577 87276 10678
rect 87696 10668 87748 10674
rect 87696 10610 87748 10616
rect 87234 10568 87290 10577
rect 87234 10503 87236 10512
rect 87288 10503 87290 10512
rect 87236 10474 87288 10480
rect 86960 10124 87012 10130
rect 86960 10066 87012 10072
rect 87708 9926 87736 10610
rect 87984 10010 88012 11630
rect 88076 11558 88104 12106
rect 88064 11552 88116 11558
rect 88064 11494 88116 11500
rect 88154 11520 88210 11529
rect 88154 11455 88210 11464
rect 87984 9982 88104 10010
rect 87696 9920 87748 9926
rect 87696 9862 87748 9868
rect 87880 9920 87932 9926
rect 87880 9862 87932 9868
rect 87972 9920 88024 9926
rect 87972 9862 88024 9868
rect 87786 9344 87842 9353
rect 87786 9279 87842 9288
rect 86408 8968 86460 8974
rect 86408 8910 86460 8916
rect 86420 7954 86448 8910
rect 86500 8900 86552 8906
rect 86500 8842 86552 8848
rect 86512 8362 86540 8842
rect 87800 8838 87828 9279
rect 87788 8832 87840 8838
rect 87788 8774 87840 8780
rect 87892 8566 87920 9862
rect 87880 8560 87932 8566
rect 87880 8502 87932 8508
rect 86500 8356 86552 8362
rect 86500 8298 86552 8304
rect 87892 7954 87920 8502
rect 86408 7948 86460 7954
rect 86408 7890 86460 7896
rect 87880 7948 87932 7954
rect 87880 7890 87932 7896
rect 87696 7880 87748 7886
rect 87696 7822 87748 7828
rect 85580 7812 85632 7818
rect 85580 7754 85632 7760
rect 85592 7206 85620 7754
rect 86224 7540 86276 7546
rect 86224 7482 86276 7488
rect 86236 7342 86264 7482
rect 86224 7336 86276 7342
rect 86224 7278 86276 7284
rect 87708 7206 87736 7822
rect 85580 7200 85632 7206
rect 85580 7142 85632 7148
rect 86408 7200 86460 7206
rect 86408 7142 86460 7148
rect 86776 7200 86828 7206
rect 86776 7142 86828 7148
rect 87696 7200 87748 7206
rect 87696 7142 87748 7148
rect 86420 6662 86448 7142
rect 86788 6934 86816 7142
rect 86776 6928 86828 6934
rect 86776 6870 86828 6876
rect 86408 6656 86460 6662
rect 86408 6598 86460 6604
rect 85500 6458 85620 6474
rect 85500 6452 85632 6458
rect 85500 6446 85580 6452
rect 85580 6394 85632 6400
rect 85592 6118 85620 6394
rect 85580 6112 85632 6118
rect 85580 6054 85632 6060
rect 86420 5846 86448 6598
rect 86408 5840 86460 5846
rect 86408 5782 86460 5788
rect 83280 5704 83332 5710
rect 83280 5646 83332 5652
rect 84292 5024 84344 5030
rect 84292 4966 84344 4972
rect 84304 4622 84332 4966
rect 87984 4826 88012 9862
rect 88076 5098 88104 9982
rect 88168 9178 88196 11455
rect 88720 11286 88748 13466
rect 88892 13184 88944 13190
rect 88890 13152 88892 13161
rect 88984 13184 89036 13190
rect 88944 13152 88946 13161
rect 88984 13126 89036 13132
rect 88890 13087 88946 13096
rect 88996 12730 89024 13126
rect 88904 12702 89024 12730
rect 88904 12646 88932 12702
rect 88892 12640 88944 12646
rect 88892 12582 88944 12588
rect 88982 12608 89038 12617
rect 88904 12170 88932 12582
rect 88982 12543 89038 12552
rect 88892 12164 88944 12170
rect 88892 12106 88944 12112
rect 88708 11280 88760 11286
rect 88708 11222 88760 11228
rect 88524 11076 88576 11082
rect 88524 11018 88576 11024
rect 88340 10736 88392 10742
rect 88340 10678 88392 10684
rect 88352 10470 88380 10678
rect 88432 10668 88484 10674
rect 88432 10610 88484 10616
rect 88340 10464 88392 10470
rect 88340 10406 88392 10412
rect 88340 9988 88392 9994
rect 88340 9930 88392 9936
rect 88246 9752 88302 9761
rect 88352 9722 88380 9930
rect 88246 9687 88302 9696
rect 88340 9716 88392 9722
rect 88260 9586 88288 9687
rect 88340 9658 88392 9664
rect 88352 9586 88380 9658
rect 88248 9580 88300 9586
rect 88248 9522 88300 9528
rect 88340 9580 88392 9586
rect 88340 9522 88392 9528
rect 88352 9178 88380 9522
rect 88156 9172 88208 9178
rect 88156 9114 88208 9120
rect 88340 9172 88392 9178
rect 88340 9114 88392 9120
rect 88340 8832 88392 8838
rect 88338 8800 88340 8809
rect 88392 8800 88394 8809
rect 88338 8735 88394 8744
rect 88444 8498 88472 10610
rect 88536 10470 88564 11018
rect 88904 10606 88932 12106
rect 88996 11898 89024 12543
rect 89088 12458 89116 15200
rect 89444 13320 89496 13326
rect 89258 13288 89314 13297
rect 89444 13262 89496 13268
rect 89258 13223 89260 13232
rect 89312 13223 89314 13232
rect 89260 13194 89312 13200
rect 89456 12918 89484 13262
rect 89444 12912 89496 12918
rect 89640 12900 89668 15200
rect 89720 13728 89772 13734
rect 89720 13670 89772 13676
rect 89732 13326 89760 13670
rect 89720 13320 89772 13326
rect 89720 13262 89772 13268
rect 89640 12872 89944 12900
rect 89444 12854 89496 12860
rect 89352 12844 89404 12850
rect 89352 12786 89404 12792
rect 89088 12430 89208 12458
rect 89180 12374 89208 12430
rect 89168 12368 89220 12374
rect 89168 12310 89220 12316
rect 89168 12232 89220 12238
rect 89168 12174 89220 12180
rect 88984 11892 89036 11898
rect 88984 11834 89036 11840
rect 89180 10674 89208 12174
rect 89260 11824 89312 11830
rect 89260 11766 89312 11772
rect 89272 11626 89300 11766
rect 89260 11620 89312 11626
rect 89260 11562 89312 11568
rect 89168 10668 89220 10674
rect 89168 10610 89220 10616
rect 88892 10600 88944 10606
rect 88892 10542 88944 10548
rect 88524 10464 88576 10470
rect 88524 10406 88576 10412
rect 88432 8492 88484 8498
rect 88432 8434 88484 8440
rect 88340 6792 88392 6798
rect 88340 6734 88392 6740
rect 88352 5234 88380 6734
rect 88432 6248 88484 6254
rect 88432 6190 88484 6196
rect 88340 5228 88392 5234
rect 88340 5170 88392 5176
rect 88064 5092 88116 5098
rect 88064 5034 88116 5040
rect 88352 4826 88380 5170
rect 87972 4820 88024 4826
rect 87972 4762 88024 4768
rect 88340 4820 88392 4826
rect 88340 4762 88392 4768
rect 84292 4616 84344 4622
rect 84292 4558 84344 4564
rect 84844 3936 84896 3942
rect 84844 3878 84896 3884
rect 84856 3466 84884 3878
rect 88444 3738 88472 6190
rect 88432 3732 88484 3738
rect 88432 3674 88484 3680
rect 84844 3460 84896 3466
rect 84844 3402 84896 3408
rect 83096 3188 83148 3194
rect 83096 3130 83148 3136
rect 88536 2990 88564 10406
rect 89076 9716 89128 9722
rect 89076 9658 89128 9664
rect 89088 9450 89116 9658
rect 89076 9444 89128 9450
rect 89076 9386 89128 9392
rect 89364 8634 89392 12786
rect 89456 12238 89484 12854
rect 89812 12776 89864 12782
rect 89732 12736 89812 12764
rect 89536 12640 89588 12646
rect 89536 12582 89588 12588
rect 89548 12306 89576 12582
rect 89536 12300 89588 12306
rect 89536 12242 89588 12248
rect 89444 12232 89496 12238
rect 89444 12174 89496 12180
rect 89732 11014 89760 12736
rect 89812 12718 89864 12724
rect 89916 12374 89944 12872
rect 89904 12368 89956 12374
rect 89904 12310 89956 12316
rect 90192 12306 90220 15200
rect 90824 13728 90876 13734
rect 90824 13670 90876 13676
rect 90836 13326 90864 13670
rect 91020 13530 91048 15286
rect 91282 15200 91338 16000
rect 91834 15200 91890 16000
rect 92386 15200 92442 16000
rect 92938 15314 92994 16000
rect 92938 15286 93256 15314
rect 92938 15200 92994 15286
rect 91008 13524 91060 13530
rect 91008 13466 91060 13472
rect 91100 13456 91152 13462
rect 91100 13398 91152 13404
rect 90548 13320 90600 13326
rect 90548 13262 90600 13268
rect 90824 13320 90876 13326
rect 90824 13262 90876 13268
rect 90560 12714 90588 13262
rect 90548 12708 90600 12714
rect 90548 12650 90600 12656
rect 90088 12300 90140 12306
rect 90088 12242 90140 12248
rect 90180 12300 90232 12306
rect 90180 12242 90232 12248
rect 89904 12164 89956 12170
rect 89904 12106 89956 12112
rect 89916 11830 89944 12106
rect 89904 11824 89956 11830
rect 89904 11766 89956 11772
rect 90100 11558 90128 12242
rect 90364 12232 90416 12238
rect 90364 12174 90416 12180
rect 89996 11552 90048 11558
rect 89996 11494 90048 11500
rect 90088 11552 90140 11558
rect 90376 11529 90404 12174
rect 90456 11688 90508 11694
rect 90456 11630 90508 11636
rect 90088 11494 90140 11500
rect 90362 11520 90418 11529
rect 90008 11370 90036 11494
rect 90362 11455 90418 11464
rect 90008 11342 90404 11370
rect 90376 11286 90404 11342
rect 90364 11280 90416 11286
rect 90364 11222 90416 11228
rect 90272 11144 90324 11150
rect 90272 11086 90324 11092
rect 89720 11008 89772 11014
rect 89720 10950 89772 10956
rect 89732 10198 89760 10950
rect 90284 10470 90312 11086
rect 90468 10674 90496 11630
rect 90456 10668 90508 10674
rect 90456 10610 90508 10616
rect 90272 10464 90324 10470
rect 90272 10406 90324 10412
rect 89720 10192 89772 10198
rect 89720 10134 89772 10140
rect 89536 10124 89588 10130
rect 89536 10066 89588 10072
rect 89444 8832 89496 8838
rect 89444 8774 89496 8780
rect 89456 8634 89484 8774
rect 89352 8628 89404 8634
rect 89352 8570 89404 8576
rect 89444 8628 89496 8634
rect 89444 8570 89496 8576
rect 88892 8424 88944 8430
rect 88892 8366 88944 8372
rect 88904 4622 88932 8366
rect 89350 7576 89406 7585
rect 89350 7511 89406 7520
rect 89364 7478 89392 7511
rect 89352 7472 89404 7478
rect 89352 7414 89404 7420
rect 89456 6458 89484 8570
rect 89444 6452 89496 6458
rect 89444 6394 89496 6400
rect 89548 6254 89576 10066
rect 90086 9752 90142 9761
rect 90468 9738 90496 10610
rect 90560 10198 90588 12650
rect 90824 12164 90876 12170
rect 90824 12106 90876 12112
rect 90640 11688 90692 11694
rect 90640 11630 90692 11636
rect 90652 11150 90680 11630
rect 90836 11286 90864 12106
rect 90824 11280 90876 11286
rect 90824 11222 90876 11228
rect 90640 11144 90692 11150
rect 90640 11086 90692 11092
rect 90652 11014 90680 11086
rect 90640 11008 90692 11014
rect 90640 10950 90692 10956
rect 90548 10192 90600 10198
rect 90548 10134 90600 10140
rect 90086 9687 90142 9696
rect 90376 9710 90496 9738
rect 90100 9518 90128 9687
rect 90088 9512 90140 9518
rect 90088 9454 90140 9460
rect 89628 9104 89680 9110
rect 89628 9046 89680 9052
rect 89718 9072 89774 9081
rect 89640 8838 89668 9046
rect 89718 9007 89774 9016
rect 89732 8974 89760 9007
rect 89720 8968 89772 8974
rect 89720 8910 89772 8916
rect 89628 8832 89680 8838
rect 89628 8774 89680 8780
rect 90088 8492 90140 8498
rect 90088 8434 90140 8440
rect 90100 8022 90128 8434
rect 90376 8430 90404 9710
rect 90456 9648 90508 9654
rect 90456 9590 90508 9596
rect 90468 9382 90496 9590
rect 90456 9376 90508 9382
rect 90454 9344 90456 9353
rect 90508 9344 90510 9353
rect 90454 9279 90510 9288
rect 90456 8900 90508 8906
rect 90456 8842 90508 8848
rect 90468 8498 90496 8842
rect 90456 8492 90508 8498
rect 90456 8434 90508 8440
rect 90364 8424 90416 8430
rect 90364 8366 90416 8372
rect 90088 8016 90140 8022
rect 90088 7958 90140 7964
rect 89628 7880 89680 7886
rect 89628 7822 89680 7828
rect 89640 6322 89668 7822
rect 89810 7576 89866 7585
rect 89810 7511 89866 7520
rect 89824 7478 89852 7511
rect 89812 7472 89864 7478
rect 89812 7414 89864 7420
rect 90560 6338 90588 10134
rect 90824 9988 90876 9994
rect 90824 9930 90876 9936
rect 90836 9178 90864 9930
rect 91112 9926 91140 13398
rect 91296 13190 91324 15200
rect 91376 13320 91428 13326
rect 91376 13262 91428 13268
rect 91284 13184 91336 13190
rect 91284 13126 91336 13132
rect 91388 12850 91416 13262
rect 91652 12912 91704 12918
rect 91652 12854 91704 12860
rect 91376 12844 91428 12850
rect 91376 12786 91428 12792
rect 91560 12096 91612 12102
rect 91560 12038 91612 12044
rect 91100 9920 91152 9926
rect 91100 9862 91152 9868
rect 90824 9172 90876 9178
rect 90824 9114 90876 9120
rect 90916 9172 90968 9178
rect 90916 9114 90968 9120
rect 90928 9081 90956 9114
rect 90914 9072 90970 9081
rect 90914 9007 90970 9016
rect 90916 8968 90968 8974
rect 90916 8910 90968 8916
rect 90732 8900 90784 8906
rect 90732 8842 90784 8848
rect 90744 8378 90772 8842
rect 90928 8566 90956 8910
rect 91112 8673 91140 9862
rect 91098 8664 91154 8673
rect 91098 8599 91154 8608
rect 90916 8560 90968 8566
rect 90916 8502 90968 8508
rect 91008 8492 91060 8498
rect 91008 8434 91060 8440
rect 90652 8350 90772 8378
rect 90916 8424 90968 8430
rect 90916 8366 90968 8372
rect 90652 8022 90680 8350
rect 90732 8288 90784 8294
rect 90732 8230 90784 8236
rect 90824 8288 90876 8294
rect 90824 8230 90876 8236
rect 90744 8022 90772 8230
rect 90640 8016 90692 8022
rect 90640 7958 90692 7964
rect 90732 8016 90784 8022
rect 90732 7958 90784 7964
rect 90836 7886 90864 8230
rect 90824 7880 90876 7886
rect 90730 7848 90786 7857
rect 90824 7822 90876 7828
rect 90730 7783 90732 7792
rect 90784 7783 90786 7792
rect 90732 7754 90784 7760
rect 90824 7744 90876 7750
rect 90822 7712 90824 7721
rect 90876 7712 90878 7721
rect 90822 7647 90878 7656
rect 90822 7576 90878 7585
rect 90822 7511 90878 7520
rect 90836 7410 90864 7511
rect 90928 7410 90956 8366
rect 91020 7886 91048 8434
rect 91008 7880 91060 7886
rect 91008 7822 91060 7828
rect 90824 7404 90876 7410
rect 90824 7346 90876 7352
rect 90916 7404 90968 7410
rect 90916 7346 90968 7352
rect 89628 6316 89680 6322
rect 90560 6310 90680 6338
rect 89628 6258 89680 6264
rect 89536 6248 89588 6254
rect 89536 6190 89588 6196
rect 90548 6248 90600 6254
rect 90548 6190 90600 6196
rect 88892 4616 88944 4622
rect 88892 4558 88944 4564
rect 90560 3534 90588 6190
rect 90652 5914 90680 6310
rect 90640 5908 90692 5914
rect 90640 5850 90692 5856
rect 91112 5030 91140 8599
rect 91376 7948 91428 7954
rect 91376 7890 91428 7896
rect 91388 7750 91416 7890
rect 91376 7744 91428 7750
rect 91376 7686 91428 7692
rect 91374 7304 91430 7313
rect 91374 7239 91430 7248
rect 91388 7206 91416 7239
rect 91376 7200 91428 7206
rect 91376 7142 91428 7148
rect 91466 6352 91522 6361
rect 91466 6287 91468 6296
rect 91520 6287 91522 6296
rect 91468 6258 91520 6264
rect 91100 5024 91152 5030
rect 91100 4966 91152 4972
rect 91572 3942 91600 12038
rect 91664 10062 91692 12854
rect 91848 12102 91876 15200
rect 92400 12986 92428 15200
rect 93228 13462 93256 15286
rect 93490 15200 93546 16000
rect 94042 15200 94098 16000
rect 94594 15200 94650 16000
rect 95146 15200 95202 16000
rect 95698 15314 95754 16000
rect 95698 15286 96016 15314
rect 95698 15200 95754 15286
rect 93216 13456 93268 13462
rect 93216 13398 93268 13404
rect 92480 13252 92532 13258
rect 92480 13194 92532 13200
rect 92388 12980 92440 12986
rect 92388 12922 92440 12928
rect 92388 12640 92440 12646
rect 92388 12582 92440 12588
rect 91836 12096 91888 12102
rect 91836 12038 91888 12044
rect 92020 11008 92072 11014
rect 92020 10950 92072 10956
rect 92032 10606 92060 10950
rect 92020 10600 92072 10606
rect 92020 10542 92072 10548
rect 92296 10600 92348 10606
rect 92296 10542 92348 10548
rect 91652 10056 91704 10062
rect 91652 9998 91704 10004
rect 92308 9518 92336 10542
rect 92400 9926 92428 12582
rect 92492 12434 92520 13194
rect 93400 12844 93452 12850
rect 93400 12786 93452 12792
rect 93412 12753 93440 12786
rect 93398 12744 93454 12753
rect 93398 12679 93454 12688
rect 93412 12646 93440 12679
rect 93216 12640 93268 12646
rect 93216 12582 93268 12588
rect 93400 12640 93452 12646
rect 93400 12582 93452 12588
rect 93228 12434 93256 12582
rect 92492 12406 92888 12434
rect 92860 11762 92888 12406
rect 93044 12406 93256 12434
rect 93044 12306 93072 12406
rect 93032 12300 93084 12306
rect 93308 12300 93360 12306
rect 93032 12242 93084 12248
rect 93136 12260 93308 12288
rect 93136 12170 93164 12260
rect 93308 12242 93360 12248
rect 93124 12164 93176 12170
rect 93124 12106 93176 12112
rect 93216 12164 93268 12170
rect 93216 12106 93268 12112
rect 92756 11756 92808 11762
rect 92756 11698 92808 11704
rect 92848 11756 92900 11762
rect 92848 11698 92900 11704
rect 92480 11280 92532 11286
rect 92480 11222 92532 11228
rect 92388 9920 92440 9926
rect 92388 9862 92440 9868
rect 92296 9512 92348 9518
rect 92296 9454 92348 9460
rect 92492 8809 92520 11222
rect 92768 10470 92796 11698
rect 92846 11248 92902 11257
rect 92846 11183 92902 11192
rect 92756 10464 92808 10470
rect 92756 10406 92808 10412
rect 92768 9489 92796 10406
rect 92860 10198 92888 11183
rect 93032 11076 93084 11082
rect 93032 11018 93084 11024
rect 93044 10606 93072 11018
rect 93032 10600 93084 10606
rect 93032 10542 93084 10548
rect 92848 10192 92900 10198
rect 92848 10134 92900 10140
rect 92754 9480 92810 9489
rect 92754 9415 92810 9424
rect 92860 9382 92888 10134
rect 92940 9512 92992 9518
rect 92940 9454 92992 9460
rect 92848 9376 92900 9382
rect 92848 9318 92900 9324
rect 92952 9042 92980 9454
rect 92940 9036 92992 9042
rect 92940 8978 92992 8984
rect 92572 8900 92624 8906
rect 92572 8842 92624 8848
rect 92478 8800 92534 8809
rect 92478 8735 92534 8744
rect 92480 8560 92532 8566
rect 92216 8498 92336 8514
rect 92480 8502 92532 8508
rect 91928 8492 91980 8498
rect 91928 8434 91980 8440
rect 92204 8492 92336 8498
rect 92256 8486 92336 8492
rect 92204 8434 92256 8440
rect 91940 8344 91968 8434
rect 92308 8430 92336 8486
rect 92388 8492 92440 8498
rect 92388 8434 92440 8440
rect 92296 8424 92348 8430
rect 92296 8366 92348 8372
rect 92204 8356 92256 8362
rect 91940 8316 92204 8344
rect 92204 8298 92256 8304
rect 92400 8294 92428 8434
rect 92388 8288 92440 8294
rect 92388 8230 92440 8236
rect 92388 7880 92440 7886
rect 92492 7868 92520 8502
rect 92440 7840 92520 7868
rect 92388 7822 92440 7828
rect 92480 7744 92532 7750
rect 92480 7686 92532 7692
rect 92204 6792 92256 6798
rect 92204 6734 92256 6740
rect 91928 6656 91980 6662
rect 91928 6598 91980 6604
rect 91836 6248 91888 6254
rect 91836 6190 91888 6196
rect 91848 5914 91876 6190
rect 91836 5908 91888 5914
rect 91836 5850 91888 5856
rect 91940 4554 91968 6598
rect 92216 6458 92244 6734
rect 92492 6730 92520 7686
rect 92480 6724 92532 6730
rect 92480 6666 92532 6672
rect 92584 6662 92612 8842
rect 92952 8106 92980 8978
rect 92952 8078 93072 8106
rect 92940 8016 92992 8022
rect 92940 7958 92992 7964
rect 92952 7868 92980 7958
rect 93044 7886 93072 8078
rect 92768 7840 92980 7868
rect 93032 7880 93084 7886
rect 92768 7834 92796 7840
rect 92676 7818 92796 7834
rect 93032 7822 93084 7828
rect 92664 7812 92796 7818
rect 92716 7806 92796 7812
rect 92664 7754 92716 7760
rect 92940 7744 92992 7750
rect 93136 7698 93164 12106
rect 93228 11150 93256 12106
rect 93400 11756 93452 11762
rect 93400 11698 93452 11704
rect 93216 11144 93268 11150
rect 93216 11086 93268 11092
rect 93228 10810 93256 11086
rect 93216 10804 93268 10810
rect 93216 10746 93268 10752
rect 93214 10296 93270 10305
rect 93214 10231 93270 10240
rect 93228 10130 93256 10231
rect 93216 10124 93268 10130
rect 93216 10066 93268 10072
rect 93214 8800 93270 8809
rect 93214 8735 93270 8744
rect 92940 7686 92992 7692
rect 92952 7206 92980 7686
rect 93044 7670 93164 7698
rect 92940 7200 92992 7206
rect 92940 7142 92992 7148
rect 92572 6656 92624 6662
rect 92572 6598 92624 6604
rect 92204 6452 92256 6458
rect 92204 6394 92256 6400
rect 92572 5228 92624 5234
rect 92572 5170 92624 5176
rect 92584 4622 92612 5170
rect 92572 4616 92624 4622
rect 92572 4558 92624 4564
rect 91928 4548 91980 4554
rect 91928 4490 91980 4496
rect 93044 4010 93072 7670
rect 93228 7562 93256 8735
rect 93308 8356 93360 8362
rect 93308 8298 93360 8304
rect 93136 7534 93256 7562
rect 93136 6202 93164 7534
rect 93320 6866 93348 8298
rect 93308 6860 93360 6866
rect 93308 6802 93360 6808
rect 93216 6724 93268 6730
rect 93216 6666 93268 6672
rect 93228 6322 93256 6666
rect 93412 6662 93440 11698
rect 93504 11626 93532 15200
rect 94056 13802 94084 15200
rect 94044 13796 94096 13802
rect 94044 13738 94096 13744
rect 94412 13320 94464 13326
rect 94412 13262 94464 13268
rect 94424 13161 94452 13262
rect 94410 13152 94466 13161
rect 94410 13087 94466 13096
rect 94320 12980 94372 12986
rect 94320 12922 94372 12928
rect 94228 12776 94280 12782
rect 94228 12718 94280 12724
rect 93676 12232 93728 12238
rect 93676 12174 93728 12180
rect 93688 11830 93716 12174
rect 93676 11824 93728 11830
rect 93676 11766 93728 11772
rect 93492 11620 93544 11626
rect 93492 11562 93544 11568
rect 93674 11384 93730 11393
rect 93674 11319 93730 11328
rect 93584 10056 93636 10062
rect 93584 9998 93636 10004
rect 93490 7576 93546 7585
rect 93490 7511 93492 7520
rect 93544 7511 93546 7520
rect 93492 7482 93544 7488
rect 93492 7404 93544 7410
rect 93492 7346 93544 7352
rect 93504 7206 93532 7346
rect 93596 7206 93624 9998
rect 93688 8906 93716 11319
rect 94240 11286 94268 12718
rect 94332 12714 94360 12922
rect 94320 12708 94372 12714
rect 94320 12650 94372 12656
rect 94608 11898 94636 15200
rect 94872 13728 94924 13734
rect 94872 13670 94924 13676
rect 94688 12708 94740 12714
rect 94688 12650 94740 12656
rect 94596 11892 94648 11898
rect 94596 11834 94648 11840
rect 94320 11756 94372 11762
rect 94320 11698 94372 11704
rect 94332 11540 94360 11698
rect 94700 11694 94728 12650
rect 94884 12646 94912 13670
rect 95160 13530 95188 15200
rect 95792 13796 95844 13802
rect 95792 13738 95844 13744
rect 95884 13796 95936 13802
rect 95884 13738 95936 13744
rect 95148 13524 95200 13530
rect 95148 13466 95200 13472
rect 95804 13462 95832 13738
rect 95792 13456 95844 13462
rect 95896 13433 95924 13738
rect 95792 13398 95844 13404
rect 95882 13424 95938 13433
rect 95056 13388 95108 13394
rect 95882 13359 95938 13368
rect 95056 13330 95108 13336
rect 95068 13190 95096 13330
rect 95896 13326 95924 13359
rect 95424 13320 95476 13326
rect 95608 13320 95660 13326
rect 95476 13280 95608 13308
rect 95424 13262 95476 13268
rect 95608 13262 95660 13268
rect 95884 13320 95936 13326
rect 95884 13262 95936 13268
rect 95056 13184 95108 13190
rect 95056 13126 95108 13132
rect 95988 12918 96016 15286
rect 96250 15200 96306 16000
rect 96802 15314 96858 16000
rect 97354 15314 97410 16000
rect 96802 15286 97120 15314
rect 96802 15200 96858 15286
rect 95332 12912 95384 12918
rect 95332 12854 95384 12860
rect 95976 12912 96028 12918
rect 95976 12854 96028 12860
rect 95240 12776 95292 12782
rect 95240 12718 95292 12724
rect 94872 12640 94924 12646
rect 94872 12582 94924 12588
rect 94780 12096 94832 12102
rect 94780 12038 94832 12044
rect 94688 11688 94740 11694
rect 94688 11630 94740 11636
rect 94412 11552 94464 11558
rect 94332 11512 94412 11540
rect 94412 11494 94464 11500
rect 94228 11280 94280 11286
rect 94228 11222 94280 11228
rect 94412 11076 94464 11082
rect 94412 11018 94464 11024
rect 94424 10810 94452 11018
rect 94792 11014 94820 12038
rect 95252 11762 95280 12718
rect 95056 11756 95108 11762
rect 95056 11698 95108 11704
rect 95240 11756 95292 11762
rect 95240 11698 95292 11704
rect 95068 11642 95096 11698
rect 95068 11614 95280 11642
rect 94780 11008 94832 11014
rect 94780 10950 94832 10956
rect 94412 10804 94464 10810
rect 94412 10746 94464 10752
rect 94792 10674 94820 10950
rect 94320 10668 94372 10674
rect 94320 10610 94372 10616
rect 94780 10668 94832 10674
rect 94780 10610 94832 10616
rect 93952 10464 94004 10470
rect 93952 10406 94004 10412
rect 93964 9994 93992 10406
rect 93860 9988 93912 9994
rect 93860 9930 93912 9936
rect 93952 9988 94004 9994
rect 93952 9930 94004 9936
rect 93872 9654 93900 9930
rect 93860 9648 93912 9654
rect 93860 9590 93912 9596
rect 93860 9376 93912 9382
rect 93860 9318 93912 9324
rect 93872 9081 93900 9318
rect 93858 9072 93914 9081
rect 93858 9007 93914 9016
rect 93676 8900 93728 8906
rect 93676 8842 93728 8848
rect 93492 7200 93544 7206
rect 93492 7142 93544 7148
rect 93584 7200 93636 7206
rect 93584 7142 93636 7148
rect 93400 6656 93452 6662
rect 93400 6598 93452 6604
rect 93216 6316 93268 6322
rect 93216 6258 93268 6264
rect 93136 6174 93256 6202
rect 93124 6112 93176 6118
rect 93124 6054 93176 6060
rect 93136 5234 93164 6054
rect 93228 5234 93256 6174
rect 93400 5568 93452 5574
rect 93400 5510 93452 5516
rect 93412 5302 93440 5510
rect 93400 5296 93452 5302
rect 93400 5238 93452 5244
rect 93124 5228 93176 5234
rect 93124 5170 93176 5176
rect 93216 5228 93268 5234
rect 93216 5170 93268 5176
rect 93032 4004 93084 4010
rect 93032 3946 93084 3952
rect 91560 3936 91612 3942
rect 91560 3878 91612 3884
rect 90548 3528 90600 3534
rect 90548 3470 90600 3476
rect 93504 3097 93532 7142
rect 93688 4826 93716 8842
rect 93768 7948 93820 7954
rect 93768 7890 93820 7896
rect 93780 7857 93808 7890
rect 93766 7848 93822 7857
rect 93766 7783 93822 7792
rect 93872 7313 93900 9007
rect 93964 7585 93992 9930
rect 94332 8498 94360 10610
rect 94872 10464 94924 10470
rect 94872 10406 94924 10412
rect 94884 10062 94912 10406
rect 94872 10056 94924 10062
rect 94872 9998 94924 10004
rect 94884 9926 94912 9998
rect 94872 9920 94924 9926
rect 94872 9862 94924 9868
rect 94504 9376 94556 9382
rect 94504 9318 94556 9324
rect 94320 8492 94372 8498
rect 94320 8434 94372 8440
rect 94044 8424 94096 8430
rect 94044 8366 94096 8372
rect 94056 7750 94084 8366
rect 94044 7744 94096 7750
rect 94044 7686 94096 7692
rect 93950 7576 94006 7585
rect 93950 7511 94006 7520
rect 93858 7304 93914 7313
rect 93858 7239 93914 7248
rect 94056 6254 94084 7686
rect 94044 6248 94096 6254
rect 94044 6190 94096 6196
rect 94332 6118 94360 8434
rect 94516 6458 94544 9318
rect 95252 9110 95280 11614
rect 95344 10470 95372 12854
rect 95516 12844 95568 12850
rect 95516 12786 95568 12792
rect 95528 10470 95556 12786
rect 96264 12442 96292 15200
rect 96436 14952 96488 14958
rect 96436 14894 96488 14900
rect 96252 12436 96304 12442
rect 96252 12378 96304 12384
rect 96160 12232 96212 12238
rect 96160 12174 96212 12180
rect 96172 11898 96200 12174
rect 96160 11892 96212 11898
rect 96160 11834 96212 11840
rect 96448 11694 96476 14894
rect 97092 13462 97120 15286
rect 97354 15286 97672 15314
rect 97354 15200 97410 15286
rect 97080 13456 97132 13462
rect 97080 13398 97132 13404
rect 96988 13320 97040 13326
rect 96986 13288 96988 13297
rect 97040 13288 97042 13297
rect 96620 13252 96672 13258
rect 96620 13194 96672 13200
rect 96896 13252 96948 13258
rect 96986 13223 97042 13232
rect 96896 13194 96948 13200
rect 96528 12096 96580 12102
rect 96528 12038 96580 12044
rect 96436 11688 96488 11694
rect 96436 11630 96488 11636
rect 96448 11286 96476 11630
rect 95608 11280 95660 11286
rect 95608 11222 95660 11228
rect 96436 11280 96488 11286
rect 96436 11222 96488 11228
rect 95332 10464 95384 10470
rect 95516 10464 95568 10470
rect 95384 10424 95464 10452
rect 95332 10406 95384 10412
rect 95330 9888 95386 9897
rect 95330 9823 95386 9832
rect 95240 9104 95292 9110
rect 95240 9046 95292 9052
rect 95344 8945 95372 9823
rect 95436 9722 95464 10424
rect 95516 10406 95568 10412
rect 95528 10305 95556 10406
rect 95514 10296 95570 10305
rect 95514 10231 95570 10240
rect 95424 9716 95476 9722
rect 95424 9658 95476 9664
rect 95528 9042 95556 10231
rect 95516 9036 95568 9042
rect 95516 8978 95568 8984
rect 95330 8936 95386 8945
rect 95330 8871 95386 8880
rect 95424 8900 95476 8906
rect 95424 8842 95476 8848
rect 95056 8832 95108 8838
rect 95056 8774 95108 8780
rect 95068 7750 95096 8774
rect 95436 8362 95464 8842
rect 95332 8356 95384 8362
rect 95332 8298 95384 8304
rect 95424 8356 95476 8362
rect 95424 8298 95476 8304
rect 95344 7886 95372 8298
rect 95332 7880 95384 7886
rect 95332 7822 95384 7828
rect 95056 7744 95108 7750
rect 95148 7744 95200 7750
rect 95056 7686 95108 7692
rect 95146 7712 95148 7721
rect 95200 7712 95202 7721
rect 95146 7647 95202 7656
rect 94504 6452 94556 6458
rect 94504 6394 94556 6400
rect 93860 6112 93912 6118
rect 93860 6054 93912 6060
rect 94320 6112 94372 6118
rect 94320 6054 94372 6060
rect 93872 5930 93900 6054
rect 93780 5902 93900 5930
rect 93780 5658 93808 5902
rect 93860 5840 93912 5846
rect 93912 5788 94084 5794
rect 93860 5782 94084 5788
rect 93872 5766 94084 5782
rect 93780 5630 93900 5658
rect 93872 5574 93900 5630
rect 94056 5574 94084 5766
rect 94136 5636 94188 5642
rect 94136 5578 94188 5584
rect 93860 5568 93912 5574
rect 93860 5510 93912 5516
rect 94044 5568 94096 5574
rect 94044 5510 94096 5516
rect 94148 5098 94176 5578
rect 94136 5092 94188 5098
rect 94136 5034 94188 5040
rect 93676 4820 93728 4826
rect 93676 4762 93728 4768
rect 94516 3738 94544 6394
rect 95332 5704 95384 5710
rect 95332 5646 95384 5652
rect 95344 5302 95372 5646
rect 95332 5296 95384 5302
rect 95332 5238 95384 5244
rect 95344 4826 95372 5238
rect 95332 4820 95384 4826
rect 95332 4762 95384 4768
rect 94504 3732 94556 3738
rect 94504 3674 94556 3680
rect 93490 3088 93546 3097
rect 93490 3023 93546 3032
rect 88524 2984 88576 2990
rect 88524 2926 88576 2932
rect 83004 2848 83056 2854
rect 83004 2790 83056 2796
rect 81452 2746 81756 2774
rect 81452 2650 81480 2746
rect 81440 2644 81492 2650
rect 81440 2586 81492 2592
rect 74540 2382 74592 2388
rect 75472 2378 75592 2394
rect 81348 2440 81400 2446
rect 81348 2382 81400 2388
rect 83016 2378 83044 2790
rect 95620 2417 95648 11222
rect 95700 9920 95752 9926
rect 95700 9862 95752 9868
rect 96160 9920 96212 9926
rect 96160 9862 96212 9868
rect 95712 9654 95740 9862
rect 95700 9648 95752 9654
rect 95700 9590 95752 9596
rect 96172 8974 96200 9862
rect 96160 8968 96212 8974
rect 96160 8910 96212 8916
rect 96540 7410 96568 12038
rect 96632 11762 96660 13194
rect 96712 13184 96764 13190
rect 96712 13126 96764 13132
rect 96804 13184 96856 13190
rect 96804 13126 96856 13132
rect 96620 11756 96672 11762
rect 96620 11698 96672 11704
rect 96724 11694 96752 13126
rect 96816 12986 96844 13126
rect 96804 12980 96856 12986
rect 96804 12922 96856 12928
rect 96908 12714 96936 13194
rect 97644 12986 97672 15286
rect 97906 15200 97962 16000
rect 98458 15200 98514 16000
rect 99010 15200 99066 16000
rect 99562 15200 99618 16000
rect 100114 15200 100170 16000
rect 100666 15200 100722 16000
rect 101218 15200 101274 16000
rect 101770 15200 101826 16000
rect 102322 15314 102378 16000
rect 102322 15286 102640 15314
rect 102322 15200 102378 15286
rect 97920 13546 97948 15200
rect 97920 13530 98040 13546
rect 97920 13524 98052 13530
rect 97920 13518 98000 13524
rect 98000 13466 98052 13472
rect 98472 13462 98500 15200
rect 98736 13796 98788 13802
rect 98736 13738 98788 13744
rect 98460 13456 98512 13462
rect 98460 13398 98512 13404
rect 97724 13320 97776 13326
rect 97724 13262 97776 13268
rect 97736 13161 97764 13262
rect 97722 13152 97778 13161
rect 97722 13087 97778 13096
rect 97632 12980 97684 12986
rect 97632 12922 97684 12928
rect 98552 12980 98604 12986
rect 98552 12922 98604 12928
rect 98460 12912 98512 12918
rect 98460 12854 98512 12860
rect 98000 12844 98052 12850
rect 98000 12786 98052 12792
rect 96896 12708 96948 12714
rect 96896 12650 96948 12656
rect 96988 12708 97040 12714
rect 96988 12650 97040 12656
rect 96802 12336 96858 12345
rect 96802 12271 96858 12280
rect 96816 11801 96844 12271
rect 97000 12238 97028 12650
rect 98012 12646 98040 12786
rect 98000 12640 98052 12646
rect 98000 12582 98052 12588
rect 98184 12368 98236 12374
rect 98184 12310 98236 12316
rect 96988 12232 97040 12238
rect 96988 12174 97040 12180
rect 98196 12170 98224 12310
rect 98184 12164 98236 12170
rect 98184 12106 98236 12112
rect 98472 11898 98500 12854
rect 98184 11892 98236 11898
rect 98184 11834 98236 11840
rect 98460 11892 98512 11898
rect 98460 11834 98512 11840
rect 96802 11792 96858 11801
rect 96802 11727 96858 11736
rect 96712 11688 96764 11694
rect 96712 11630 96764 11636
rect 96816 11286 96844 11727
rect 96804 11280 96856 11286
rect 96804 11222 96856 11228
rect 98196 11218 98224 11834
rect 98472 11801 98500 11834
rect 98458 11792 98514 11801
rect 98458 11727 98514 11736
rect 98184 11212 98236 11218
rect 98184 11154 98236 11160
rect 98276 11076 98328 11082
rect 98276 11018 98328 11024
rect 98288 10470 98316 11018
rect 97080 10464 97132 10470
rect 97080 10406 97132 10412
rect 98276 10464 98328 10470
rect 98276 10406 98328 10412
rect 98368 10464 98420 10470
rect 98368 10406 98420 10412
rect 97092 10062 97120 10406
rect 98288 10062 98316 10406
rect 98380 10130 98408 10406
rect 98368 10124 98420 10130
rect 98368 10066 98420 10072
rect 97080 10056 97132 10062
rect 97080 9998 97132 10004
rect 98276 10056 98328 10062
rect 98276 9998 98328 10004
rect 97092 7698 97120 9998
rect 98092 9920 98144 9926
rect 98092 9862 98144 9868
rect 98104 9722 98132 9862
rect 98092 9716 98144 9722
rect 98092 9658 98144 9664
rect 97356 9444 97408 9450
rect 97356 9386 97408 9392
rect 97000 7670 97120 7698
rect 96896 7540 96948 7546
rect 96896 7482 96948 7488
rect 96528 7404 96580 7410
rect 96528 7346 96580 7352
rect 96804 7404 96856 7410
rect 96804 7346 96856 7352
rect 96816 6866 96844 7346
rect 96908 7342 96936 7482
rect 96896 7336 96948 7342
rect 96896 7278 96948 7284
rect 97000 7274 97028 7670
rect 97368 7546 97396 9386
rect 98092 9104 98144 9110
rect 97644 9064 98092 9092
rect 97644 8838 97672 9064
rect 98092 9046 98144 9052
rect 98000 8968 98052 8974
rect 97736 8916 98000 8922
rect 97736 8910 98052 8916
rect 97736 8906 98040 8910
rect 97724 8900 98040 8906
rect 97776 8894 98040 8900
rect 97724 8842 97776 8848
rect 97632 8832 97684 8838
rect 97632 8774 97684 8780
rect 97540 8288 97592 8294
rect 97540 8230 97592 8236
rect 97356 7540 97408 7546
rect 97356 7482 97408 7488
rect 97448 7540 97500 7546
rect 97448 7482 97500 7488
rect 97368 7410 97396 7482
rect 97356 7404 97408 7410
rect 97356 7346 97408 7352
rect 96988 7268 97040 7274
rect 96988 7210 97040 7216
rect 96804 6860 96856 6866
rect 96804 6802 96856 6808
rect 96896 6860 96948 6866
rect 96896 6802 96948 6808
rect 96908 6662 96936 6802
rect 96896 6656 96948 6662
rect 96896 6598 96948 6604
rect 96620 6248 96672 6254
rect 96620 6190 96672 6196
rect 96632 6118 96660 6190
rect 96620 6112 96672 6118
rect 96620 6054 96672 6060
rect 96632 5914 96660 6054
rect 96620 5908 96672 5914
rect 96620 5850 96672 5856
rect 96632 4690 96660 5850
rect 96712 5228 96764 5234
rect 96712 5170 96764 5176
rect 96620 4684 96672 4690
rect 96620 4626 96672 4632
rect 96252 3528 96304 3534
rect 96252 3470 96304 3476
rect 96264 3194 96292 3470
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96724 2961 96752 5170
rect 97000 3058 97028 7210
rect 97460 7206 97488 7482
rect 97552 7206 97580 8230
rect 98012 7868 98040 8894
rect 98184 8832 98236 8838
rect 98184 8774 98236 8780
rect 98196 8498 98224 8774
rect 98184 8492 98236 8498
rect 98184 8434 98236 8440
rect 98092 7880 98144 7886
rect 98012 7840 98092 7868
rect 97816 7744 97868 7750
rect 98012 7698 98040 7840
rect 98092 7822 98144 7828
rect 97868 7692 98040 7698
rect 97816 7686 98040 7692
rect 97828 7670 98040 7686
rect 97448 7200 97500 7206
rect 97448 7142 97500 7148
rect 97540 7200 97592 7206
rect 97540 7142 97592 7148
rect 97356 6656 97408 6662
rect 97356 6598 97408 6604
rect 97368 6322 97396 6598
rect 97356 6316 97408 6322
rect 97356 6258 97408 6264
rect 98196 4826 98224 8434
rect 98276 8288 98328 8294
rect 98276 8230 98328 8236
rect 98288 8022 98316 8230
rect 98276 8016 98328 8022
rect 98276 7958 98328 7964
rect 98564 7834 98592 12922
rect 98748 12442 98776 13738
rect 99024 13190 99052 15200
rect 99576 13818 99604 15200
rect 99484 13790 99604 13818
rect 99484 13410 99512 13790
rect 99562 13628 99870 13637
rect 99562 13626 99568 13628
rect 99624 13626 99648 13628
rect 99704 13626 99728 13628
rect 99784 13626 99808 13628
rect 99864 13626 99870 13628
rect 99624 13574 99626 13626
rect 99806 13574 99808 13626
rect 99562 13572 99568 13574
rect 99624 13572 99648 13574
rect 99704 13572 99728 13574
rect 99784 13572 99808 13574
rect 99864 13572 99870 13574
rect 99562 13563 99870 13572
rect 99484 13382 99604 13410
rect 99472 13320 99524 13326
rect 99472 13262 99524 13268
rect 99012 13184 99064 13190
rect 99012 13126 99064 13132
rect 99380 12776 99432 12782
rect 99380 12718 99432 12724
rect 99288 12640 99340 12646
rect 99288 12582 99340 12588
rect 98736 12436 98788 12442
rect 98736 12378 98788 12384
rect 99300 12238 99328 12582
rect 99288 12232 99340 12238
rect 99288 12174 99340 12180
rect 99012 11756 99064 11762
rect 99012 11698 99064 11704
rect 98736 11144 98788 11150
rect 98736 11086 98788 11092
rect 98644 11008 98696 11014
rect 98644 10950 98696 10956
rect 98472 7818 98592 7834
rect 98460 7812 98592 7818
rect 98512 7806 98592 7812
rect 98460 7754 98512 7760
rect 98184 4820 98236 4826
rect 98184 4762 98236 4768
rect 98552 4548 98604 4554
rect 98552 4490 98604 4496
rect 98564 4282 98592 4490
rect 98552 4276 98604 4282
rect 98552 4218 98604 4224
rect 96988 3052 97040 3058
rect 96988 2994 97040 3000
rect 96710 2952 96766 2961
rect 96710 2887 96766 2896
rect 98656 2854 98684 10950
rect 98748 9654 98776 11086
rect 98828 11008 98880 11014
rect 98828 10950 98880 10956
rect 98840 10742 98868 10950
rect 98828 10736 98880 10742
rect 98828 10678 98880 10684
rect 98828 10600 98880 10606
rect 98828 10542 98880 10548
rect 98840 10198 98868 10542
rect 98828 10192 98880 10198
rect 98828 10134 98880 10140
rect 98840 9738 98868 10134
rect 98840 9722 98960 9738
rect 98840 9716 98972 9722
rect 98840 9710 98920 9716
rect 98920 9658 98972 9664
rect 98736 9648 98788 9654
rect 98736 9590 98788 9596
rect 99024 3670 99052 11698
rect 99392 11694 99420 12718
rect 99380 11688 99432 11694
rect 99378 11656 99380 11665
rect 99432 11656 99434 11665
rect 99378 11591 99434 11600
rect 99484 11014 99512 13262
rect 99576 12714 99604 13382
rect 100024 13320 100076 13326
rect 99930 13288 99986 13297
rect 100024 13262 100076 13268
rect 99930 13223 99986 13232
rect 99564 12708 99616 12714
rect 99564 12650 99616 12656
rect 99562 12540 99870 12549
rect 99562 12538 99568 12540
rect 99624 12538 99648 12540
rect 99704 12538 99728 12540
rect 99784 12538 99808 12540
rect 99864 12538 99870 12540
rect 99624 12486 99626 12538
rect 99806 12486 99808 12538
rect 99562 12484 99568 12486
rect 99624 12484 99648 12486
rect 99704 12484 99728 12486
rect 99784 12484 99808 12486
rect 99864 12484 99870 12486
rect 99562 12475 99870 12484
rect 99944 12442 99972 13223
rect 100036 12986 100064 13262
rect 100128 12986 100156 15200
rect 100298 13152 100354 13161
rect 100298 13087 100354 13096
rect 100024 12980 100076 12986
rect 100024 12922 100076 12928
rect 100116 12980 100168 12986
rect 100116 12922 100168 12928
rect 100116 12844 100168 12850
rect 100116 12786 100168 12792
rect 99932 12436 99984 12442
rect 99984 12406 100064 12434
rect 99932 12378 99984 12384
rect 99932 11892 99984 11898
rect 99932 11834 99984 11840
rect 99562 11452 99870 11461
rect 99562 11450 99568 11452
rect 99624 11450 99648 11452
rect 99704 11450 99728 11452
rect 99784 11450 99808 11452
rect 99864 11450 99870 11452
rect 99624 11398 99626 11450
rect 99806 11398 99808 11450
rect 99562 11396 99568 11398
rect 99624 11396 99648 11398
rect 99704 11396 99728 11398
rect 99784 11396 99808 11398
rect 99864 11396 99870 11398
rect 99562 11387 99870 11396
rect 99472 11008 99524 11014
rect 99472 10950 99524 10956
rect 99562 10364 99870 10373
rect 99562 10362 99568 10364
rect 99624 10362 99648 10364
rect 99704 10362 99728 10364
rect 99784 10362 99808 10364
rect 99864 10362 99870 10364
rect 99624 10310 99626 10362
rect 99806 10310 99808 10362
rect 99562 10308 99568 10310
rect 99624 10308 99648 10310
rect 99704 10308 99728 10310
rect 99784 10308 99808 10310
rect 99864 10308 99870 10310
rect 99562 10299 99870 10308
rect 99472 9988 99524 9994
rect 99472 9930 99524 9936
rect 99380 9580 99432 9586
rect 99380 9522 99432 9528
rect 99392 9110 99420 9522
rect 99380 9104 99432 9110
rect 99380 9046 99432 9052
rect 99484 8974 99512 9930
rect 99562 9276 99870 9285
rect 99562 9274 99568 9276
rect 99624 9274 99648 9276
rect 99704 9274 99728 9276
rect 99784 9274 99808 9276
rect 99864 9274 99870 9276
rect 99624 9222 99626 9274
rect 99806 9222 99808 9274
rect 99562 9220 99568 9222
rect 99624 9220 99648 9222
rect 99704 9220 99728 9222
rect 99784 9220 99808 9222
rect 99864 9220 99870 9222
rect 99562 9211 99870 9220
rect 99748 9104 99800 9110
rect 99944 9058 99972 11834
rect 99800 9052 99972 9058
rect 99748 9046 99972 9052
rect 99760 9030 99972 9046
rect 99472 8968 99524 8974
rect 99472 8910 99524 8916
rect 99380 8832 99432 8838
rect 99380 8774 99432 8780
rect 99196 7812 99248 7818
rect 99196 7754 99248 7760
rect 99208 7342 99236 7754
rect 99196 7336 99248 7342
rect 99196 7278 99248 7284
rect 99392 6730 99420 8774
rect 99562 8188 99870 8197
rect 99562 8186 99568 8188
rect 99624 8186 99648 8188
rect 99704 8186 99728 8188
rect 99784 8186 99808 8188
rect 99864 8186 99870 8188
rect 99624 8134 99626 8186
rect 99806 8134 99808 8186
rect 99562 8132 99568 8134
rect 99624 8132 99648 8134
rect 99704 8132 99728 8134
rect 99784 8132 99808 8134
rect 99864 8132 99870 8134
rect 99562 8123 99870 8132
rect 99562 7100 99870 7109
rect 99562 7098 99568 7100
rect 99624 7098 99648 7100
rect 99704 7098 99728 7100
rect 99784 7098 99808 7100
rect 99864 7098 99870 7100
rect 99624 7046 99626 7098
rect 99806 7046 99808 7098
rect 99562 7044 99568 7046
rect 99624 7044 99648 7046
rect 99704 7044 99728 7046
rect 99784 7044 99808 7046
rect 99864 7044 99870 7046
rect 99562 7035 99870 7044
rect 99380 6724 99432 6730
rect 99380 6666 99432 6672
rect 99562 6012 99870 6021
rect 99562 6010 99568 6012
rect 99624 6010 99648 6012
rect 99704 6010 99728 6012
rect 99784 6010 99808 6012
rect 99864 6010 99870 6012
rect 99624 5958 99626 6010
rect 99806 5958 99808 6010
rect 99562 5956 99568 5958
rect 99624 5956 99648 5958
rect 99704 5956 99728 5958
rect 99784 5956 99808 5958
rect 99864 5956 99870 5958
rect 99562 5947 99870 5956
rect 99932 5840 99984 5846
rect 99932 5782 99984 5788
rect 99944 5574 99972 5782
rect 99932 5568 99984 5574
rect 99932 5510 99984 5516
rect 99944 5273 99972 5510
rect 99930 5264 99986 5273
rect 99930 5199 99986 5208
rect 100036 5137 100064 12406
rect 100128 8022 100156 12786
rect 100208 12776 100260 12782
rect 100208 12718 100260 12724
rect 100220 11898 100248 12718
rect 100312 12238 100340 13087
rect 100392 12912 100444 12918
rect 100392 12854 100444 12860
rect 100300 12232 100352 12238
rect 100300 12174 100352 12180
rect 100208 11892 100260 11898
rect 100208 11834 100260 11840
rect 100312 8242 100340 12174
rect 100404 12102 100432 12854
rect 100680 12714 100708 15200
rect 100760 14000 100812 14006
rect 100760 13942 100812 13948
rect 100668 12708 100720 12714
rect 100668 12650 100720 12656
rect 100392 12096 100444 12102
rect 100392 12038 100444 12044
rect 100404 8430 100432 12038
rect 100668 11552 100720 11558
rect 100668 11494 100720 11500
rect 100680 11121 100708 11494
rect 100666 11112 100722 11121
rect 100666 11047 100722 11056
rect 100680 8945 100708 11047
rect 100772 10266 100800 13942
rect 101232 13462 101260 15200
rect 101220 13456 101272 13462
rect 101220 13398 101272 13404
rect 101784 12986 101812 15200
rect 102324 13796 102376 13802
rect 102324 13738 102376 13744
rect 102336 13326 102364 13738
rect 101864 13320 101916 13326
rect 101864 13262 101916 13268
rect 102324 13320 102376 13326
rect 102324 13262 102376 13268
rect 102508 13320 102560 13326
rect 102508 13262 102560 13268
rect 101772 12980 101824 12986
rect 101772 12922 101824 12928
rect 101312 12844 101364 12850
rect 101312 12786 101364 12792
rect 101036 12164 101088 12170
rect 101036 12106 101088 12112
rect 101048 11626 101076 12106
rect 101324 12102 101352 12786
rect 101876 12434 101904 13262
rect 102048 12436 102100 12442
rect 101876 12406 101996 12434
rect 101404 12368 101456 12374
rect 101404 12310 101456 12316
rect 101312 12096 101364 12102
rect 101312 12038 101364 12044
rect 101036 11620 101088 11626
rect 101036 11562 101088 11568
rect 101416 11150 101444 12310
rect 101588 12300 101640 12306
rect 101588 12242 101640 12248
rect 101496 12096 101548 12102
rect 101496 12038 101548 12044
rect 101404 11144 101456 11150
rect 101404 11086 101456 11092
rect 101128 11008 101180 11014
rect 101128 10950 101180 10956
rect 100852 10804 100904 10810
rect 100852 10746 100904 10752
rect 100864 10470 100892 10746
rect 101140 10538 101168 10950
rect 101128 10532 101180 10538
rect 101128 10474 101180 10480
rect 100852 10464 100904 10470
rect 100852 10406 100904 10412
rect 100760 10260 100812 10266
rect 100760 10202 100812 10208
rect 100772 9994 100800 10202
rect 101128 10192 101180 10198
rect 101128 10134 101180 10140
rect 101140 9994 101168 10134
rect 100760 9988 100812 9994
rect 100760 9930 100812 9936
rect 101128 9988 101180 9994
rect 101128 9930 101180 9936
rect 101220 9444 101272 9450
rect 101220 9386 101272 9392
rect 101232 9178 101260 9386
rect 101036 9172 101088 9178
rect 101036 9114 101088 9120
rect 101220 9172 101272 9178
rect 101220 9114 101272 9120
rect 100666 8936 100722 8945
rect 100666 8871 100722 8880
rect 101048 8498 101076 9114
rect 101036 8492 101088 8498
rect 101036 8434 101088 8440
rect 100392 8424 100444 8430
rect 100392 8366 100444 8372
rect 100312 8214 100432 8242
rect 100116 8016 100168 8022
rect 100116 7958 100168 7964
rect 100300 7744 100352 7750
rect 100404 7721 100432 8214
rect 100300 7686 100352 7692
rect 100390 7712 100446 7721
rect 100312 6225 100340 7686
rect 100390 7647 100446 7656
rect 100758 6896 100814 6905
rect 100758 6831 100814 6840
rect 100772 6254 100800 6831
rect 100760 6248 100812 6254
rect 100298 6216 100354 6225
rect 100760 6190 100812 6196
rect 100852 6248 100904 6254
rect 100852 6190 100904 6196
rect 100298 6151 100354 6160
rect 100022 5128 100078 5137
rect 100022 5063 100078 5072
rect 99562 4924 99870 4933
rect 99562 4922 99568 4924
rect 99624 4922 99648 4924
rect 99704 4922 99728 4924
rect 99784 4922 99808 4924
rect 99864 4922 99870 4924
rect 99624 4870 99626 4922
rect 99806 4870 99808 4922
rect 99562 4868 99568 4870
rect 99624 4868 99648 4870
rect 99704 4868 99728 4870
rect 99784 4868 99808 4870
rect 99864 4868 99870 4870
rect 99562 4859 99870 4868
rect 99562 3836 99870 3845
rect 99562 3834 99568 3836
rect 99624 3834 99648 3836
rect 99704 3834 99728 3836
rect 99784 3834 99808 3836
rect 99864 3834 99870 3836
rect 99624 3782 99626 3834
rect 99806 3782 99808 3834
rect 99562 3780 99568 3782
rect 99624 3780 99648 3782
rect 99704 3780 99728 3782
rect 99784 3780 99808 3782
rect 99864 3780 99870 3782
rect 99562 3771 99870 3780
rect 99012 3664 99064 3670
rect 99012 3606 99064 3612
rect 100864 2922 100892 6190
rect 100944 6112 100996 6118
rect 100944 6054 100996 6060
rect 100956 5642 100984 6054
rect 101312 5908 101364 5914
rect 101312 5850 101364 5856
rect 101324 5710 101352 5850
rect 101508 5778 101536 12038
rect 101600 11830 101628 12242
rect 101968 12102 101996 12406
rect 102048 12378 102100 12384
rect 101956 12096 102008 12102
rect 101956 12038 102008 12044
rect 101588 11824 101640 11830
rect 101588 11766 101640 11772
rect 101968 11762 101996 12038
rect 101772 11756 101824 11762
rect 101772 11698 101824 11704
rect 101956 11756 102008 11762
rect 101956 11698 102008 11704
rect 101680 11280 101732 11286
rect 101680 11222 101732 11228
rect 101692 8362 101720 11222
rect 101680 8356 101732 8362
rect 101680 8298 101732 8304
rect 101588 6860 101640 6866
rect 101588 6802 101640 6808
rect 101600 6730 101628 6802
rect 101588 6724 101640 6730
rect 101588 6666 101640 6672
rect 101600 6322 101628 6666
rect 101588 6316 101640 6322
rect 101588 6258 101640 6264
rect 101496 5772 101548 5778
rect 101496 5714 101548 5720
rect 101312 5704 101364 5710
rect 101312 5646 101364 5652
rect 100944 5636 100996 5642
rect 100944 5578 100996 5584
rect 101324 5166 101352 5646
rect 101312 5160 101364 5166
rect 101312 5102 101364 5108
rect 101692 4622 101720 8298
rect 101680 4616 101732 4622
rect 101680 4558 101732 4564
rect 101784 4486 101812 11698
rect 101862 10296 101918 10305
rect 101862 10231 101918 10240
rect 101876 10198 101904 10231
rect 101864 10192 101916 10198
rect 101864 10134 101916 10140
rect 101876 8294 101904 10134
rect 101864 8288 101916 8294
rect 101864 8230 101916 8236
rect 101864 6316 101916 6322
rect 101864 6258 101916 6264
rect 101876 6089 101904 6258
rect 101862 6080 101918 6089
rect 101862 6015 101918 6024
rect 101956 5568 102008 5574
rect 101956 5510 102008 5516
rect 101772 4480 101824 4486
rect 101772 4422 101824 4428
rect 100852 2916 100904 2922
rect 100852 2858 100904 2864
rect 98644 2848 98696 2854
rect 98644 2790 98696 2796
rect 99562 2748 99870 2757
rect 99562 2746 99568 2748
rect 99624 2746 99648 2748
rect 99704 2746 99728 2748
rect 99784 2746 99808 2748
rect 99864 2746 99870 2748
rect 99624 2694 99626 2746
rect 99806 2694 99808 2746
rect 99562 2692 99568 2694
rect 99624 2692 99648 2694
rect 99704 2692 99728 2694
rect 99784 2692 99808 2694
rect 99864 2692 99870 2694
rect 99562 2683 99870 2692
rect 95606 2408 95662 2417
rect 45376 2372 45428 2378
rect 45376 2314 45428 2320
rect 75460 2372 75592 2378
rect 75512 2366 75592 2372
rect 83004 2372 83056 2378
rect 75460 2314 75512 2320
rect 95606 2343 95662 2352
rect 83004 2314 83056 2320
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 32404 2304 32456 2310
rect 32404 2246 32456 2252
rect 31772 2038 31800 2246
rect 32416 2106 32444 2246
rect 40394 2204 40702 2213
rect 40394 2202 40400 2204
rect 40456 2202 40480 2204
rect 40536 2202 40560 2204
rect 40616 2202 40640 2204
rect 40696 2202 40702 2204
rect 40456 2150 40458 2202
rect 40638 2150 40640 2202
rect 40394 2148 40400 2150
rect 40456 2148 40480 2150
rect 40536 2148 40560 2150
rect 40616 2148 40640 2150
rect 40696 2148 40702 2150
rect 40394 2139 40702 2148
rect 79839 2204 80147 2213
rect 79839 2202 79845 2204
rect 79901 2202 79925 2204
rect 79981 2202 80005 2204
rect 80061 2202 80085 2204
rect 80141 2202 80147 2204
rect 79901 2150 79903 2202
rect 80083 2150 80085 2202
rect 79839 2148 79845 2150
rect 79901 2148 79925 2150
rect 79981 2148 80005 2150
rect 80061 2148 80085 2150
rect 80141 2148 80147 2150
rect 79839 2139 80147 2148
rect 32404 2100 32456 2106
rect 32404 2042 32456 2048
rect 15568 2032 15620 2038
rect 1674 2000 1730 2009
rect 15568 1974 15620 1980
rect 31760 2032 31812 2038
rect 31760 1974 31812 1980
rect 1674 1935 1730 1944
rect 101968 1086 101996 5510
rect 102060 3738 102088 12378
rect 102324 12096 102376 12102
rect 102324 12038 102376 12044
rect 102232 11212 102284 11218
rect 102232 11154 102284 11160
rect 102244 10810 102272 11154
rect 102140 10804 102192 10810
rect 102140 10746 102192 10752
rect 102232 10804 102284 10810
rect 102232 10746 102284 10752
rect 102152 6458 102180 10746
rect 102244 10266 102272 10746
rect 102336 10742 102364 12038
rect 102324 10736 102376 10742
rect 102324 10678 102376 10684
rect 102232 10260 102284 10266
rect 102232 10202 102284 10208
rect 102520 6905 102548 13262
rect 102612 12986 102640 15286
rect 102874 15200 102930 16000
rect 103426 15200 103482 16000
rect 103978 15200 104034 16000
rect 104530 15314 104586 16000
rect 104530 15286 104848 15314
rect 104530 15200 104586 15286
rect 102888 13530 102916 15200
rect 103440 13546 103468 15200
rect 102876 13524 102928 13530
rect 103440 13518 103560 13546
rect 102876 13466 102928 13472
rect 103532 13462 103560 13518
rect 103520 13456 103572 13462
rect 103520 13398 103572 13404
rect 103060 13320 103112 13326
rect 103060 13262 103112 13268
rect 103072 13190 103100 13262
rect 102968 13184 103020 13190
rect 102968 13126 103020 13132
rect 103060 13184 103112 13190
rect 103060 13126 103112 13132
rect 102600 12980 102652 12986
rect 102600 12922 102652 12928
rect 102980 12238 103008 13126
rect 103992 12986 104020 15200
rect 104256 13932 104308 13938
rect 104256 13874 104308 13880
rect 104164 13728 104216 13734
rect 104164 13670 104216 13676
rect 104176 13394 104204 13670
rect 104164 13388 104216 13394
rect 104164 13330 104216 13336
rect 104072 13320 104124 13326
rect 104072 13262 104124 13268
rect 103980 12980 104032 12986
rect 103980 12922 104032 12928
rect 104084 12918 104112 13262
rect 103888 12912 103940 12918
rect 103888 12854 103940 12860
rect 104072 12912 104124 12918
rect 104072 12854 104124 12860
rect 103900 12782 103928 12854
rect 103612 12776 103664 12782
rect 103888 12776 103940 12782
rect 103612 12718 103664 12724
rect 103886 12744 103888 12753
rect 103940 12744 103942 12753
rect 102968 12232 103020 12238
rect 102968 12174 103020 12180
rect 103060 12232 103112 12238
rect 103060 12174 103112 12180
rect 103072 11898 103100 12174
rect 103624 12102 103652 12718
rect 103886 12679 103942 12688
rect 103796 12640 103848 12646
rect 103796 12582 103848 12588
rect 103612 12096 103664 12102
rect 103612 12038 103664 12044
rect 103060 11892 103112 11898
rect 103060 11834 103112 11840
rect 103520 11892 103572 11898
rect 103520 11834 103572 11840
rect 103428 11552 103480 11558
rect 103428 11494 103480 11500
rect 103440 11150 103468 11494
rect 103428 11144 103480 11150
rect 103428 11086 103480 11092
rect 103336 11008 103388 11014
rect 103336 10950 103388 10956
rect 103348 10674 103376 10950
rect 103440 10742 103468 11086
rect 103532 11082 103560 11834
rect 103520 11076 103572 11082
rect 103520 11018 103572 11024
rect 103428 10736 103480 10742
rect 103428 10678 103480 10684
rect 103336 10668 103388 10674
rect 103336 10610 103388 10616
rect 102876 10260 102928 10266
rect 102876 10202 102928 10208
rect 102888 9994 102916 10202
rect 103440 10130 103468 10678
rect 103428 10124 103480 10130
rect 103428 10066 103480 10072
rect 102876 9988 102928 9994
rect 102876 9930 102928 9936
rect 103428 9988 103480 9994
rect 103428 9930 103480 9936
rect 103440 9382 103468 9930
rect 103244 9376 103296 9382
rect 103244 9318 103296 9324
rect 103428 9376 103480 9382
rect 103428 9318 103480 9324
rect 103256 9178 103284 9318
rect 103244 9172 103296 9178
rect 103244 9114 103296 9120
rect 102506 6896 102562 6905
rect 102506 6831 102562 6840
rect 102140 6452 102192 6458
rect 102140 6394 102192 6400
rect 103440 5914 103468 9318
rect 103624 6866 103652 12038
rect 103808 11218 103836 12582
rect 104268 11898 104296 13874
rect 104348 13796 104400 13802
rect 104348 13738 104400 13744
rect 104360 12434 104388 13738
rect 104820 13530 104848 15286
rect 105082 15200 105138 16000
rect 105634 15200 105690 16000
rect 106186 15200 106242 16000
rect 106738 15200 106794 16000
rect 107290 15200 107346 16000
rect 107842 15200 107898 16000
rect 108394 15200 108450 16000
rect 108946 15200 109002 16000
rect 109498 15314 109554 16000
rect 110050 15314 110106 16000
rect 109498 15286 109816 15314
rect 109498 15200 109554 15286
rect 104808 13524 104860 13530
rect 104808 13466 104860 13472
rect 104808 12980 104860 12986
rect 104808 12922 104860 12928
rect 104820 12646 104848 12922
rect 104900 12844 104952 12850
rect 104900 12786 104952 12792
rect 104808 12640 104860 12646
rect 104808 12582 104860 12588
rect 104624 12436 104676 12442
rect 104360 12406 104480 12434
rect 104348 12232 104400 12238
rect 104348 12174 104400 12180
rect 104360 12073 104388 12174
rect 104346 12064 104402 12073
rect 104346 11999 104402 12008
rect 104256 11892 104308 11898
rect 104256 11834 104308 11840
rect 103796 11212 103848 11218
rect 103796 11154 103848 11160
rect 103808 10810 103836 11154
rect 103796 10804 103848 10810
rect 103796 10746 103848 10752
rect 104348 10736 104400 10742
rect 104348 10678 104400 10684
rect 104072 10600 104124 10606
rect 104072 10542 104124 10548
rect 104084 10130 104112 10542
rect 104162 10432 104218 10441
rect 104162 10367 104218 10376
rect 104072 10124 104124 10130
rect 104072 10066 104124 10072
rect 104176 9897 104204 10367
rect 104360 10266 104388 10678
rect 104348 10260 104400 10266
rect 104348 10202 104400 10208
rect 104162 9888 104218 9897
rect 104162 9823 104218 9832
rect 104452 9586 104480 12406
rect 104624 12378 104676 12384
rect 104636 12238 104664 12378
rect 104624 12232 104676 12238
rect 104624 12174 104676 12180
rect 104716 11892 104768 11898
rect 104716 11834 104768 11840
rect 104532 10600 104584 10606
rect 104532 10542 104584 10548
rect 104544 10266 104572 10542
rect 104532 10260 104584 10266
rect 104532 10202 104584 10208
rect 104544 9926 104572 10202
rect 104728 10169 104756 11834
rect 104714 10160 104770 10169
rect 104714 10095 104770 10104
rect 104532 9920 104584 9926
rect 104532 9862 104584 9868
rect 104256 9580 104308 9586
rect 104256 9522 104308 9528
rect 104440 9580 104492 9586
rect 104440 9522 104492 9528
rect 104624 9580 104676 9586
rect 104624 9522 104676 9528
rect 104268 8362 104296 9522
rect 104452 9110 104480 9522
rect 104440 9104 104492 9110
rect 104440 9046 104492 9052
rect 104636 9042 104664 9522
rect 104624 9036 104676 9042
rect 104624 8978 104676 8984
rect 104636 8906 104664 8978
rect 104624 8900 104676 8906
rect 104624 8842 104676 8848
rect 104256 8356 104308 8362
rect 104256 8298 104308 8304
rect 104728 7993 104756 10095
rect 104808 9920 104860 9926
rect 104912 9874 104940 12786
rect 105096 12442 105124 15200
rect 105648 12442 105676 15200
rect 105728 12776 105780 12782
rect 105728 12718 105780 12724
rect 105084 12436 105136 12442
rect 105084 12378 105136 12384
rect 105636 12436 105688 12442
rect 105636 12378 105688 12384
rect 105636 12096 105688 12102
rect 105636 12038 105688 12044
rect 105176 11008 105228 11014
rect 105176 10950 105228 10956
rect 105188 10305 105216 10950
rect 104990 10296 105046 10305
rect 104990 10231 105046 10240
rect 105174 10296 105230 10305
rect 105174 10231 105230 10240
rect 105004 9994 105032 10231
rect 104992 9988 105044 9994
rect 104992 9930 105044 9936
rect 104860 9868 104940 9874
rect 104808 9862 104940 9868
rect 104820 9846 104940 9862
rect 104714 7984 104770 7993
rect 104714 7919 104770 7928
rect 104912 7818 104940 9846
rect 105648 9586 105676 12038
rect 105740 11082 105768 12718
rect 106200 12628 106228 15200
rect 106648 13796 106700 13802
rect 106648 13738 106700 13744
rect 106660 13530 106688 13738
rect 106648 13524 106700 13530
rect 106648 13466 106700 13472
rect 106372 13184 106424 13190
rect 106372 13126 106424 13132
rect 106280 12640 106332 12646
rect 106200 12600 106280 12628
rect 106280 12582 106332 12588
rect 106384 12434 106412 13126
rect 106752 12442 106780 15200
rect 106832 13796 106884 13802
rect 106832 13738 106884 13744
rect 106740 12436 106792 12442
rect 106384 12406 106504 12434
rect 106372 12300 106424 12306
rect 106372 12242 106424 12248
rect 106188 12232 106240 12238
rect 106188 12174 106240 12180
rect 105820 12096 105872 12102
rect 105818 12064 105820 12073
rect 105872 12064 105874 12073
rect 105818 11999 105874 12008
rect 106200 11898 106228 12174
rect 106188 11892 106240 11898
rect 106188 11834 106240 11840
rect 106384 11626 106412 12242
rect 106372 11620 106424 11626
rect 106372 11562 106424 11568
rect 106476 11218 106504 12406
rect 106740 12378 106792 12384
rect 106464 11212 106516 11218
rect 106464 11154 106516 11160
rect 106648 11212 106700 11218
rect 106648 11154 106700 11160
rect 105820 11144 105872 11150
rect 105820 11086 105872 11092
rect 105728 11076 105780 11082
rect 105728 11018 105780 11024
rect 105636 9580 105688 9586
rect 105636 9522 105688 9528
rect 105360 9376 105412 9382
rect 105360 9318 105412 9324
rect 105452 9376 105504 9382
rect 105452 9318 105504 9324
rect 105372 7886 105400 9318
rect 105360 7880 105412 7886
rect 105360 7822 105412 7828
rect 104900 7812 104952 7818
rect 104900 7754 104952 7760
rect 103612 6860 103664 6866
rect 103612 6802 103664 6808
rect 105464 6798 105492 9318
rect 105740 6798 105768 11018
rect 105832 9586 105860 11086
rect 106372 11076 106424 11082
rect 106372 11018 106424 11024
rect 105912 11008 105964 11014
rect 105912 10950 105964 10956
rect 105924 10198 105952 10950
rect 105912 10192 105964 10198
rect 105912 10134 105964 10140
rect 105820 9580 105872 9586
rect 105820 9522 105872 9528
rect 105452 6792 105504 6798
rect 105452 6734 105504 6740
rect 105728 6792 105780 6798
rect 105728 6734 105780 6740
rect 106384 6662 106412 11018
rect 106462 6760 106518 6769
rect 106462 6695 106518 6704
rect 106372 6656 106424 6662
rect 106372 6598 106424 6604
rect 106476 6458 106504 6695
rect 106464 6452 106516 6458
rect 106464 6394 106516 6400
rect 105176 6316 105228 6322
rect 105176 6258 105228 6264
rect 105084 6180 105136 6186
rect 105084 6122 105136 6128
rect 103428 5908 103480 5914
rect 103428 5850 103480 5856
rect 105096 5846 105124 6122
rect 105084 5840 105136 5846
rect 105084 5782 105136 5788
rect 105188 5234 105216 6258
rect 106096 6248 106148 6254
rect 106096 6190 106148 6196
rect 106108 5778 106136 6190
rect 106660 5846 106688 11154
rect 106740 11144 106792 11150
rect 106740 11086 106792 11092
rect 106752 7818 106780 11086
rect 106844 10266 106872 13738
rect 107016 13320 107068 13326
rect 107016 13262 107068 13268
rect 107028 12986 107056 13262
rect 107304 12986 107332 15200
rect 107476 14408 107528 14414
rect 107476 14350 107528 14356
rect 107016 12980 107068 12986
rect 107016 12922 107068 12928
rect 107292 12980 107344 12986
rect 107292 12922 107344 12928
rect 106924 12844 106976 12850
rect 106924 12786 106976 12792
rect 106936 11540 106964 12786
rect 107028 12782 107056 12922
rect 107016 12776 107068 12782
rect 107016 12718 107068 12724
rect 107292 12436 107344 12442
rect 107292 12378 107344 12384
rect 107304 12322 107332 12378
rect 107212 12294 107332 12322
rect 107212 11626 107240 12294
rect 107292 12232 107344 12238
rect 107292 12174 107344 12180
rect 107304 11626 107332 12174
rect 107488 11762 107516 14350
rect 107856 13530 107884 15200
rect 107660 13524 107712 13530
rect 107660 13466 107712 13472
rect 107844 13524 107896 13530
rect 107844 13466 107896 13472
rect 107672 12646 107700 13466
rect 108408 12986 108436 15200
rect 108960 13530 108988 15200
rect 109316 14816 109368 14822
rect 109316 14758 109368 14764
rect 108948 13524 109000 13530
rect 108948 13466 109000 13472
rect 109040 13320 109092 13326
rect 109040 13262 109092 13268
rect 108580 13252 108632 13258
rect 108580 13194 108632 13200
rect 108396 12980 108448 12986
rect 108396 12922 108448 12928
rect 108120 12844 108172 12850
rect 108120 12786 108172 12792
rect 107660 12640 107712 12646
rect 107660 12582 107712 12588
rect 107568 12232 107620 12238
rect 107568 12174 107620 12180
rect 107476 11756 107528 11762
rect 107476 11698 107528 11704
rect 107200 11620 107252 11626
rect 107200 11562 107252 11568
rect 107292 11620 107344 11626
rect 107292 11562 107344 11568
rect 107016 11552 107068 11558
rect 106936 11512 107016 11540
rect 107016 11494 107068 11500
rect 107384 11552 107436 11558
rect 107384 11494 107436 11500
rect 106832 10260 106884 10266
rect 106832 10202 106884 10208
rect 106740 7812 106792 7818
rect 106740 7754 106792 7760
rect 107028 7342 107056 11494
rect 107396 11082 107424 11494
rect 107488 11354 107516 11698
rect 107580 11694 107608 12174
rect 107936 12096 107988 12102
rect 107936 12038 107988 12044
rect 108028 12096 108080 12102
rect 108028 12038 108080 12044
rect 107568 11688 107620 11694
rect 107568 11630 107620 11636
rect 107580 11354 107608 11630
rect 107476 11348 107528 11354
rect 107476 11290 107528 11296
rect 107568 11348 107620 11354
rect 107568 11290 107620 11296
rect 107384 11076 107436 11082
rect 107384 11018 107436 11024
rect 107580 10742 107608 11290
rect 107842 10840 107898 10849
rect 107752 10804 107804 10810
rect 107842 10775 107898 10784
rect 107752 10746 107804 10752
rect 107568 10736 107620 10742
rect 107764 10713 107792 10746
rect 107568 10678 107620 10684
rect 107750 10704 107806 10713
rect 107476 10668 107528 10674
rect 107476 10610 107528 10616
rect 107488 10538 107516 10610
rect 107476 10532 107528 10538
rect 107476 10474 107528 10480
rect 107580 10266 107608 10678
rect 107750 10639 107806 10648
rect 107856 10606 107884 10775
rect 107844 10600 107896 10606
rect 107764 10560 107844 10588
rect 107764 10266 107792 10560
rect 107844 10542 107896 10548
rect 107844 10464 107896 10470
rect 107844 10406 107896 10412
rect 107568 10260 107620 10266
rect 107568 10202 107620 10208
rect 107752 10260 107804 10266
rect 107752 10202 107804 10208
rect 107750 10160 107806 10169
rect 107476 10124 107528 10130
rect 107750 10095 107806 10104
rect 107476 10066 107528 10072
rect 107200 9376 107252 9382
rect 107200 9318 107252 9324
rect 107292 9376 107344 9382
rect 107292 9318 107344 9324
rect 107212 8974 107240 9318
rect 107200 8968 107252 8974
rect 107200 8910 107252 8916
rect 107304 8430 107332 9318
rect 107488 9110 107516 10066
rect 107764 9994 107792 10095
rect 107752 9988 107804 9994
rect 107752 9930 107804 9936
rect 107856 9761 107884 10406
rect 107842 9752 107898 9761
rect 107842 9687 107898 9696
rect 107844 9580 107896 9586
rect 107844 9522 107896 9528
rect 107660 9512 107712 9518
rect 107660 9454 107712 9460
rect 107476 9104 107528 9110
rect 107476 9046 107528 9052
rect 107568 8968 107620 8974
rect 107568 8910 107620 8916
rect 107580 8498 107608 8910
rect 107672 8673 107700 9454
rect 107856 8673 107884 9522
rect 107948 8906 107976 12038
rect 108040 9654 108068 12038
rect 108028 9648 108080 9654
rect 108028 9590 108080 9596
rect 107936 8900 107988 8906
rect 107936 8842 107988 8848
rect 107658 8664 107714 8673
rect 107658 8599 107714 8608
rect 107842 8664 107898 8673
rect 107842 8599 107898 8608
rect 107568 8492 107620 8498
rect 107568 8434 107620 8440
rect 107936 8492 107988 8498
rect 107936 8434 107988 8440
rect 107292 8424 107344 8430
rect 107292 8366 107344 8372
rect 107384 8424 107436 8430
rect 107384 8366 107436 8372
rect 107292 7812 107344 7818
rect 107292 7754 107344 7760
rect 107200 7744 107252 7750
rect 107200 7686 107252 7692
rect 107016 7336 107068 7342
rect 107016 7278 107068 7284
rect 106924 6860 106976 6866
rect 106924 6802 106976 6808
rect 106936 5953 106964 6802
rect 107016 6656 107068 6662
rect 107016 6598 107068 6604
rect 107028 6322 107056 6598
rect 107106 6488 107162 6497
rect 107106 6423 107162 6432
rect 107016 6316 107068 6322
rect 107016 6258 107068 6264
rect 107120 6254 107148 6423
rect 107212 6390 107240 7686
rect 107200 6384 107252 6390
rect 107200 6326 107252 6332
rect 107108 6248 107160 6254
rect 107108 6190 107160 6196
rect 106922 5944 106978 5953
rect 106922 5879 106978 5888
rect 106648 5840 106700 5846
rect 106648 5782 106700 5788
rect 106096 5772 106148 5778
rect 106096 5714 106148 5720
rect 105176 5228 105228 5234
rect 105176 5170 105228 5176
rect 104624 5160 104676 5166
rect 104624 5102 104676 5108
rect 104636 4826 104664 5102
rect 104624 4820 104676 4826
rect 104624 4762 104676 4768
rect 105188 4214 105216 5170
rect 105268 4616 105320 4622
rect 105268 4558 105320 4564
rect 105280 4214 105308 4558
rect 105176 4208 105228 4214
rect 105176 4150 105228 4156
rect 105268 4208 105320 4214
rect 105268 4150 105320 4156
rect 102968 3936 103020 3942
rect 102968 3878 103020 3884
rect 102048 3732 102100 3738
rect 102048 3674 102100 3680
rect 102980 3466 103008 3878
rect 105188 3602 105216 4150
rect 106556 4140 106608 4146
rect 106556 4082 106608 4088
rect 106004 3936 106056 3942
rect 106002 3904 106004 3913
rect 106056 3904 106058 3913
rect 106002 3839 106058 3848
rect 105176 3596 105228 3602
rect 105176 3538 105228 3544
rect 102968 3460 103020 3466
rect 102968 3402 103020 3408
rect 106464 3392 106516 3398
rect 106464 3334 106516 3340
rect 106476 2990 106504 3334
rect 106464 2984 106516 2990
rect 106464 2926 106516 2932
rect 106568 1970 106596 4082
rect 107304 2650 107332 7754
rect 107396 6730 107424 8366
rect 107948 8129 107976 8434
rect 107934 8120 107990 8129
rect 107934 8055 107990 8064
rect 107384 6724 107436 6730
rect 107384 6666 107436 6672
rect 107844 6384 107896 6390
rect 107396 6332 107844 6338
rect 107396 6326 107896 6332
rect 107396 6322 107884 6326
rect 107384 6316 107884 6322
rect 107436 6310 107884 6316
rect 107384 6258 107436 6264
rect 107672 5710 107700 6310
rect 107660 5704 107712 5710
rect 107382 5672 107438 5681
rect 107660 5646 107712 5652
rect 107382 5607 107384 5616
rect 107436 5607 107438 5616
rect 107384 5578 107436 5584
rect 108040 5574 108068 9590
rect 108028 5568 108080 5574
rect 108028 5510 108080 5516
rect 108132 4826 108160 12786
rect 108592 11150 108620 13194
rect 109052 12850 109080 13262
rect 109040 12844 109092 12850
rect 109040 12786 109092 12792
rect 108960 12714 109264 12730
rect 108948 12708 109264 12714
rect 109000 12702 109264 12708
rect 108948 12650 109000 12656
rect 109132 12640 109184 12646
rect 109052 12588 109132 12594
rect 109052 12582 109184 12588
rect 109052 12566 109172 12582
rect 109052 12434 109080 12566
rect 109052 12406 109172 12434
rect 108672 12368 108724 12374
rect 108672 12310 108724 12316
rect 108684 12220 108712 12310
rect 108684 12192 108896 12220
rect 108672 11892 108724 11898
rect 108672 11834 108724 11840
rect 108684 11694 108712 11834
rect 108868 11762 108896 12192
rect 108764 11756 108816 11762
rect 108764 11698 108816 11704
rect 108856 11756 108908 11762
rect 108856 11698 108908 11704
rect 108672 11688 108724 11694
rect 108672 11630 108724 11636
rect 108776 11354 108804 11698
rect 109040 11552 109092 11558
rect 109040 11494 109092 11500
rect 108764 11348 108816 11354
rect 108764 11290 108816 11296
rect 108304 11144 108356 11150
rect 108304 11086 108356 11092
rect 108580 11144 108632 11150
rect 108580 11086 108632 11092
rect 108212 10668 108264 10674
rect 108212 10610 108264 10616
rect 108224 9926 108252 10610
rect 108212 9920 108264 9926
rect 108212 9862 108264 9868
rect 108212 8832 108264 8838
rect 108212 8774 108264 8780
rect 108120 4820 108172 4826
rect 108120 4762 108172 4768
rect 107660 4004 107712 4010
rect 107660 3946 107712 3952
rect 107672 3058 107700 3946
rect 108224 3738 108252 8774
rect 108316 6746 108344 11086
rect 109052 11082 109080 11494
rect 109144 11150 109172 12406
rect 109236 11286 109264 12702
rect 109224 11280 109276 11286
rect 109224 11222 109276 11228
rect 109132 11144 109184 11150
rect 109132 11086 109184 11092
rect 109040 11076 109092 11082
rect 109040 11018 109092 11024
rect 109038 10840 109094 10849
rect 108948 10804 109000 10810
rect 109038 10775 109040 10784
rect 108948 10746 109000 10752
rect 109092 10775 109094 10784
rect 109040 10746 109092 10752
rect 108960 10690 108988 10746
rect 108960 10662 109080 10690
rect 108488 10464 108540 10470
rect 108488 10406 108540 10412
rect 108396 10056 108448 10062
rect 108396 9998 108448 10004
rect 108408 9450 108436 9998
rect 108396 9444 108448 9450
rect 108396 9386 108448 9392
rect 108408 6866 108436 9386
rect 108500 8498 108528 10406
rect 108672 9988 108724 9994
rect 108672 9930 108724 9936
rect 108684 9450 108712 9930
rect 108764 9920 108816 9926
rect 108764 9862 108816 9868
rect 108672 9444 108724 9450
rect 108672 9386 108724 9392
rect 108672 8560 108724 8566
rect 108672 8502 108724 8508
rect 108488 8492 108540 8498
rect 108488 8434 108540 8440
rect 108684 8294 108712 8502
rect 108672 8288 108724 8294
rect 108672 8230 108724 8236
rect 108396 6860 108448 6866
rect 108396 6802 108448 6808
rect 108316 6718 108436 6746
rect 108212 3732 108264 3738
rect 108212 3674 108264 3680
rect 108304 3392 108356 3398
rect 108304 3334 108356 3340
rect 108316 3126 108344 3334
rect 108408 3126 108436 6718
rect 108776 6458 108804 9862
rect 109052 9674 109080 10662
rect 109144 10606 109172 11086
rect 109132 10600 109184 10606
rect 109132 10542 109184 10548
rect 109052 9646 109264 9674
rect 109236 8906 109264 9646
rect 108948 8900 109000 8906
rect 108948 8842 109000 8848
rect 109224 8900 109276 8906
rect 109224 8842 109276 8848
rect 108854 7848 108910 7857
rect 108854 7783 108910 7792
rect 108868 7546 108896 7783
rect 108856 7540 108908 7546
rect 108856 7482 108908 7488
rect 108960 6934 108988 8842
rect 109132 8492 109184 8498
rect 109132 8434 109184 8440
rect 109144 7886 109172 8434
rect 109132 7880 109184 7886
rect 109132 7822 109184 7828
rect 108948 6928 109000 6934
rect 108948 6870 109000 6876
rect 108856 6860 108908 6866
rect 108856 6802 108908 6808
rect 108868 6458 108896 6802
rect 108764 6452 108816 6458
rect 108764 6394 108816 6400
rect 108856 6452 108908 6458
rect 108856 6394 108908 6400
rect 108868 5914 108896 6394
rect 108856 5908 108908 5914
rect 108856 5850 108908 5856
rect 108488 5772 108540 5778
rect 108488 5714 108540 5720
rect 108500 4622 108528 5714
rect 109144 5234 109172 7822
rect 109132 5228 109184 5234
rect 109132 5170 109184 5176
rect 108488 4616 108540 4622
rect 108488 4558 108540 4564
rect 109224 4548 109276 4554
rect 109224 4490 109276 4496
rect 109236 4457 109264 4490
rect 109222 4448 109278 4457
rect 109222 4383 109278 4392
rect 109328 4146 109356 14758
rect 109592 13728 109644 13734
rect 109592 13670 109644 13676
rect 109684 13728 109736 13734
rect 109684 13670 109736 13676
rect 109408 12912 109460 12918
rect 109408 12854 109460 12860
rect 109420 12646 109448 12854
rect 109408 12640 109460 12646
rect 109408 12582 109460 12588
rect 109408 12164 109460 12170
rect 109408 12106 109460 12112
rect 109420 5794 109448 12106
rect 109604 11354 109632 13670
rect 109696 13326 109724 13670
rect 109788 13462 109816 15286
rect 110050 15286 110276 15314
rect 110050 15200 110106 15286
rect 109776 13456 109828 13462
rect 109776 13398 109828 13404
rect 109684 13320 109736 13326
rect 109684 13262 109736 13268
rect 110052 13320 110104 13326
rect 110052 13262 110104 13268
rect 109684 11892 109736 11898
rect 109684 11834 109736 11840
rect 109696 11558 109724 11834
rect 109684 11552 109736 11558
rect 109684 11494 109736 11500
rect 109592 11348 109644 11354
rect 109592 11290 109644 11296
rect 109592 11144 109644 11150
rect 109592 11086 109644 11092
rect 109604 8498 109632 11086
rect 109592 8492 109644 8498
rect 109592 8434 109644 8440
rect 109420 5766 109540 5794
rect 109512 4826 109540 5766
rect 109500 4820 109552 4826
rect 109500 4762 109552 4768
rect 109316 4140 109368 4146
rect 109316 4082 109368 4088
rect 109040 4072 109092 4078
rect 109040 4014 109092 4020
rect 109052 3534 109080 4014
rect 109040 3528 109092 3534
rect 109040 3470 109092 3476
rect 109328 3194 109356 4082
rect 109696 4010 109724 11494
rect 110064 9382 110092 13262
rect 110248 12442 110276 15286
rect 110602 15200 110658 16000
rect 111154 15314 111210 16000
rect 111154 15286 111472 15314
rect 111154 15200 111210 15286
rect 110616 13530 110644 15200
rect 110604 13524 110656 13530
rect 110604 13466 110656 13472
rect 111444 13462 111472 15286
rect 111706 15200 111762 16000
rect 112258 15200 112314 16000
rect 112810 15200 112866 16000
rect 113362 15314 113418 16000
rect 113362 15286 113680 15314
rect 113362 15200 113418 15286
rect 111432 13456 111484 13462
rect 111432 13398 111484 13404
rect 110512 13388 110564 13394
rect 110512 13330 110564 13336
rect 110420 13184 110472 13190
rect 110418 13152 110420 13161
rect 110472 13152 110474 13161
rect 110418 13087 110474 13096
rect 110328 12708 110380 12714
rect 110328 12650 110380 12656
rect 110236 12436 110288 12442
rect 110236 12378 110288 12384
rect 110340 9994 110368 12650
rect 110420 12640 110472 12646
rect 110420 12582 110472 12588
rect 110432 12481 110460 12582
rect 110418 12472 110474 12481
rect 110418 12407 110474 12416
rect 110420 11552 110472 11558
rect 110420 11494 110472 11500
rect 110432 11082 110460 11494
rect 110420 11076 110472 11082
rect 110420 11018 110472 11024
rect 110420 10600 110472 10606
rect 110420 10542 110472 10548
rect 110432 10062 110460 10542
rect 110420 10056 110472 10062
rect 110420 9998 110472 10004
rect 110328 9988 110380 9994
rect 110328 9930 110380 9936
rect 110052 9376 110104 9382
rect 110052 9318 110104 9324
rect 110064 8265 110092 9318
rect 110050 8256 110106 8265
rect 110050 8191 110106 8200
rect 110524 8106 110552 13330
rect 111340 13320 111392 13326
rect 111340 13262 111392 13268
rect 111352 12646 111380 13262
rect 110972 12640 111024 12646
rect 110972 12582 111024 12588
rect 111340 12640 111392 12646
rect 111340 12582 111392 12588
rect 110880 12232 110932 12238
rect 110880 12174 110932 12180
rect 110892 10810 110920 12174
rect 110604 10804 110656 10810
rect 110604 10746 110656 10752
rect 110880 10804 110932 10810
rect 110880 10746 110932 10752
rect 110616 10674 110644 10746
rect 110984 10674 111012 12582
rect 111720 12442 111748 15200
rect 112272 12986 112300 15200
rect 112824 13530 112852 15200
rect 112812 13524 112864 13530
rect 112812 13466 112864 13472
rect 112824 13394 113036 13410
rect 112824 13388 113048 13394
rect 112824 13382 112996 13388
rect 112444 13320 112496 13326
rect 112496 13268 112668 13274
rect 112444 13262 112668 13268
rect 112456 13258 112668 13262
rect 112456 13252 112680 13258
rect 112456 13246 112628 13252
rect 112628 13194 112680 13200
rect 112260 12980 112312 12986
rect 112260 12922 112312 12928
rect 112444 12776 112496 12782
rect 112444 12718 112496 12724
rect 111708 12436 111760 12442
rect 111708 12378 111760 12384
rect 112352 12436 112404 12442
rect 112456 12434 112484 12718
rect 112456 12406 112576 12434
rect 112352 12378 112404 12384
rect 111248 12232 111300 12238
rect 111248 12174 111300 12180
rect 111064 12096 111116 12102
rect 111064 12038 111116 12044
rect 111076 11218 111104 12038
rect 111156 11280 111208 11286
rect 111156 11222 111208 11228
rect 111064 11212 111116 11218
rect 111064 11154 111116 11160
rect 111064 11008 111116 11014
rect 111064 10950 111116 10956
rect 110604 10668 110656 10674
rect 110604 10610 110656 10616
rect 110880 10668 110932 10674
rect 110880 10610 110932 10616
rect 110972 10668 111024 10674
rect 110972 10610 111024 10616
rect 110696 10600 110748 10606
rect 110696 10542 110748 10548
rect 110604 10464 110656 10470
rect 110708 10452 110736 10542
rect 110656 10424 110736 10452
rect 110788 10464 110840 10470
rect 110604 10406 110656 10412
rect 110788 10406 110840 10412
rect 110696 10192 110748 10198
rect 110696 10134 110748 10140
rect 110604 10056 110656 10062
rect 110604 9998 110656 10004
rect 110432 8078 110552 8106
rect 110432 8022 110460 8078
rect 110420 8016 110472 8022
rect 110420 7958 110472 7964
rect 109776 7812 109828 7818
rect 109776 7754 109828 7760
rect 109868 7812 109920 7818
rect 109868 7754 109920 7760
rect 109788 7018 109816 7754
rect 109880 7206 109908 7754
rect 110616 7478 110644 9998
rect 110708 9926 110736 10134
rect 110696 9920 110748 9926
rect 110696 9862 110748 9868
rect 110800 9586 110828 10406
rect 110892 9926 110920 10610
rect 111076 10554 111104 10950
rect 110984 10526 111104 10554
rect 110880 9920 110932 9926
rect 110880 9862 110932 9868
rect 110788 9580 110840 9586
rect 110788 9522 110840 9528
rect 110788 9376 110840 9382
rect 110788 9318 110840 9324
rect 110800 8838 110828 9318
rect 110788 8832 110840 8838
rect 110788 8774 110840 8780
rect 110696 7744 110748 7750
rect 110696 7686 110748 7692
rect 110604 7472 110656 7478
rect 110604 7414 110656 7420
rect 110326 7304 110382 7313
rect 110326 7239 110328 7248
rect 110380 7239 110382 7248
rect 110328 7210 110380 7216
rect 109868 7200 109920 7206
rect 109868 7142 109920 7148
rect 110052 7200 110104 7206
rect 110052 7142 110104 7148
rect 110064 7018 110092 7142
rect 110616 7041 110644 7414
rect 110708 7410 110736 7686
rect 110696 7404 110748 7410
rect 110696 7346 110748 7352
rect 109788 6990 110092 7018
rect 109776 5228 109828 5234
rect 109776 5170 109828 5176
rect 109788 4622 109816 5170
rect 109776 4616 109828 4622
rect 109776 4558 109828 4564
rect 109684 4004 109736 4010
rect 109684 3946 109736 3952
rect 110064 3534 110092 6990
rect 110602 7032 110658 7041
rect 110602 6967 110658 6976
rect 110616 6934 110644 6967
rect 110604 6928 110656 6934
rect 110604 6870 110656 6876
rect 110604 6792 110656 6798
rect 110604 6734 110656 6740
rect 110696 6792 110748 6798
rect 110696 6734 110748 6740
rect 110616 6633 110644 6734
rect 110602 6624 110658 6633
rect 110602 6559 110658 6568
rect 110708 6390 110736 6734
rect 110696 6384 110748 6390
rect 110696 6326 110748 6332
rect 110892 5166 110920 9862
rect 110984 9382 111012 10526
rect 110972 9376 111024 9382
rect 110972 9318 111024 9324
rect 110972 7880 111024 7886
rect 110972 7822 111024 7828
rect 111064 7880 111116 7886
rect 111064 7822 111116 7828
rect 110984 7342 111012 7822
rect 110972 7336 111024 7342
rect 110972 7278 111024 7284
rect 111076 6934 111104 7822
rect 111064 6928 111116 6934
rect 111064 6870 111116 6876
rect 110880 5160 110932 5166
rect 110880 5102 110932 5108
rect 110328 4276 110380 4282
rect 110328 4218 110380 4224
rect 109592 3528 109644 3534
rect 109592 3470 109644 3476
rect 110052 3528 110104 3534
rect 110052 3470 110104 3476
rect 109316 3188 109368 3194
rect 109316 3130 109368 3136
rect 108304 3120 108356 3126
rect 108304 3062 108356 3068
rect 108396 3120 108448 3126
rect 108396 3062 108448 3068
rect 107660 3052 107712 3058
rect 107660 2994 107712 3000
rect 107292 2644 107344 2650
rect 107292 2586 107344 2592
rect 108316 2009 108344 3062
rect 109604 2650 109632 3470
rect 110144 3460 110196 3466
rect 110144 3402 110196 3408
rect 110052 3392 110104 3398
rect 110052 3334 110104 3340
rect 110064 2922 110092 3334
rect 110156 3194 110184 3402
rect 110144 3188 110196 3194
rect 110144 3130 110196 3136
rect 110052 2916 110104 2922
rect 110052 2858 110104 2864
rect 110156 2774 110184 3130
rect 110340 2922 110368 4218
rect 111168 4146 111196 11222
rect 111260 11014 111288 12174
rect 111616 12096 111668 12102
rect 111616 12038 111668 12044
rect 111628 11150 111656 12038
rect 112364 11898 112392 12378
rect 112548 12170 112576 12406
rect 112536 12164 112588 12170
rect 112536 12106 112588 12112
rect 112352 11892 112404 11898
rect 112352 11834 112404 11840
rect 112076 11756 112128 11762
rect 112076 11698 112128 11704
rect 112168 11756 112220 11762
rect 112168 11698 112220 11704
rect 112088 11354 112116 11698
rect 112076 11348 112128 11354
rect 112076 11290 112128 11296
rect 111616 11144 111668 11150
rect 111616 11086 111668 11092
rect 112180 11082 112208 11698
rect 112548 11626 112576 12106
rect 112536 11620 112588 11626
rect 112536 11562 112588 11568
rect 111708 11076 111760 11082
rect 111708 11018 111760 11024
rect 112168 11076 112220 11082
rect 112168 11018 112220 11024
rect 111248 11008 111300 11014
rect 111248 10950 111300 10956
rect 111260 10198 111288 10950
rect 111524 10804 111576 10810
rect 111524 10746 111576 10752
rect 111536 10674 111564 10746
rect 111432 10668 111484 10674
rect 111432 10610 111484 10616
rect 111524 10668 111576 10674
rect 111720 10656 111748 11018
rect 111800 10668 111852 10674
rect 111720 10628 111800 10656
rect 111524 10610 111576 10616
rect 111800 10610 111852 10616
rect 111444 10470 111472 10610
rect 111340 10464 111392 10470
rect 111340 10406 111392 10412
rect 111432 10464 111484 10470
rect 111432 10406 111484 10412
rect 111248 10192 111300 10198
rect 111248 10134 111300 10140
rect 111248 9376 111300 9382
rect 111248 9318 111300 9324
rect 111156 4140 111208 4146
rect 111156 4082 111208 4088
rect 110972 4072 111024 4078
rect 110972 4014 111024 4020
rect 110984 3602 111012 4014
rect 110972 3596 111024 3602
rect 110972 3538 111024 3544
rect 110328 2916 110380 2922
rect 110328 2858 110380 2864
rect 110156 2746 110276 2774
rect 109592 2644 109644 2650
rect 109592 2586 109644 2592
rect 108302 2000 108358 2009
rect 106556 1964 106608 1970
rect 108302 1935 108358 1944
rect 106556 1906 106608 1912
rect 110248 1358 110276 2746
rect 111260 2446 111288 9318
rect 111352 8974 111380 10406
rect 111536 10062 111564 10610
rect 111616 10532 111668 10538
rect 111616 10474 111668 10480
rect 111628 10169 111656 10474
rect 111614 10160 111670 10169
rect 111614 10095 111670 10104
rect 111524 10056 111576 10062
rect 111524 9998 111576 10004
rect 111616 10056 111668 10062
rect 111616 9998 111668 10004
rect 111340 8968 111392 8974
rect 111340 8910 111392 8916
rect 111628 7478 111656 9998
rect 112076 8288 112128 8294
rect 112076 8230 112128 8236
rect 112088 8090 112116 8230
rect 112180 8090 112208 11018
rect 112548 10266 112576 11562
rect 112720 11552 112772 11558
rect 112720 11494 112772 11500
rect 112732 10810 112760 11494
rect 112720 10804 112772 10810
rect 112720 10746 112772 10752
rect 112536 10260 112588 10266
rect 112536 10202 112588 10208
rect 112626 9616 112682 9625
rect 112626 9551 112682 9560
rect 112352 8968 112404 8974
rect 112352 8910 112404 8916
rect 112364 8566 112392 8910
rect 112352 8560 112404 8566
rect 112352 8502 112404 8508
rect 112534 8120 112590 8129
rect 112076 8084 112128 8090
rect 112076 8026 112128 8032
rect 112168 8084 112220 8090
rect 112534 8055 112590 8064
rect 112168 8026 112220 8032
rect 111616 7472 111668 7478
rect 111616 7414 111668 7420
rect 111340 7336 111392 7342
rect 111340 7278 111392 7284
rect 111352 6934 111380 7278
rect 111340 6928 111392 6934
rect 111340 6870 111392 6876
rect 111524 6928 111576 6934
rect 111524 6870 111576 6876
rect 111352 6458 111380 6870
rect 111432 6792 111484 6798
rect 111432 6734 111484 6740
rect 111340 6452 111392 6458
rect 111340 6394 111392 6400
rect 111444 6390 111472 6734
rect 111432 6384 111484 6390
rect 111432 6326 111484 6332
rect 111536 2854 111564 6870
rect 111616 6724 111668 6730
rect 111616 6666 111668 6672
rect 111628 6458 111656 6666
rect 111616 6452 111668 6458
rect 111616 6394 111668 6400
rect 111984 6384 112036 6390
rect 111984 6326 112036 6332
rect 111892 6112 111944 6118
rect 111892 6054 111944 6060
rect 111904 5098 111932 6054
rect 111996 5953 112024 6326
rect 111982 5944 112038 5953
rect 111982 5879 112038 5888
rect 112180 5642 112208 8026
rect 112548 8022 112576 8055
rect 112536 8016 112588 8022
rect 112536 7958 112588 7964
rect 112444 7336 112496 7342
rect 112442 7304 112444 7313
rect 112640 7313 112668 9551
rect 112720 8492 112772 8498
rect 112720 8434 112772 8440
rect 112732 7886 112760 8434
rect 112824 8362 112852 13382
rect 112996 13330 113048 13336
rect 112996 13252 113048 13258
rect 112996 13194 113048 13200
rect 113088 13252 113140 13258
rect 113088 13194 113140 13200
rect 113008 12434 113036 13194
rect 113100 13161 113128 13194
rect 113180 13184 113232 13190
rect 113086 13152 113142 13161
rect 113180 13126 113232 13132
rect 113086 13087 113142 13096
rect 113008 12406 113128 12434
rect 112904 10804 112956 10810
rect 112904 10746 112956 10752
rect 112916 10062 112944 10746
rect 112996 10192 113048 10198
rect 112996 10134 113048 10140
rect 112904 10056 112956 10062
rect 112904 9998 112956 10004
rect 112812 8356 112864 8362
rect 112812 8298 112864 8304
rect 112720 7880 112772 7886
rect 112720 7822 112772 7828
rect 112904 7880 112956 7886
rect 112904 7822 112956 7828
rect 112916 7342 112944 7822
rect 113008 7818 113036 10134
rect 113100 9926 113128 12406
rect 113192 11218 113220 13126
rect 113652 12986 113680 15286
rect 113914 15200 113970 16000
rect 114466 15200 114522 16000
rect 115018 15314 115074 16000
rect 115018 15286 115244 15314
rect 115018 15200 115074 15286
rect 113928 13530 113956 15200
rect 114192 14748 114244 14754
rect 114192 14690 114244 14696
rect 113916 13524 113968 13530
rect 113916 13466 113968 13472
rect 113640 12980 113692 12986
rect 113640 12922 113692 12928
rect 113272 12912 113324 12918
rect 113272 12854 113324 12860
rect 113284 11898 113312 12854
rect 113548 12776 113600 12782
rect 113548 12718 113600 12724
rect 113560 12102 113588 12718
rect 113548 12096 113600 12102
rect 113548 12038 113600 12044
rect 113272 11892 113324 11898
rect 113272 11834 113324 11840
rect 113180 11212 113232 11218
rect 113180 11154 113232 11160
rect 113364 11212 113416 11218
rect 113364 11154 113416 11160
rect 113088 9920 113140 9926
rect 113086 9888 113088 9897
rect 113140 9888 113142 9897
rect 113086 9823 113142 9832
rect 113272 9512 113324 9518
rect 113272 9454 113324 9460
rect 113284 8838 113312 9454
rect 113272 8832 113324 8838
rect 113272 8774 113324 8780
rect 113376 8129 113404 11154
rect 113454 10704 113510 10713
rect 113454 10639 113510 10648
rect 113468 10470 113496 10639
rect 113456 10464 113508 10470
rect 113456 10406 113508 10412
rect 113560 10169 113588 12038
rect 113640 11756 113692 11762
rect 113640 11698 113692 11704
rect 113546 10160 113602 10169
rect 113546 10095 113602 10104
rect 113548 10056 113600 10062
rect 113548 9998 113600 10004
rect 113560 9926 113588 9998
rect 113548 9920 113600 9926
rect 113548 9862 113600 9868
rect 113560 9722 113588 9862
rect 113548 9716 113600 9722
rect 113548 9658 113600 9664
rect 113362 8120 113418 8129
rect 113362 8055 113418 8064
rect 113088 7880 113140 7886
rect 113088 7822 113140 7828
rect 113270 7848 113326 7857
rect 112996 7812 113048 7818
rect 112996 7754 113048 7760
rect 112904 7336 112956 7342
rect 112496 7304 112498 7313
rect 112442 7239 112498 7248
rect 112626 7304 112682 7313
rect 112904 7278 112956 7284
rect 112626 7239 112682 7248
rect 112720 7200 112772 7206
rect 112720 7142 112772 7148
rect 112904 7200 112956 7206
rect 112904 7142 112956 7148
rect 112168 5636 112220 5642
rect 112168 5578 112220 5584
rect 111892 5092 111944 5098
rect 111892 5034 111944 5040
rect 112168 5024 112220 5030
rect 112168 4966 112220 4972
rect 112180 4486 112208 4966
rect 112168 4480 112220 4486
rect 112168 4422 112220 4428
rect 112732 4185 112760 7142
rect 112916 6934 112944 7142
rect 112904 6928 112956 6934
rect 112904 6870 112956 6876
rect 113100 6866 113128 7822
rect 113270 7783 113326 7792
rect 113284 7342 113312 7783
rect 113272 7336 113324 7342
rect 113272 7278 113324 7284
rect 113088 6860 113140 6866
rect 113088 6802 113140 6808
rect 113548 5568 113600 5574
rect 113548 5510 113600 5516
rect 113560 5166 113588 5510
rect 113548 5160 113600 5166
rect 113548 5102 113600 5108
rect 113548 4480 113600 4486
rect 113548 4422 113600 4428
rect 112718 4176 112774 4185
rect 112718 4111 112774 4120
rect 111616 4004 111668 4010
rect 111616 3946 111668 3952
rect 111628 3398 111656 3946
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111524 2848 111576 2854
rect 111524 2790 111576 2796
rect 112732 2650 112760 4111
rect 112720 2644 112772 2650
rect 112720 2586 112772 2592
rect 111248 2440 111300 2446
rect 111248 2382 111300 2388
rect 110236 1352 110288 1358
rect 110236 1294 110288 1300
rect 101956 1080 102008 1086
rect 101956 1022 102008 1028
rect 113560 1018 113588 4422
rect 113652 2650 113680 11698
rect 113824 11348 113876 11354
rect 113824 11290 113876 11296
rect 113732 10668 113784 10674
rect 113732 10610 113784 10616
rect 113744 9722 113772 10610
rect 113836 10470 113864 11290
rect 113824 10464 113876 10470
rect 113824 10406 113876 10412
rect 113916 9988 113968 9994
rect 113916 9930 113968 9936
rect 113732 9716 113784 9722
rect 113732 9658 113784 9664
rect 113824 9648 113876 9654
rect 113824 9590 113876 9596
rect 113836 9518 113864 9590
rect 113824 9512 113876 9518
rect 113824 9454 113876 9460
rect 113824 6112 113876 6118
rect 113824 6054 113876 6060
rect 113732 5704 113784 5710
rect 113730 5672 113732 5681
rect 113784 5672 113786 5681
rect 113730 5607 113786 5616
rect 113732 5568 113784 5574
rect 113732 5510 113784 5516
rect 113744 4690 113772 5510
rect 113836 5234 113864 6054
rect 113824 5228 113876 5234
rect 113824 5170 113876 5176
rect 113732 4684 113784 4690
rect 113732 4626 113784 4632
rect 113732 4276 113784 4282
rect 113732 4218 113784 4224
rect 113744 4078 113772 4218
rect 113732 4072 113784 4078
rect 113732 4014 113784 4020
rect 113928 3738 113956 9930
rect 114100 9920 114152 9926
rect 114100 9862 114152 9868
rect 114008 9376 114060 9382
rect 114008 9318 114060 9324
rect 114020 6769 114048 9318
rect 114112 7410 114140 9862
rect 114204 9382 114232 14690
rect 114480 13462 114508 15200
rect 114468 13456 114520 13462
rect 114468 13398 114520 13404
rect 114468 13320 114520 13326
rect 114468 13262 114520 13268
rect 114652 13320 114704 13326
rect 114652 13262 114704 13268
rect 114480 12714 114508 13262
rect 114468 12708 114520 12714
rect 114468 12650 114520 12656
rect 114560 12640 114612 12646
rect 114560 12582 114612 12588
rect 114284 12300 114336 12306
rect 114284 12242 114336 12248
rect 114296 12102 114324 12242
rect 114572 12102 114600 12582
rect 114284 12096 114336 12102
rect 114284 12038 114336 12044
rect 114560 12096 114612 12102
rect 114560 12038 114612 12044
rect 114192 9376 114244 9382
rect 114192 9318 114244 9324
rect 114192 8424 114244 8430
rect 114192 8366 114244 8372
rect 114100 7404 114152 7410
rect 114100 7346 114152 7352
rect 114006 6760 114062 6769
rect 114006 6695 114062 6704
rect 114100 5364 114152 5370
rect 114100 5306 114152 5312
rect 114112 4622 114140 5306
rect 114100 4616 114152 4622
rect 114100 4558 114152 4564
rect 114204 4214 114232 8366
rect 114192 4208 114244 4214
rect 114192 4150 114244 4156
rect 113916 3732 113968 3738
rect 113916 3674 113968 3680
rect 113640 2644 113692 2650
rect 113640 2586 113692 2592
rect 114296 1737 114324 12038
rect 114572 11354 114600 12038
rect 114560 11348 114612 11354
rect 114560 11290 114612 11296
rect 114560 10668 114612 10674
rect 114560 10610 114612 10616
rect 114468 9172 114520 9178
rect 114468 9114 114520 9120
rect 114480 8809 114508 9114
rect 114466 8800 114522 8809
rect 114466 8735 114522 8744
rect 114466 7032 114522 7041
rect 114466 6967 114522 6976
rect 114480 6934 114508 6967
rect 114468 6928 114520 6934
rect 114468 6870 114520 6876
rect 114480 2650 114508 6870
rect 114572 6866 114600 10610
rect 114560 6860 114612 6866
rect 114560 6802 114612 6808
rect 114560 6316 114612 6322
rect 114560 6258 114612 6264
rect 114572 5846 114600 6258
rect 114664 6186 114692 13262
rect 114744 13184 114796 13190
rect 114744 13126 114796 13132
rect 114756 12782 114784 13126
rect 114744 12776 114796 12782
rect 114744 12718 114796 12724
rect 114836 12232 114888 12238
rect 114836 12174 114888 12180
rect 114848 11898 114876 12174
rect 115216 12102 115244 15286
rect 115570 15200 115626 16000
rect 116122 15314 116178 16000
rect 116122 15286 116348 15314
rect 116122 15200 116178 15286
rect 115584 13530 115612 15200
rect 115664 13796 115716 13802
rect 115664 13738 115716 13744
rect 115572 13524 115624 13530
rect 115572 13466 115624 13472
rect 115676 13326 115704 13738
rect 115664 13320 115716 13326
rect 115664 13262 115716 13268
rect 115676 12968 115704 13262
rect 115676 12940 115888 12968
rect 115662 12880 115718 12889
rect 115860 12850 115888 12940
rect 115662 12815 115718 12824
rect 115756 12844 115808 12850
rect 115296 12164 115348 12170
rect 115296 12106 115348 12112
rect 115204 12096 115256 12102
rect 115204 12038 115256 12044
rect 114836 11892 114888 11898
rect 114836 11834 114888 11840
rect 115204 11348 115256 11354
rect 115204 11290 115256 11296
rect 114744 10056 114796 10062
rect 114744 9998 114796 10004
rect 114756 9518 114784 9998
rect 114926 9616 114982 9625
rect 114926 9551 114982 9560
rect 114744 9512 114796 9518
rect 114744 9454 114796 9460
rect 114756 7834 114784 9454
rect 114940 9178 114968 9551
rect 114928 9172 114980 9178
rect 114928 9114 114980 9120
rect 114756 7806 114968 7834
rect 114836 7744 114888 7750
rect 114742 7712 114798 7721
rect 114836 7686 114888 7692
rect 114742 7647 114798 7656
rect 114756 6769 114784 7647
rect 114848 6798 114876 7686
rect 114940 7206 114968 7806
rect 114928 7200 114980 7206
rect 114928 7142 114980 7148
rect 114836 6792 114888 6798
rect 114742 6760 114798 6769
rect 114836 6734 114888 6740
rect 114742 6695 114798 6704
rect 114652 6180 114704 6186
rect 114652 6122 114704 6128
rect 114848 6066 114876 6734
rect 114940 6322 114968 7142
rect 115020 6792 115072 6798
rect 115020 6734 115072 6740
rect 115032 6662 115060 6734
rect 115020 6656 115072 6662
rect 115020 6598 115072 6604
rect 114928 6316 114980 6322
rect 114928 6258 114980 6264
rect 114848 6038 115152 6066
rect 114560 5840 114612 5846
rect 114560 5782 114612 5788
rect 115124 4758 115152 6038
rect 115112 4752 115164 4758
rect 115112 4694 115164 4700
rect 114652 4548 114704 4554
rect 114652 4490 114704 4496
rect 114664 4146 114692 4490
rect 114652 4140 114704 4146
rect 114652 4082 114704 4088
rect 114836 3392 114888 3398
rect 114836 3334 114888 3340
rect 114848 3194 114876 3334
rect 114836 3188 114888 3194
rect 114836 3130 114888 3136
rect 114848 3058 114876 3130
rect 114836 3052 114888 3058
rect 114836 2994 114888 3000
rect 114468 2644 114520 2650
rect 114468 2586 114520 2592
rect 114480 1834 114508 2586
rect 114468 1828 114520 1834
rect 114468 1770 114520 1776
rect 114282 1728 114338 1737
rect 114282 1663 114338 1672
rect 115216 1290 115244 11290
rect 115308 11218 115336 12106
rect 115676 11762 115704 12815
rect 115756 12786 115808 12792
rect 115848 12844 115900 12850
rect 115848 12786 115900 12792
rect 115664 11756 115716 11762
rect 115664 11698 115716 11704
rect 115480 11688 115532 11694
rect 115480 11630 115532 11636
rect 115492 11286 115520 11630
rect 115480 11280 115532 11286
rect 115480 11222 115532 11228
rect 115296 11212 115348 11218
rect 115296 11154 115348 11160
rect 115308 10810 115336 11154
rect 115388 11076 115440 11082
rect 115388 11018 115440 11024
rect 115296 10804 115348 10810
rect 115296 10746 115348 10752
rect 115400 9518 115428 11018
rect 115676 10810 115704 11698
rect 115768 11218 115796 12786
rect 116124 12640 116176 12646
rect 116122 12608 116124 12617
rect 116176 12608 116178 12617
rect 116122 12543 116178 12552
rect 116320 12102 116348 15286
rect 116674 15200 116730 16000
rect 117226 15200 117282 16000
rect 117778 15200 117834 16000
rect 118330 15200 118386 16000
rect 118882 15314 118938 16000
rect 119434 15314 119490 16000
rect 118882 15286 119200 15314
rect 118882 15200 118938 15286
rect 116688 13530 116716 15200
rect 116950 13696 117006 13705
rect 116950 13631 117006 13640
rect 116676 13524 116728 13530
rect 116676 13466 116728 13472
rect 116584 13320 116636 13326
rect 116584 13262 116636 13268
rect 116596 12850 116624 13262
rect 116584 12844 116636 12850
rect 116584 12786 116636 12792
rect 116964 12434 116992 13631
rect 117240 13394 117268 15200
rect 117228 13388 117280 13394
rect 117228 13330 117280 13336
rect 117320 13320 117372 13326
rect 117148 13268 117320 13274
rect 117148 13262 117372 13268
rect 117148 13258 117360 13262
rect 117136 13252 117360 13258
rect 117188 13246 117360 13252
rect 117136 13194 117188 13200
rect 117320 13184 117372 13190
rect 117320 13126 117372 13132
rect 116872 12406 116992 12434
rect 117332 12434 117360 13126
rect 117792 12986 117820 15200
rect 118056 14884 118108 14890
rect 118056 14826 118108 14832
rect 117964 13388 118016 13394
rect 117964 13330 118016 13336
rect 117688 12980 117740 12986
rect 117688 12922 117740 12928
rect 117780 12980 117832 12986
rect 117780 12922 117832 12928
rect 117332 12406 117452 12434
rect 116492 12232 116544 12238
rect 116492 12174 116544 12180
rect 116308 12096 116360 12102
rect 116308 12038 116360 12044
rect 116400 12096 116452 12102
rect 116504 12073 116532 12174
rect 116400 12038 116452 12044
rect 116490 12064 116546 12073
rect 116412 11762 116440 12038
rect 116490 11999 116546 12008
rect 116400 11756 116452 11762
rect 116400 11698 116452 11704
rect 115848 11552 115900 11558
rect 115848 11494 115900 11500
rect 115860 11218 115888 11494
rect 115940 11280 115992 11286
rect 115940 11222 115992 11228
rect 116584 11280 116636 11286
rect 116584 11222 116636 11228
rect 115756 11212 115808 11218
rect 115756 11154 115808 11160
rect 115848 11212 115900 11218
rect 115848 11154 115900 11160
rect 115664 10804 115716 10810
rect 115664 10746 115716 10752
rect 115664 10600 115716 10606
rect 115664 10542 115716 10548
rect 115572 10124 115624 10130
rect 115572 10066 115624 10072
rect 115584 9926 115612 10066
rect 115480 9920 115532 9926
rect 115480 9862 115532 9868
rect 115572 9920 115624 9926
rect 115572 9862 115624 9868
rect 115388 9512 115440 9518
rect 115388 9454 115440 9460
rect 115388 9376 115440 9382
rect 115388 9318 115440 9324
rect 115294 9208 115350 9217
rect 115294 9143 115350 9152
rect 115308 8566 115336 9143
rect 115296 8560 115348 8566
rect 115296 8502 115348 8508
rect 115294 8392 115350 8401
rect 115400 8378 115428 9318
rect 115350 8350 115428 8378
rect 115294 8327 115350 8336
rect 115308 4049 115336 8327
rect 115492 7818 115520 9862
rect 115570 9344 115626 9353
rect 115570 9279 115626 9288
rect 115584 9178 115612 9279
rect 115572 9172 115624 9178
rect 115572 9114 115624 9120
rect 115570 8664 115626 8673
rect 115570 8599 115626 8608
rect 115584 8498 115612 8599
rect 115572 8492 115624 8498
rect 115572 8434 115624 8440
rect 115480 7812 115532 7818
rect 115480 7754 115532 7760
rect 115480 6860 115532 6866
rect 115480 6802 115532 6808
rect 115388 6724 115440 6730
rect 115388 6666 115440 6672
rect 115400 6497 115428 6666
rect 115492 6633 115520 6802
rect 115478 6624 115534 6633
rect 115478 6559 115534 6568
rect 115386 6488 115442 6497
rect 115386 6423 115442 6432
rect 115386 6352 115442 6361
rect 115386 6287 115442 6296
rect 115400 5846 115428 6287
rect 115388 5840 115440 5846
rect 115388 5782 115440 5788
rect 115400 5681 115428 5782
rect 115386 5672 115442 5681
rect 115386 5607 115442 5616
rect 115480 5024 115532 5030
rect 115480 4966 115532 4972
rect 115388 4548 115440 4554
rect 115388 4490 115440 4496
rect 115400 4457 115428 4490
rect 115386 4448 115442 4457
rect 115386 4383 115442 4392
rect 115294 4040 115350 4049
rect 115294 3975 115350 3984
rect 115492 3058 115520 4966
rect 115572 4480 115624 4486
rect 115572 4422 115624 4428
rect 115584 4146 115612 4422
rect 115572 4140 115624 4146
rect 115572 4082 115624 4088
rect 115480 3052 115532 3058
rect 115480 2994 115532 3000
rect 115584 1698 115612 4082
rect 115676 3194 115704 10542
rect 115768 4146 115796 11154
rect 115952 11014 115980 11222
rect 115940 11008 115992 11014
rect 115940 10950 115992 10956
rect 116308 11008 116360 11014
rect 116308 10950 116360 10956
rect 115848 10464 115900 10470
rect 115848 10406 115900 10412
rect 115860 10130 115888 10406
rect 115848 10124 115900 10130
rect 115848 10066 115900 10072
rect 115952 10062 115980 10950
rect 116030 10840 116086 10849
rect 116030 10775 116086 10784
rect 116216 10804 116268 10810
rect 115940 10056 115992 10062
rect 115940 9998 115992 10004
rect 115848 9988 115900 9994
rect 115848 9930 115900 9936
rect 115860 9761 115888 9930
rect 115846 9752 115902 9761
rect 115846 9687 115902 9696
rect 115848 9512 115900 9518
rect 115848 9454 115900 9460
rect 115860 9178 115888 9454
rect 115848 9172 115900 9178
rect 115848 9114 115900 9120
rect 115952 9058 115980 9998
rect 116044 9994 116072 10775
rect 116216 10746 116268 10752
rect 116228 10606 116256 10746
rect 116216 10600 116268 10606
rect 116216 10542 116268 10548
rect 116032 9988 116084 9994
rect 116032 9930 116084 9936
rect 116320 9654 116348 10950
rect 116596 9654 116624 11222
rect 116308 9648 116360 9654
rect 116308 9590 116360 9596
rect 116584 9648 116636 9654
rect 116584 9590 116636 9596
rect 115860 9030 116072 9058
rect 115860 8838 115888 9030
rect 115848 8832 115900 8838
rect 115848 8774 115900 8780
rect 115938 8528 115994 8537
rect 115938 8463 115994 8472
rect 115952 8294 115980 8463
rect 116044 8294 116072 9030
rect 116872 8809 116900 12406
rect 117228 12232 117280 12238
rect 117228 12174 117280 12180
rect 116950 11112 117006 11121
rect 117240 11082 117268 12174
rect 117318 11792 117374 11801
rect 117318 11727 117374 11736
rect 117332 11558 117360 11727
rect 117424 11558 117452 12406
rect 117320 11552 117372 11558
rect 117320 11494 117372 11500
rect 117412 11552 117464 11558
rect 117412 11494 117464 11500
rect 117424 11336 117452 11494
rect 117332 11308 117452 11336
rect 117332 11082 117360 11308
rect 117504 11280 117556 11286
rect 117424 11240 117504 11268
rect 117424 11150 117452 11240
rect 117504 11222 117556 11228
rect 117412 11144 117464 11150
rect 117412 11086 117464 11092
rect 117504 11144 117556 11150
rect 117504 11086 117556 11092
rect 116950 11047 117006 11056
rect 117228 11076 117280 11082
rect 116964 10742 116992 11047
rect 117228 11018 117280 11024
rect 117320 11076 117372 11082
rect 117320 11018 117372 11024
rect 116952 10736 117004 10742
rect 117332 10690 117360 11018
rect 116952 10678 117004 10684
rect 117240 10662 117360 10690
rect 117240 10062 117268 10662
rect 117320 10600 117372 10606
rect 117320 10542 117372 10548
rect 117228 10056 117280 10062
rect 117228 9998 117280 10004
rect 116950 9752 117006 9761
rect 117332 9722 117360 10542
rect 117412 9920 117464 9926
rect 117412 9862 117464 9868
rect 116950 9687 117006 9696
rect 117320 9716 117372 9722
rect 116964 8838 116992 9687
rect 117320 9658 117372 9664
rect 117136 9512 117188 9518
rect 117136 9454 117188 9460
rect 117148 8838 117176 9454
rect 117228 8900 117280 8906
rect 117228 8842 117280 8848
rect 116952 8832 117004 8838
rect 116858 8800 116914 8809
rect 116952 8774 117004 8780
rect 117136 8832 117188 8838
rect 117240 8809 117268 8842
rect 117136 8774 117188 8780
rect 117226 8800 117282 8809
rect 116858 8735 116914 8744
rect 116676 8424 116728 8430
rect 116676 8366 116728 8372
rect 116766 8392 116822 8401
rect 115940 8288 115992 8294
rect 115940 8230 115992 8236
rect 116032 8288 116084 8294
rect 116032 8230 116084 8236
rect 115848 6316 115900 6322
rect 115848 6258 115900 6264
rect 115860 6118 115888 6258
rect 115848 6112 115900 6118
rect 115848 6054 115900 6060
rect 116044 5370 116072 8230
rect 116214 7848 116270 7857
rect 116214 7783 116216 7792
rect 116268 7783 116270 7792
rect 116308 7812 116360 7818
rect 116216 7754 116268 7760
rect 116308 7754 116360 7760
rect 116320 6866 116348 7754
rect 116688 6934 116716 8366
rect 116766 8327 116822 8336
rect 116780 7546 116808 8327
rect 116768 7540 116820 7546
rect 116768 7482 116820 7488
rect 116676 6928 116728 6934
rect 116676 6870 116728 6876
rect 116872 6866 116900 8735
rect 116964 7410 116992 8774
rect 117148 8022 117176 8774
rect 117226 8735 117282 8744
rect 117320 8628 117372 8634
rect 117320 8570 117372 8576
rect 117332 8498 117360 8570
rect 117320 8492 117372 8498
rect 117320 8434 117372 8440
rect 117136 8016 117188 8022
rect 117136 7958 117188 7964
rect 117148 7886 117176 7958
rect 117424 7886 117452 9862
rect 117516 9382 117544 11086
rect 117700 10810 117728 12922
rect 117976 12714 118004 13330
rect 117964 12708 118016 12714
rect 117964 12650 118016 12656
rect 118068 12594 118096 14826
rect 118344 13530 118372 15200
rect 119068 14680 119120 14686
rect 119068 14622 119120 14628
rect 118332 13524 118384 13530
rect 118332 13466 118384 13472
rect 118792 12844 118844 12850
rect 118792 12786 118844 12792
rect 117976 12566 118096 12594
rect 118148 12640 118200 12646
rect 118148 12582 118200 12588
rect 117976 12306 118004 12566
rect 118160 12434 118188 12582
rect 118068 12406 118188 12434
rect 118516 12436 118568 12442
rect 117964 12300 118016 12306
rect 117964 12242 118016 12248
rect 117780 11144 117832 11150
rect 117780 11086 117832 11092
rect 117688 10804 117740 10810
rect 117688 10746 117740 10752
rect 117504 9376 117556 9382
rect 117504 9318 117556 9324
rect 117504 8628 117556 8634
rect 117504 8570 117556 8576
rect 117516 8430 117544 8570
rect 117504 8424 117556 8430
rect 117504 8366 117556 8372
rect 117596 8424 117648 8430
rect 117596 8366 117648 8372
rect 117504 8288 117556 8294
rect 117608 8242 117636 8366
rect 117556 8236 117636 8242
rect 117504 8230 117636 8236
rect 117516 8214 117636 8230
rect 117608 7954 117636 8214
rect 117792 7970 117820 11086
rect 117872 10668 117924 10674
rect 117872 10610 117924 10616
rect 117884 10470 117912 10610
rect 117872 10464 117924 10470
rect 117872 10406 117924 10412
rect 117964 9920 118016 9926
rect 117964 9862 118016 9868
rect 117976 9586 118004 9862
rect 117964 9580 118016 9586
rect 117964 9522 118016 9528
rect 118068 9466 118096 12406
rect 118568 12396 118648 12424
rect 118516 12378 118568 12384
rect 118516 12232 118568 12238
rect 118516 12174 118568 12180
rect 118240 11756 118292 11762
rect 118240 11698 118292 11704
rect 118148 11552 118200 11558
rect 118148 11494 118200 11500
rect 117596 7948 117648 7954
rect 117596 7890 117648 7896
rect 117700 7942 117820 7970
rect 117976 9438 118096 9466
rect 117136 7880 117188 7886
rect 117136 7822 117188 7828
rect 117412 7880 117464 7886
rect 117412 7822 117464 7828
rect 117044 7744 117096 7750
rect 117044 7686 117096 7692
rect 116952 7404 117004 7410
rect 116952 7346 117004 7352
rect 116308 6860 116360 6866
rect 116308 6802 116360 6808
rect 116860 6860 116912 6866
rect 116860 6802 116912 6808
rect 116124 6248 116176 6254
rect 116124 6190 116176 6196
rect 116032 5364 116084 5370
rect 116032 5306 116084 5312
rect 116044 5166 116072 5306
rect 116032 5160 116084 5166
rect 116032 5102 116084 5108
rect 115848 5092 115900 5098
rect 115848 5034 115900 5040
rect 115860 4486 115888 5034
rect 116136 4690 116164 6190
rect 116768 6180 116820 6186
rect 116768 6122 116820 6128
rect 116780 5914 116808 6122
rect 116768 5908 116820 5914
rect 116768 5850 116820 5856
rect 117056 5846 117084 7686
rect 117148 6458 117176 7822
rect 117412 7200 117464 7206
rect 117412 7142 117464 7148
rect 117424 7041 117452 7142
rect 117410 7032 117466 7041
rect 117410 6967 117466 6976
rect 117136 6452 117188 6458
rect 117136 6394 117188 6400
rect 117044 5840 117096 5846
rect 116950 5808 117006 5817
rect 117044 5782 117096 5788
rect 117148 5778 117176 6394
rect 117410 5944 117466 5953
rect 117410 5879 117412 5888
rect 117464 5879 117466 5888
rect 117412 5850 117464 5856
rect 116950 5743 117006 5752
rect 117136 5772 117188 5778
rect 116964 5302 116992 5743
rect 117136 5714 117188 5720
rect 117148 5302 117176 5714
rect 117424 5642 117452 5850
rect 117412 5636 117464 5642
rect 117412 5578 117464 5584
rect 116952 5296 117004 5302
rect 116952 5238 117004 5244
rect 117136 5296 117188 5302
rect 117136 5238 117188 5244
rect 117226 4856 117282 4865
rect 117226 4791 117228 4800
rect 117280 4791 117282 4800
rect 117228 4762 117280 4768
rect 116124 4684 116176 4690
rect 116124 4626 116176 4632
rect 116768 4684 116820 4690
rect 116768 4626 116820 4632
rect 115848 4480 115900 4486
rect 115848 4422 115900 4428
rect 115756 4140 115808 4146
rect 115756 4082 115808 4088
rect 116780 4078 116808 4626
rect 117700 4554 117728 7942
rect 117780 5160 117832 5166
rect 117780 5102 117832 5108
rect 117872 5160 117924 5166
rect 117872 5102 117924 5108
rect 117792 4826 117820 5102
rect 117780 4820 117832 4826
rect 117780 4762 117832 4768
rect 117792 4729 117820 4762
rect 117884 4758 117912 5102
rect 117872 4752 117924 4758
rect 117778 4720 117834 4729
rect 117872 4694 117924 4700
rect 117778 4655 117834 4664
rect 117688 4548 117740 4554
rect 117688 4490 117740 4496
rect 116768 4072 116820 4078
rect 116768 4014 116820 4020
rect 116780 3602 116808 4014
rect 117780 3936 117832 3942
rect 117780 3878 117832 3884
rect 116768 3596 116820 3602
rect 116768 3538 116820 3544
rect 117792 3534 117820 3878
rect 117976 3738 118004 9438
rect 118160 8974 118188 11494
rect 118252 10033 118280 11698
rect 118528 11694 118556 12174
rect 118516 11688 118568 11694
rect 118516 11630 118568 11636
rect 118528 11558 118556 11630
rect 118516 11552 118568 11558
rect 118516 11494 118568 11500
rect 118424 11348 118476 11354
rect 118424 11290 118476 11296
rect 118436 11218 118464 11290
rect 118620 11286 118648 12396
rect 118700 11892 118752 11898
rect 118700 11834 118752 11840
rect 118712 11694 118740 11834
rect 118700 11688 118752 11694
rect 118700 11630 118752 11636
rect 118608 11280 118660 11286
rect 118608 11222 118660 11228
rect 118424 11212 118476 11218
rect 118424 11154 118476 11160
rect 118514 10704 118570 10713
rect 118514 10639 118570 10648
rect 118608 10668 118660 10674
rect 118528 10266 118556 10639
rect 118608 10610 118660 10616
rect 118516 10260 118568 10266
rect 118516 10202 118568 10208
rect 118620 10062 118648 10610
rect 118804 10198 118832 12786
rect 118884 12096 118936 12102
rect 119080 12073 119108 14622
rect 119172 13462 119200 15286
rect 119434 15286 119752 15314
rect 119434 15200 119490 15286
rect 119160 13456 119212 13462
rect 119160 13398 119212 13404
rect 119160 13184 119212 13190
rect 119160 13126 119212 13132
rect 119172 12646 119200 13126
rect 119284 13084 119592 13093
rect 119284 13082 119290 13084
rect 119346 13082 119370 13084
rect 119426 13082 119450 13084
rect 119506 13082 119530 13084
rect 119586 13082 119592 13084
rect 119346 13030 119348 13082
rect 119528 13030 119530 13082
rect 119284 13028 119290 13030
rect 119346 13028 119370 13030
rect 119426 13028 119450 13030
rect 119506 13028 119530 13030
rect 119586 13028 119592 13030
rect 119284 13019 119592 13028
rect 119724 12986 119752 15286
rect 119986 15200 120042 16000
rect 120538 15200 120594 16000
rect 121090 15200 121146 16000
rect 121642 15200 121698 16000
rect 122194 15200 122250 16000
rect 122746 15200 122802 16000
rect 123298 15200 123354 16000
rect 123850 15200 123906 16000
rect 124402 15314 124458 16000
rect 124954 15314 125010 16000
rect 124402 15286 124720 15314
rect 124402 15200 124458 15286
rect 119896 13320 119948 13326
rect 119896 13262 119948 13268
rect 119712 12980 119764 12986
rect 119712 12922 119764 12928
rect 119252 12844 119304 12850
rect 119252 12786 119304 12792
rect 119264 12646 119292 12786
rect 119160 12640 119212 12646
rect 119160 12582 119212 12588
rect 119252 12640 119304 12646
rect 119252 12582 119304 12588
rect 118884 12038 118936 12044
rect 119066 12064 119122 12073
rect 118896 11937 118924 12038
rect 119066 11999 119122 12008
rect 118882 11928 118938 11937
rect 119080 11898 119108 11999
rect 118882 11863 118938 11872
rect 119068 11892 119120 11898
rect 119068 11834 119120 11840
rect 119172 11694 119200 12582
rect 119908 12434 119936 13262
rect 120000 13002 120028 15200
rect 120172 13728 120224 13734
rect 120172 13670 120224 13676
rect 120000 12986 120120 13002
rect 120000 12980 120132 12986
rect 120000 12974 120080 12980
rect 120080 12922 120132 12928
rect 120184 12850 120212 13670
rect 120552 13530 120580 15200
rect 120540 13524 120592 13530
rect 120540 13466 120592 13472
rect 120816 13320 120868 13326
rect 120816 13262 120868 13268
rect 120908 13320 120960 13326
rect 120908 13262 120960 13268
rect 120632 12912 120684 12918
rect 120828 12889 120856 13262
rect 120920 13025 120948 13262
rect 120906 13016 120962 13025
rect 121104 12986 121132 15200
rect 121366 14104 121422 14113
rect 121366 14039 121422 14048
rect 121380 13394 121408 14039
rect 121368 13388 121420 13394
rect 121368 13330 121420 13336
rect 121458 13288 121514 13297
rect 121458 13223 121514 13232
rect 120906 12951 120962 12960
rect 121092 12980 121144 12986
rect 121092 12922 121144 12928
rect 120632 12854 120684 12860
rect 120814 12880 120870 12889
rect 120172 12844 120224 12850
rect 120172 12786 120224 12792
rect 120172 12708 120224 12714
rect 120172 12650 120224 12656
rect 119816 12406 119936 12434
rect 119284 11996 119592 12005
rect 119284 11994 119290 11996
rect 119346 11994 119370 11996
rect 119426 11994 119450 11996
rect 119506 11994 119530 11996
rect 119586 11994 119592 11996
rect 119346 11942 119348 11994
rect 119528 11942 119530 11994
rect 119284 11940 119290 11942
rect 119346 11940 119370 11942
rect 119426 11940 119450 11942
rect 119506 11940 119530 11942
rect 119586 11940 119592 11942
rect 119284 11931 119592 11940
rect 119436 11892 119488 11898
rect 119436 11834 119488 11840
rect 119160 11688 119212 11694
rect 119160 11630 119212 11636
rect 118884 11620 118936 11626
rect 118884 11562 118936 11568
rect 118792 10192 118844 10198
rect 118792 10134 118844 10140
rect 118608 10056 118660 10062
rect 118238 10024 118294 10033
rect 118608 9998 118660 10004
rect 118238 9959 118294 9968
rect 118332 9988 118384 9994
rect 118332 9930 118384 9936
rect 118344 9382 118372 9930
rect 118332 9376 118384 9382
rect 118332 9318 118384 9324
rect 118344 9178 118372 9318
rect 118332 9172 118384 9178
rect 118332 9114 118384 9120
rect 118148 8968 118200 8974
rect 118148 8910 118200 8916
rect 118424 8900 118476 8906
rect 118424 8842 118476 8848
rect 118332 8424 118384 8430
rect 118436 8401 118464 8842
rect 118516 8424 118568 8430
rect 118332 8366 118384 8372
rect 118422 8392 118478 8401
rect 118148 6656 118200 6662
rect 118148 6598 118200 6604
rect 118056 5228 118108 5234
rect 118056 5170 118108 5176
rect 118068 4554 118096 5170
rect 118160 5098 118188 6598
rect 118240 6112 118292 6118
rect 118240 6054 118292 6060
rect 118148 5092 118200 5098
rect 118148 5034 118200 5040
rect 118148 4752 118200 4758
rect 118148 4694 118200 4700
rect 118056 4548 118108 4554
rect 118056 4490 118108 4496
rect 118160 4486 118188 4694
rect 118148 4480 118200 4486
rect 118148 4422 118200 4428
rect 118252 4146 118280 6054
rect 118344 5234 118372 8366
rect 118516 8366 118568 8372
rect 118422 8327 118478 8336
rect 118424 7472 118476 7478
rect 118424 7414 118476 7420
rect 118436 5370 118464 7414
rect 118424 5364 118476 5370
rect 118424 5306 118476 5312
rect 118332 5228 118384 5234
rect 118332 5170 118384 5176
rect 118436 4146 118464 5306
rect 118240 4140 118292 4146
rect 118240 4082 118292 4088
rect 118424 4140 118476 4146
rect 118424 4082 118476 4088
rect 118252 3777 118280 4082
rect 118528 4026 118556 8366
rect 118608 7948 118660 7954
rect 118608 7890 118660 7896
rect 118620 6866 118648 7890
rect 118700 7880 118752 7886
rect 118700 7822 118752 7828
rect 118608 6860 118660 6866
rect 118608 6802 118660 6808
rect 118712 6798 118740 7822
rect 118700 6792 118752 6798
rect 118700 6734 118752 6740
rect 118608 5704 118660 5710
rect 118608 5646 118660 5652
rect 118620 4146 118648 5646
rect 118896 5370 118924 11562
rect 119448 11354 119476 11834
rect 119620 11552 119672 11558
rect 119620 11494 119672 11500
rect 119632 11354 119660 11494
rect 119436 11348 119488 11354
rect 119436 11290 119488 11296
rect 119620 11348 119672 11354
rect 119620 11290 119672 11296
rect 119160 11076 119212 11082
rect 119160 11018 119212 11024
rect 119620 11076 119672 11082
rect 119620 11018 119672 11024
rect 118974 10840 119030 10849
rect 118974 10775 119030 10784
rect 118988 10198 119016 10775
rect 119172 10606 119200 11018
rect 119284 10908 119592 10917
rect 119284 10906 119290 10908
rect 119346 10906 119370 10908
rect 119426 10906 119450 10908
rect 119506 10906 119530 10908
rect 119586 10906 119592 10908
rect 119346 10854 119348 10906
rect 119528 10854 119530 10906
rect 119284 10852 119290 10854
rect 119346 10852 119370 10854
rect 119426 10852 119450 10854
rect 119506 10852 119530 10854
rect 119586 10852 119592 10854
rect 119284 10843 119592 10852
rect 119160 10600 119212 10606
rect 119160 10542 119212 10548
rect 118976 10192 119028 10198
rect 119172 10146 119200 10542
rect 118976 10134 119028 10140
rect 119080 10118 119200 10146
rect 118976 8832 119028 8838
rect 118976 8774 119028 8780
rect 118988 8537 119016 8774
rect 118974 8528 119030 8537
rect 118974 8463 118976 8472
rect 119028 8463 119030 8472
rect 118976 8434 119028 8440
rect 119080 8344 119108 10118
rect 119160 10056 119212 10062
rect 119160 9998 119212 10004
rect 119172 9761 119200 9998
rect 119284 9820 119592 9829
rect 119284 9818 119290 9820
rect 119346 9818 119370 9820
rect 119426 9818 119450 9820
rect 119506 9818 119530 9820
rect 119586 9818 119592 9820
rect 119346 9766 119348 9818
rect 119528 9766 119530 9818
rect 119284 9764 119290 9766
rect 119346 9764 119370 9766
rect 119426 9764 119450 9766
rect 119506 9764 119530 9766
rect 119586 9764 119592 9766
rect 119158 9752 119214 9761
rect 119284 9755 119592 9764
rect 119158 9687 119214 9696
rect 119632 8974 119660 11018
rect 119816 9382 119844 12406
rect 119896 12096 119948 12102
rect 119896 12038 119948 12044
rect 119804 9376 119856 9382
rect 119804 9318 119856 9324
rect 119620 8968 119672 8974
rect 119620 8910 119672 8916
rect 119160 8832 119212 8838
rect 119158 8800 119160 8809
rect 119212 8800 119214 8809
rect 119158 8735 119214 8744
rect 119284 8732 119592 8741
rect 119284 8730 119290 8732
rect 119346 8730 119370 8732
rect 119426 8730 119450 8732
rect 119506 8730 119530 8732
rect 119586 8730 119592 8732
rect 119346 8678 119348 8730
rect 119528 8678 119530 8730
rect 119284 8676 119290 8678
rect 119346 8676 119370 8678
rect 119426 8676 119450 8678
rect 119506 8676 119530 8678
rect 119586 8676 119592 8678
rect 119284 8667 119592 8676
rect 119160 8424 119212 8430
rect 119160 8366 119212 8372
rect 118988 8316 119108 8344
rect 118988 7206 119016 8316
rect 119068 7404 119120 7410
rect 119068 7346 119120 7352
rect 118976 7200 119028 7206
rect 118976 7142 119028 7148
rect 118988 5710 119016 7142
rect 119080 6390 119108 7346
rect 119068 6384 119120 6390
rect 119068 6326 119120 6332
rect 118976 5704 119028 5710
rect 118976 5646 119028 5652
rect 118700 5364 118752 5370
rect 118700 5306 118752 5312
rect 118884 5364 118936 5370
rect 118884 5306 118936 5312
rect 118712 4865 118740 5306
rect 118698 4856 118754 4865
rect 118698 4791 118754 4800
rect 118792 4276 118844 4282
rect 118792 4218 118844 4224
rect 118608 4140 118660 4146
rect 118608 4082 118660 4088
rect 118436 3998 118556 4026
rect 118238 3768 118294 3777
rect 117964 3732 118016 3738
rect 118238 3703 118294 3712
rect 117964 3674 118016 3680
rect 117780 3528 117832 3534
rect 117780 3470 117832 3476
rect 116952 3460 117004 3466
rect 116952 3402 117004 3408
rect 117688 3460 117740 3466
rect 117688 3402 117740 3408
rect 116964 3194 116992 3402
rect 115664 3188 115716 3194
rect 115664 3130 115716 3136
rect 116952 3188 117004 3194
rect 116952 3130 117004 3136
rect 117700 2854 117728 3402
rect 118252 3398 118280 3703
rect 118240 3392 118292 3398
rect 118240 3334 118292 3340
rect 118436 3058 118464 3998
rect 118804 3641 118832 4218
rect 118988 4010 119016 5646
rect 119068 5092 119120 5098
rect 119068 5034 119120 5040
rect 119080 4826 119108 5034
rect 119172 5012 119200 8366
rect 119436 8356 119488 8362
rect 119436 8298 119488 8304
rect 119448 8022 119476 8298
rect 119436 8016 119488 8022
rect 119436 7958 119488 7964
rect 119284 7644 119592 7653
rect 119284 7642 119290 7644
rect 119346 7642 119370 7644
rect 119426 7642 119450 7644
rect 119506 7642 119530 7644
rect 119586 7642 119592 7644
rect 119346 7590 119348 7642
rect 119528 7590 119530 7642
rect 119284 7588 119290 7590
rect 119346 7588 119370 7590
rect 119426 7588 119450 7590
rect 119506 7588 119530 7590
rect 119586 7588 119592 7590
rect 119284 7579 119592 7588
rect 119284 6556 119592 6565
rect 119284 6554 119290 6556
rect 119346 6554 119370 6556
rect 119426 6554 119450 6556
rect 119506 6554 119530 6556
rect 119586 6554 119592 6556
rect 119346 6502 119348 6554
rect 119528 6502 119530 6554
rect 119284 6500 119290 6502
rect 119346 6500 119370 6502
rect 119426 6500 119450 6502
rect 119506 6500 119530 6502
rect 119586 6500 119592 6502
rect 119284 6491 119592 6500
rect 119712 6112 119764 6118
rect 119712 6054 119764 6060
rect 119284 5468 119592 5477
rect 119284 5466 119290 5468
rect 119346 5466 119370 5468
rect 119426 5466 119450 5468
rect 119506 5466 119530 5468
rect 119586 5466 119592 5468
rect 119346 5414 119348 5466
rect 119528 5414 119530 5466
rect 119284 5412 119290 5414
rect 119346 5412 119370 5414
rect 119426 5412 119450 5414
rect 119506 5412 119530 5414
rect 119586 5412 119592 5414
rect 119284 5403 119592 5412
rect 119252 5024 119304 5030
rect 119172 4984 119252 5012
rect 119252 4966 119304 4972
rect 119068 4820 119120 4826
rect 119068 4762 119120 4768
rect 119264 4690 119292 4966
rect 119252 4684 119304 4690
rect 119252 4626 119304 4632
rect 119172 4542 119292 4570
rect 119172 4214 119200 4542
rect 119264 4486 119292 4542
rect 119252 4480 119304 4486
rect 119252 4422 119304 4428
rect 119284 4380 119592 4389
rect 119284 4378 119290 4380
rect 119346 4378 119370 4380
rect 119426 4378 119450 4380
rect 119506 4378 119530 4380
rect 119586 4378 119592 4380
rect 119346 4326 119348 4378
rect 119528 4326 119530 4378
rect 119284 4324 119290 4326
rect 119346 4324 119370 4326
rect 119426 4324 119450 4326
rect 119506 4324 119530 4326
rect 119586 4324 119592 4326
rect 119284 4315 119592 4324
rect 119160 4208 119212 4214
rect 119160 4150 119212 4156
rect 118976 4004 119028 4010
rect 118976 3946 119028 3952
rect 119252 3936 119304 3942
rect 119252 3878 119304 3884
rect 119264 3777 119292 3878
rect 119250 3768 119306 3777
rect 119250 3703 119306 3712
rect 118790 3632 118846 3641
rect 118790 3567 118846 3576
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 118516 3120 118568 3126
rect 118516 3062 118568 3068
rect 118424 3052 118476 3058
rect 118424 2994 118476 3000
rect 117596 2848 117648 2854
rect 117594 2816 117596 2825
rect 117688 2848 117740 2854
rect 117648 2816 117650 2825
rect 117688 2790 117740 2796
rect 117594 2751 117650 2760
rect 118528 2689 118556 3062
rect 118514 2680 118570 2689
rect 118514 2615 118570 2624
rect 118804 2446 118832 3470
rect 119724 3398 119752 6054
rect 119712 3392 119764 3398
rect 119712 3334 119764 3340
rect 119284 3292 119592 3301
rect 119284 3290 119290 3292
rect 119346 3290 119370 3292
rect 119426 3290 119450 3292
rect 119506 3290 119530 3292
rect 119586 3290 119592 3292
rect 119346 3238 119348 3290
rect 119528 3238 119530 3290
rect 119284 3236 119290 3238
rect 119346 3236 119370 3238
rect 119426 3236 119450 3238
rect 119506 3236 119530 3238
rect 119586 3236 119592 3238
rect 119284 3227 119592 3236
rect 119160 3188 119212 3194
rect 119160 3130 119212 3136
rect 119172 2854 119200 3130
rect 119160 2848 119212 2854
rect 119160 2790 119212 2796
rect 119344 2848 119396 2854
rect 119344 2790 119396 2796
rect 118792 2440 118844 2446
rect 117410 2408 117466 2417
rect 118792 2382 118844 2388
rect 119356 2378 119384 2790
rect 117410 2343 117466 2352
rect 119344 2372 119396 2378
rect 117424 2310 117452 2343
rect 119344 2314 119396 2320
rect 117412 2304 117464 2310
rect 117412 2246 117464 2252
rect 119284 2204 119592 2213
rect 119284 2202 119290 2204
rect 119346 2202 119370 2204
rect 119426 2202 119450 2204
rect 119506 2202 119530 2204
rect 119586 2202 119592 2204
rect 119346 2150 119348 2202
rect 119528 2150 119530 2202
rect 119284 2148 119290 2150
rect 119346 2148 119370 2150
rect 119426 2148 119450 2150
rect 119506 2148 119530 2150
rect 119586 2148 119592 2150
rect 119284 2139 119592 2148
rect 115572 1692 115624 1698
rect 115572 1634 115624 1640
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 119816 1154 119844 9318
rect 119908 8242 119936 12038
rect 120184 11937 120212 12650
rect 120262 12472 120318 12481
rect 120262 12407 120318 12416
rect 120644 12434 120672 12854
rect 121472 12850 121500 13223
rect 120814 12815 120870 12824
rect 121460 12844 121512 12850
rect 121460 12786 121512 12792
rect 121656 12442 121684 15200
rect 122104 13796 122156 13802
rect 122104 13738 122156 13744
rect 122012 13388 122064 13394
rect 122012 13330 122064 13336
rect 122024 12782 122052 13330
rect 122116 13326 122144 13738
rect 122208 13410 122236 15200
rect 122760 13530 122788 15200
rect 123024 13864 123076 13870
rect 123024 13806 123076 13812
rect 122748 13524 122800 13530
rect 122748 13466 122800 13472
rect 122208 13382 122512 13410
rect 122104 13320 122156 13326
rect 122104 13262 122156 13268
rect 122378 13152 122434 13161
rect 122378 13087 122434 13096
rect 122012 12776 122064 12782
rect 122012 12718 122064 12724
rect 121644 12436 121696 12442
rect 120170 11928 120226 11937
rect 120170 11863 120226 11872
rect 120184 11150 120212 11863
rect 120172 11144 120224 11150
rect 120172 11086 120224 11092
rect 120172 10736 120224 10742
rect 120172 10678 120224 10684
rect 120184 10470 120212 10678
rect 120172 10464 120224 10470
rect 120172 10406 120224 10412
rect 119988 9920 120040 9926
rect 119988 9862 120040 9868
rect 120000 9382 120028 9862
rect 119988 9376 120040 9382
rect 119988 9318 120040 9324
rect 120000 8430 120028 9318
rect 120276 8922 120304 12407
rect 120644 12406 120856 12434
rect 120448 12232 120500 12238
rect 120448 12174 120500 12180
rect 120460 11558 120488 12174
rect 120828 12102 120856 12406
rect 121644 12378 121696 12384
rect 121828 12436 121880 12442
rect 121828 12378 121880 12384
rect 121840 12238 121868 12378
rect 121828 12232 121880 12238
rect 121828 12174 121880 12180
rect 120816 12096 120868 12102
rect 120814 12064 120816 12073
rect 120868 12064 120870 12073
rect 120814 11999 120870 12008
rect 121642 11792 121698 11801
rect 121184 11756 121236 11762
rect 121642 11727 121698 11736
rect 121184 11698 121236 11704
rect 120448 11552 120500 11558
rect 120448 11494 120500 11500
rect 120540 11552 120592 11558
rect 120540 11494 120592 11500
rect 120552 10674 120580 11494
rect 121000 11348 121052 11354
rect 121000 11290 121052 11296
rect 121012 11150 121040 11290
rect 121196 11257 121224 11698
rect 121368 11688 121420 11694
rect 121368 11630 121420 11636
rect 121380 11393 121408 11630
rect 121366 11384 121422 11393
rect 121366 11319 121422 11328
rect 121182 11248 121238 11257
rect 121182 11183 121238 11192
rect 121000 11144 121052 11150
rect 121000 11086 121052 11092
rect 121012 10690 121040 11086
rect 120540 10668 120592 10674
rect 121012 10662 121132 10690
rect 120540 10610 120592 10616
rect 120356 10464 120408 10470
rect 120354 10432 120356 10441
rect 121000 10464 121052 10470
rect 120408 10432 120410 10441
rect 121000 10406 121052 10412
rect 120354 10367 120410 10376
rect 120724 10124 120776 10130
rect 120724 10066 120776 10072
rect 120736 10033 120764 10066
rect 120722 10024 120778 10033
rect 120448 9988 120500 9994
rect 120722 9959 120778 9968
rect 120448 9930 120500 9936
rect 120276 8894 120396 8922
rect 120460 8906 120488 9930
rect 121012 9722 121040 10406
rect 121104 10062 121132 10662
rect 121092 10056 121144 10062
rect 121092 9998 121144 10004
rect 121000 9716 121052 9722
rect 121000 9658 121052 9664
rect 121104 9586 121132 9998
rect 121092 9580 121144 9586
rect 121092 9522 121144 9528
rect 121380 9382 121408 11319
rect 121552 9920 121604 9926
rect 121552 9862 121604 9868
rect 121368 9376 121420 9382
rect 121368 9318 121420 9324
rect 120724 9104 120776 9110
rect 120724 9046 120776 9052
rect 120264 8832 120316 8838
rect 120264 8774 120316 8780
rect 120170 8528 120226 8537
rect 120170 8463 120226 8472
rect 119988 8424 120040 8430
rect 119988 8366 120040 8372
rect 120184 8294 120212 8463
rect 120172 8288 120224 8294
rect 119908 8214 120120 8242
rect 120172 8230 120224 8236
rect 119988 7200 120040 7206
rect 119988 7142 120040 7148
rect 120000 7002 120028 7142
rect 119988 6996 120040 7002
rect 119988 6938 120040 6944
rect 119896 6248 119948 6254
rect 119896 6190 119948 6196
rect 119908 3534 119936 6190
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 120000 2553 120028 6938
rect 120092 6497 120120 8214
rect 120172 6656 120224 6662
rect 120172 6598 120224 6604
rect 120078 6488 120134 6497
rect 120078 6423 120134 6432
rect 120184 5302 120212 6598
rect 120172 5296 120224 5302
rect 120172 5238 120224 5244
rect 120080 3936 120132 3942
rect 120080 3878 120132 3884
rect 120092 2990 120120 3878
rect 120080 2984 120132 2990
rect 120080 2926 120132 2932
rect 120170 2816 120226 2825
rect 120276 2774 120304 8774
rect 120368 4486 120396 8894
rect 120448 8900 120500 8906
rect 120448 8842 120500 8848
rect 120736 8673 120764 9046
rect 120908 8968 120960 8974
rect 120908 8910 120960 8916
rect 120722 8664 120778 8673
rect 120722 8599 120778 8608
rect 120632 6996 120684 7002
rect 120632 6938 120684 6944
rect 120540 6452 120592 6458
rect 120540 6394 120592 6400
rect 120552 5914 120580 6394
rect 120540 5908 120592 5914
rect 120540 5850 120592 5856
rect 120356 4480 120408 4486
rect 120354 4448 120356 4457
rect 120408 4448 120410 4457
rect 120354 4383 120410 4392
rect 120644 2990 120672 6938
rect 120816 6792 120868 6798
rect 120816 6734 120868 6740
rect 120828 5914 120856 6734
rect 120816 5908 120868 5914
rect 120816 5850 120868 5856
rect 120920 2990 120948 8910
rect 121368 8832 121420 8838
rect 121420 8792 121500 8820
rect 121368 8774 121420 8780
rect 121472 8294 121500 8792
rect 121460 8288 121512 8294
rect 121460 8230 121512 8236
rect 121366 8120 121422 8129
rect 121276 8084 121328 8090
rect 121366 8055 121422 8064
rect 121276 8026 121328 8032
rect 121092 6656 121144 6662
rect 121092 6598 121144 6604
rect 121000 4004 121052 4010
rect 121000 3946 121052 3952
rect 121012 3602 121040 3946
rect 121000 3596 121052 3602
rect 121000 3538 121052 3544
rect 121104 3126 121132 6598
rect 121184 5704 121236 5710
rect 121184 5646 121236 5652
rect 121196 4486 121224 5646
rect 121184 4480 121236 4486
rect 121184 4422 121236 4428
rect 121196 3942 121224 4422
rect 121184 3936 121236 3942
rect 121184 3878 121236 3884
rect 121288 3466 121316 8026
rect 121380 5574 121408 8055
rect 121472 7818 121500 8230
rect 121460 7812 121512 7818
rect 121460 7754 121512 7760
rect 121564 6662 121592 9862
rect 121656 7936 121684 11727
rect 122024 11694 122052 12718
rect 122392 12646 122420 13087
rect 122484 12646 122512 13382
rect 122380 12640 122432 12646
rect 122380 12582 122432 12588
rect 122472 12640 122524 12646
rect 122472 12582 122524 12588
rect 122748 12300 122800 12306
rect 122748 12242 122800 12248
rect 122012 11688 122064 11694
rect 122012 11630 122064 11636
rect 121920 11552 121972 11558
rect 121920 11494 121972 11500
rect 121932 11150 121960 11494
rect 121920 11144 121972 11150
rect 121920 11086 121972 11092
rect 121828 11008 121880 11014
rect 122024 10996 122052 11630
rect 122760 11558 122788 12242
rect 122838 12200 122894 12209
rect 122838 12135 122894 12144
rect 122748 11552 122800 11558
rect 122748 11494 122800 11500
rect 122564 11144 122616 11150
rect 122564 11086 122616 11092
rect 122656 11144 122708 11150
rect 122656 11086 122708 11092
rect 122104 11076 122156 11082
rect 122104 11018 122156 11024
rect 121880 10968 122052 10996
rect 121828 10950 121880 10956
rect 121734 10432 121790 10441
rect 121734 10367 121790 10376
rect 121748 9518 121776 10367
rect 121932 10130 121960 10968
rect 122116 10674 122144 11018
rect 122104 10668 122156 10674
rect 122104 10610 122156 10616
rect 122288 10668 122340 10674
rect 122576 10656 122604 11086
rect 122668 10810 122696 11086
rect 122656 10804 122708 10810
rect 122656 10746 122708 10752
rect 122576 10628 122696 10656
rect 122288 10610 122340 10616
rect 122300 10198 122328 10610
rect 122380 10600 122432 10606
rect 122380 10542 122432 10548
rect 122288 10192 122340 10198
rect 122288 10134 122340 10140
rect 122392 10130 122420 10542
rect 122564 10532 122616 10538
rect 122564 10474 122616 10480
rect 122576 10266 122604 10474
rect 122564 10260 122616 10266
rect 122564 10202 122616 10208
rect 121920 10124 121972 10130
rect 121920 10066 121972 10072
rect 122380 10124 122432 10130
rect 122380 10066 122432 10072
rect 121932 9586 121960 10066
rect 122564 10056 122616 10062
rect 122564 9998 122616 10004
rect 122668 10010 122696 10628
rect 122760 10130 122788 11494
rect 122852 10470 122880 12135
rect 123036 11218 123064 13806
rect 123312 12986 123340 15200
rect 123484 13252 123536 13258
rect 123484 13194 123536 13200
rect 123208 12980 123260 12986
rect 123208 12922 123260 12928
rect 123300 12980 123352 12986
rect 123300 12922 123352 12928
rect 123220 11558 123248 12922
rect 123392 12912 123444 12918
rect 123392 12854 123444 12860
rect 123298 12472 123354 12481
rect 123298 12407 123354 12416
rect 123208 11552 123260 11558
rect 123208 11494 123260 11500
rect 123024 11212 123076 11218
rect 123024 11154 123076 11160
rect 122932 11008 122984 11014
rect 122932 10950 122984 10956
rect 122944 10810 122972 10950
rect 122932 10804 122984 10810
rect 122932 10746 122984 10752
rect 123220 10713 123248 11494
rect 123206 10704 123262 10713
rect 123206 10639 123262 10648
rect 122840 10464 122892 10470
rect 122840 10406 122892 10412
rect 122932 10260 122984 10266
rect 122932 10202 122984 10208
rect 122748 10124 122800 10130
rect 122748 10066 122800 10072
rect 122840 10056 122892 10062
rect 122668 10004 122840 10010
rect 122944 10033 122972 10202
rect 122668 9998 122892 10004
rect 122930 10024 122986 10033
rect 121920 9580 121972 9586
rect 121920 9522 121972 9528
rect 121736 9512 121788 9518
rect 121736 9454 121788 9460
rect 121932 9466 121960 9522
rect 121932 9438 122052 9466
rect 121920 9104 121972 9110
rect 121826 9072 121882 9081
rect 121920 9046 121972 9052
rect 121826 9007 121882 9016
rect 121840 8974 121868 9007
rect 121828 8968 121880 8974
rect 121828 8910 121880 8916
rect 121932 8634 121960 9046
rect 121920 8628 121972 8634
rect 121920 8570 121972 8576
rect 122024 8362 122052 9438
rect 122380 8832 122432 8838
rect 122378 8800 122380 8809
rect 122472 8832 122524 8838
rect 122432 8800 122434 8809
rect 122472 8774 122524 8780
rect 122378 8735 122434 8744
rect 122012 8356 122064 8362
rect 122012 8298 122064 8304
rect 121828 8016 121880 8022
rect 121828 7958 121880 7964
rect 121656 7908 121776 7936
rect 121644 7812 121696 7818
rect 121644 7754 121696 7760
rect 121656 7342 121684 7754
rect 121644 7336 121696 7342
rect 121644 7278 121696 7284
rect 121656 6866 121684 7278
rect 121748 7274 121776 7908
rect 121736 7268 121788 7274
rect 121736 7210 121788 7216
rect 121840 7177 121868 7958
rect 122484 7818 122512 8774
rect 122472 7812 122524 7818
rect 122472 7754 122524 7760
rect 122012 7200 122064 7206
rect 121826 7168 121882 7177
rect 122012 7142 122064 7148
rect 122472 7200 122524 7206
rect 122472 7142 122524 7148
rect 121826 7103 121882 7112
rect 122024 6934 122052 7142
rect 122012 6928 122064 6934
rect 122012 6870 122064 6876
rect 121644 6860 121696 6866
rect 121644 6802 121696 6808
rect 121552 6656 121604 6662
rect 121552 6598 121604 6604
rect 121644 6656 121696 6662
rect 121644 6598 121696 6604
rect 121656 6458 121684 6598
rect 121644 6452 121696 6458
rect 121644 6394 121696 6400
rect 121920 6452 121972 6458
rect 121920 6394 121972 6400
rect 121828 6384 121880 6390
rect 121828 6326 121880 6332
rect 121840 6254 121868 6326
rect 121828 6248 121880 6254
rect 121828 6190 121880 6196
rect 121736 5840 121788 5846
rect 121736 5782 121788 5788
rect 121748 5710 121776 5782
rect 121736 5704 121788 5710
rect 121736 5646 121788 5652
rect 121368 5568 121420 5574
rect 121840 5556 121868 6190
rect 121932 5914 121960 6394
rect 122484 5914 122512 7142
rect 122576 6866 122604 9998
rect 122668 9982 122880 9998
rect 122564 6860 122616 6866
rect 122564 6802 122616 6808
rect 122656 6792 122708 6798
rect 122656 6734 122708 6740
rect 122564 6316 122616 6322
rect 122564 6258 122616 6264
rect 122576 5914 122604 6258
rect 121920 5908 121972 5914
rect 121920 5850 121972 5856
rect 122472 5908 122524 5914
rect 122472 5850 122524 5856
rect 122564 5908 122616 5914
rect 122564 5850 122616 5856
rect 121368 5510 121420 5516
rect 121748 5528 121868 5556
rect 121748 5166 121776 5528
rect 121828 5296 121880 5302
rect 121828 5238 121880 5244
rect 121736 5160 121788 5166
rect 121736 5102 121788 5108
rect 121840 4826 121868 5238
rect 122484 4826 122512 5850
rect 122564 5568 122616 5574
rect 122564 5510 122616 5516
rect 121828 4820 121880 4826
rect 121828 4762 121880 4768
rect 122472 4820 122524 4826
rect 122472 4762 122524 4768
rect 122012 3936 122064 3942
rect 122012 3878 122064 3884
rect 121276 3460 121328 3466
rect 121276 3402 121328 3408
rect 122024 3126 122052 3878
rect 122576 3398 122604 5510
rect 122668 5370 122696 6734
rect 122760 6390 122788 9982
rect 122930 9959 122986 9968
rect 123312 9450 123340 12407
rect 123404 10198 123432 12854
rect 123496 12434 123524 13194
rect 123864 12434 123892 15200
rect 124312 14272 124364 14278
rect 124312 14214 124364 14220
rect 124324 13190 124352 14214
rect 124692 13462 124720 15286
rect 124954 15286 125272 15314
rect 124954 15200 125010 15286
rect 124680 13456 124732 13462
rect 124680 13398 124732 13404
rect 124772 13388 124824 13394
rect 124772 13330 124824 13336
rect 124784 13297 124812 13330
rect 124770 13288 124826 13297
rect 124770 13223 124826 13232
rect 124312 13184 124364 13190
rect 124404 13184 124456 13190
rect 124312 13126 124364 13132
rect 124402 13152 124404 13161
rect 124456 13152 124458 13161
rect 124402 13087 124458 13096
rect 124862 12880 124918 12889
rect 124312 12844 124364 12850
rect 124862 12815 124918 12824
rect 124312 12786 124364 12792
rect 124324 12434 124352 12786
rect 123496 12406 123616 12434
rect 123864 12406 124076 12434
rect 124324 12406 124444 12434
rect 123392 10192 123444 10198
rect 123392 10134 123444 10140
rect 123588 9994 123616 12406
rect 124048 12322 124076 12406
rect 124048 12294 124352 12322
rect 123852 12232 123904 12238
rect 123850 12200 123852 12209
rect 123904 12200 123906 12209
rect 123760 12164 123812 12170
rect 123850 12135 123906 12144
rect 123760 12106 123812 12112
rect 123668 11552 123720 11558
rect 123668 11494 123720 11500
rect 123680 11257 123708 11494
rect 123666 11248 123722 11257
rect 123666 11183 123722 11192
rect 123668 11008 123720 11014
rect 123668 10950 123720 10956
rect 123680 10470 123708 10950
rect 123772 10674 123800 12106
rect 123864 11694 123892 12135
rect 124324 12102 124352 12294
rect 124312 12096 124364 12102
rect 124312 12038 124364 12044
rect 124310 11792 124366 11801
rect 124310 11727 124366 11736
rect 123852 11688 123904 11694
rect 123852 11630 123904 11636
rect 124220 11552 124272 11558
rect 123942 11520 123998 11529
rect 124324 11540 124352 11727
rect 124272 11512 124352 11540
rect 124220 11494 124272 11500
rect 123942 11455 123998 11464
rect 123760 10668 123812 10674
rect 123760 10610 123812 10616
rect 123668 10464 123720 10470
rect 123668 10406 123720 10412
rect 123760 10464 123812 10470
rect 123760 10406 123812 10412
rect 123576 9988 123628 9994
rect 123576 9930 123628 9936
rect 123300 9444 123352 9450
rect 123300 9386 123352 9392
rect 123588 8922 123616 9930
rect 123496 8894 123616 8922
rect 122930 8528 122986 8537
rect 122840 8492 122892 8498
rect 122930 8463 122986 8472
rect 123300 8492 123352 8498
rect 122840 8434 122892 8440
rect 122852 7750 122880 8434
rect 122840 7744 122892 7750
rect 122840 7686 122892 7692
rect 122838 7032 122894 7041
rect 122838 6967 122894 6976
rect 122748 6384 122800 6390
rect 122748 6326 122800 6332
rect 122746 6080 122802 6089
rect 122852 6066 122880 6967
rect 122802 6038 122880 6066
rect 122746 6015 122802 6024
rect 122656 5364 122708 5370
rect 122656 5306 122708 5312
rect 122840 5092 122892 5098
rect 122840 5034 122892 5040
rect 122746 4720 122802 4729
rect 122746 4655 122748 4664
rect 122800 4655 122802 4664
rect 122748 4626 122800 4632
rect 122852 4622 122880 5034
rect 122840 4616 122892 4622
rect 122840 4558 122892 4564
rect 122944 4298 122972 8463
rect 123300 8434 123352 8440
rect 123024 8424 123076 8430
rect 123024 8366 123076 8372
rect 123036 8022 123064 8366
rect 123312 8294 123340 8434
rect 123300 8288 123352 8294
rect 123300 8230 123352 8236
rect 123024 8016 123076 8022
rect 123024 7958 123076 7964
rect 123300 8016 123352 8022
rect 123300 7958 123352 7964
rect 123208 7744 123260 7750
rect 123208 7686 123260 7692
rect 123116 7472 123168 7478
rect 123116 7414 123168 7420
rect 123128 6934 123156 7414
rect 123116 6928 123168 6934
rect 123116 6870 123168 6876
rect 123024 6792 123076 6798
rect 123024 6734 123076 6740
rect 123036 6202 123064 6734
rect 123036 6186 123156 6202
rect 123036 6180 123168 6186
rect 123036 6174 123116 6180
rect 123036 5778 123064 6174
rect 123116 6122 123168 6128
rect 123024 5772 123076 5778
rect 123024 5714 123076 5720
rect 123024 5636 123076 5642
rect 123024 5578 123076 5584
rect 122760 4270 122972 4298
rect 122760 4146 122788 4270
rect 122748 4140 122800 4146
rect 122748 4082 122800 4088
rect 122840 4140 122892 4146
rect 122840 4082 122892 4088
rect 122852 4026 122880 4082
rect 122760 4010 122880 4026
rect 122748 4004 122880 4010
rect 122800 3998 122880 4004
rect 122748 3946 122800 3952
rect 122944 3602 122972 4270
rect 123036 3670 123064 5578
rect 123114 5536 123170 5545
rect 123114 5471 123170 5480
rect 123128 5370 123156 5471
rect 123116 5364 123168 5370
rect 123116 5306 123168 5312
rect 123024 3664 123076 3670
rect 123024 3606 123076 3612
rect 122932 3596 122984 3602
rect 122932 3538 122984 3544
rect 122564 3392 122616 3398
rect 122564 3334 122616 3340
rect 123024 3392 123076 3398
rect 123024 3334 123076 3340
rect 121092 3120 121144 3126
rect 121092 3062 121144 3068
rect 122012 3120 122064 3126
rect 122012 3062 122064 3068
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 120908 2984 120960 2990
rect 120908 2926 120960 2932
rect 120644 2774 120672 2926
rect 120226 2760 120304 2774
rect 120170 2751 120304 2760
rect 120184 2746 120304 2751
rect 120552 2746 120672 2774
rect 121104 2774 121132 3062
rect 122196 2984 122248 2990
rect 122196 2926 122248 2932
rect 121104 2746 121224 2774
rect 119986 2544 120042 2553
rect 119986 2479 120042 2488
rect 120184 2106 120212 2746
rect 120552 2446 120580 2746
rect 120540 2440 120592 2446
rect 120540 2382 120592 2388
rect 120816 2304 120868 2310
rect 120816 2246 120868 2252
rect 120172 2100 120224 2106
rect 120172 2042 120224 2048
rect 120828 1630 120856 2246
rect 120816 1624 120868 1630
rect 120816 1566 120868 1572
rect 121196 1222 121224 2746
rect 122208 2582 122236 2926
rect 123036 2689 123064 3334
rect 123022 2680 123078 2689
rect 123022 2615 123078 2624
rect 122196 2576 122248 2582
rect 122196 2518 122248 2524
rect 121368 2304 121420 2310
rect 121368 2246 121420 2252
rect 121380 2038 121408 2246
rect 121368 2032 121420 2038
rect 121368 1974 121420 1980
rect 123036 1766 123064 2615
rect 123024 1760 123076 1766
rect 123024 1702 123076 1708
rect 123220 1329 123248 7686
rect 123312 7342 123340 7958
rect 123300 7336 123352 7342
rect 123300 7278 123352 7284
rect 123300 6656 123352 6662
rect 123300 6598 123352 6604
rect 123312 6254 123340 6598
rect 123300 6248 123352 6254
rect 123300 6190 123352 6196
rect 123300 4140 123352 4146
rect 123496 4128 123524 8894
rect 123574 8664 123630 8673
rect 123574 8599 123630 8608
rect 123588 8498 123616 8599
rect 123576 8492 123628 8498
rect 123576 8434 123628 8440
rect 123680 7342 123708 10406
rect 123772 10198 123800 10406
rect 123760 10192 123812 10198
rect 123760 10134 123812 10140
rect 123852 9376 123904 9382
rect 123852 9318 123904 9324
rect 123760 8968 123812 8974
rect 123760 8910 123812 8916
rect 123772 8809 123800 8910
rect 123864 8838 123892 9318
rect 123852 8832 123904 8838
rect 123758 8800 123814 8809
rect 123852 8774 123904 8780
rect 123758 8735 123814 8744
rect 123668 7336 123720 7342
rect 123668 7278 123720 7284
rect 123852 6452 123904 6458
rect 123852 6394 123904 6400
rect 123864 6186 123892 6394
rect 123956 6254 123984 11455
rect 124232 11393 124260 11494
rect 124218 11384 124274 11393
rect 124218 11319 124274 11328
rect 124310 11248 124366 11257
rect 124310 11183 124366 11192
rect 124220 9104 124272 9110
rect 124220 9046 124272 9052
rect 124128 8288 124180 8294
rect 124128 8230 124180 8236
rect 124036 8084 124088 8090
rect 124036 8026 124088 8032
rect 124048 7818 124076 8026
rect 124036 7812 124088 7818
rect 124036 7754 124088 7760
rect 124140 7177 124168 8230
rect 124232 7886 124260 9046
rect 124220 7880 124272 7886
rect 124220 7822 124272 7828
rect 124324 7410 124352 11183
rect 124416 9926 124444 12406
rect 124876 12102 124904 12815
rect 125244 12646 125272 15286
rect 125506 15200 125562 16000
rect 126058 15200 126114 16000
rect 126610 15314 126666 16000
rect 126610 15286 126928 15314
rect 126610 15200 126666 15286
rect 125520 13530 125548 15200
rect 125690 14512 125746 14521
rect 125690 14447 125746 14456
rect 125508 13524 125560 13530
rect 125508 13466 125560 13472
rect 125600 13388 125652 13394
rect 125600 13330 125652 13336
rect 125324 13320 125376 13326
rect 125322 13288 125324 13297
rect 125376 13288 125378 13297
rect 125322 13223 125378 13232
rect 125324 12980 125376 12986
rect 125324 12922 125376 12928
rect 125232 12640 125284 12646
rect 125232 12582 125284 12588
rect 125336 12209 125364 12922
rect 125612 12434 125640 13330
rect 125520 12406 125640 12434
rect 125520 12238 125548 12406
rect 125600 12368 125652 12374
rect 125704 12322 125732 14447
rect 125876 14340 125928 14346
rect 125876 14282 125928 14288
rect 125652 12316 125732 12322
rect 125600 12310 125732 12316
rect 125612 12294 125732 12310
rect 125508 12232 125560 12238
rect 125322 12200 125378 12209
rect 125508 12174 125560 12180
rect 125322 12135 125378 12144
rect 124864 12096 124916 12102
rect 124864 12038 124916 12044
rect 124772 11144 124824 11150
rect 124772 11086 124824 11092
rect 124784 10985 124812 11086
rect 124770 10976 124826 10985
rect 124770 10911 124826 10920
rect 124404 9920 124456 9926
rect 124404 9862 124456 9868
rect 124416 9761 124444 9862
rect 124402 9752 124458 9761
rect 124402 9687 124458 9696
rect 124404 9580 124456 9586
rect 124404 9522 124456 9528
rect 124416 9489 124444 9522
rect 124402 9480 124458 9489
rect 124402 9415 124458 9424
rect 124404 8832 124456 8838
rect 124404 8774 124456 8780
rect 124416 8537 124444 8774
rect 124402 8528 124458 8537
rect 124402 8463 124458 8472
rect 124404 7948 124456 7954
rect 124404 7890 124456 7896
rect 124416 7478 124444 7890
rect 124876 7721 124904 12038
rect 125140 11892 125192 11898
rect 125140 11834 125192 11840
rect 124954 11792 125010 11801
rect 124954 11727 125010 11736
rect 125048 11756 125100 11762
rect 124968 11626 124996 11727
rect 125048 11698 125100 11704
rect 124956 11620 125008 11626
rect 124956 11562 125008 11568
rect 124954 11384 125010 11393
rect 124954 11319 125010 11328
rect 124968 8090 124996 11319
rect 125060 11014 125088 11698
rect 125152 11694 125180 11834
rect 125140 11688 125192 11694
rect 125140 11630 125192 11636
rect 125336 11132 125364 12135
rect 125506 11928 125562 11937
rect 125612 11898 125640 12294
rect 125506 11863 125562 11872
rect 125600 11892 125652 11898
rect 125520 11558 125548 11863
rect 125600 11834 125652 11840
rect 125508 11552 125560 11558
rect 125508 11494 125560 11500
rect 125692 11280 125744 11286
rect 125692 11222 125744 11228
rect 125407 11144 125459 11150
rect 125336 11104 125407 11132
rect 125407 11086 125459 11092
rect 125600 11144 125652 11150
rect 125600 11086 125652 11092
rect 125232 11076 125284 11082
rect 125284 11036 125364 11064
rect 125232 11018 125284 11024
rect 125048 11008 125100 11014
rect 125048 10950 125100 10956
rect 125232 10668 125284 10674
rect 125232 10610 125284 10616
rect 125140 8424 125192 8430
rect 125140 8366 125192 8372
rect 124956 8084 125008 8090
rect 124956 8026 125008 8032
rect 124862 7712 124918 7721
rect 124862 7647 124918 7656
rect 124404 7472 124456 7478
rect 124404 7414 124456 7420
rect 124312 7404 124364 7410
rect 124312 7346 124364 7352
rect 124220 7200 124272 7206
rect 124126 7168 124182 7177
rect 124048 7126 124126 7154
rect 123944 6248 123996 6254
rect 123944 6190 123996 6196
rect 123852 6180 123904 6186
rect 123852 6122 123904 6128
rect 123352 4100 123524 4128
rect 123300 4082 123352 4088
rect 123496 3602 123524 4100
rect 123300 3596 123352 3602
rect 123300 3538 123352 3544
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 123312 2650 123340 3538
rect 123390 3088 123446 3097
rect 123390 3023 123446 3032
rect 123404 2854 123432 3023
rect 123864 2854 123892 6122
rect 123956 5778 123984 6190
rect 123944 5772 123996 5778
rect 123944 5714 123996 5720
rect 124048 5030 124076 7126
rect 124220 7142 124272 7148
rect 124126 7103 124182 7112
rect 124232 7002 124260 7142
rect 124968 7018 124996 8026
rect 124220 6996 124272 7002
rect 124968 6990 125088 7018
rect 124220 6938 124272 6944
rect 124956 6860 125008 6866
rect 124956 6802 125008 6808
rect 124864 6792 124916 6798
rect 124864 6734 124916 6740
rect 124876 6322 124904 6734
rect 124864 6316 124916 6322
rect 124864 6258 124916 6264
rect 124402 6216 124458 6225
rect 124402 6151 124404 6160
rect 124456 6151 124458 6160
rect 124404 6122 124456 6128
rect 124220 6112 124272 6118
rect 124220 6054 124272 6060
rect 124232 5234 124260 6054
rect 124586 5808 124642 5817
rect 124968 5778 124996 6802
rect 124586 5743 124642 5752
rect 124956 5772 125008 5778
rect 124600 5574 124628 5743
rect 124956 5714 125008 5720
rect 125060 5658 125088 6990
rect 124968 5630 125088 5658
rect 124588 5568 124640 5574
rect 124588 5510 124640 5516
rect 124220 5228 124272 5234
rect 124220 5170 124272 5176
rect 124036 5024 124088 5030
rect 124036 4966 124088 4972
rect 124128 4684 124180 4690
rect 124128 4626 124180 4632
rect 123944 4616 123996 4622
rect 123944 4558 123996 4564
rect 123956 4146 123984 4558
rect 124140 4486 124168 4626
rect 124128 4480 124180 4486
rect 124128 4422 124180 4428
rect 124864 4480 124916 4486
rect 124864 4422 124916 4428
rect 123944 4140 123996 4146
rect 123944 4082 123996 4088
rect 123944 3596 123996 3602
rect 123944 3538 123996 3544
rect 123956 2854 123984 3538
rect 123392 2848 123444 2854
rect 123392 2790 123444 2796
rect 123852 2848 123904 2854
rect 123852 2790 123904 2796
rect 123944 2848 123996 2854
rect 123944 2790 123996 2796
rect 123300 2644 123352 2650
rect 123300 2586 123352 2592
rect 123852 2304 123904 2310
rect 123852 2246 123904 2252
rect 124404 2304 124456 2310
rect 124404 2246 124456 2252
rect 123864 1970 123892 2246
rect 124416 2106 124444 2246
rect 124404 2100 124456 2106
rect 124404 2042 124456 2048
rect 123852 1964 123904 1970
rect 123852 1906 123904 1912
rect 124416 1834 124444 2042
rect 124876 1970 124904 4422
rect 124968 2774 124996 5630
rect 125048 5568 125100 5574
rect 125048 5510 125100 5516
rect 125060 5302 125088 5510
rect 125048 5296 125100 5302
rect 125048 5238 125100 5244
rect 125152 5166 125180 8366
rect 125244 6866 125272 10610
rect 125232 6860 125284 6866
rect 125232 6802 125284 6808
rect 125232 6316 125284 6322
rect 125232 6258 125284 6264
rect 125048 5160 125100 5166
rect 125048 5102 125100 5108
rect 125140 5160 125192 5166
rect 125140 5102 125192 5108
rect 125060 4282 125088 5102
rect 125048 4276 125100 4282
rect 125244 4264 125272 6258
rect 125336 4758 125364 11036
rect 125612 10606 125640 11086
rect 125704 11082 125732 11222
rect 125692 11076 125744 11082
rect 125692 11018 125744 11024
rect 125784 11076 125836 11082
rect 125784 11018 125836 11024
rect 125690 10840 125746 10849
rect 125690 10775 125692 10784
rect 125744 10775 125746 10784
rect 125692 10746 125744 10752
rect 125692 10668 125744 10674
rect 125692 10610 125744 10616
rect 125600 10600 125652 10606
rect 125600 10542 125652 10548
rect 125600 10464 125652 10470
rect 125600 10406 125652 10412
rect 125612 10033 125640 10406
rect 125598 10024 125654 10033
rect 125598 9959 125654 9968
rect 125704 9674 125732 10610
rect 125612 9646 125732 9674
rect 125612 9382 125640 9646
rect 125692 9512 125744 9518
rect 125692 9454 125744 9460
rect 125600 9376 125652 9382
rect 125600 9318 125652 9324
rect 125704 8838 125732 9454
rect 125416 8832 125468 8838
rect 125416 8774 125468 8780
rect 125692 8832 125744 8838
rect 125692 8774 125744 8780
rect 125428 7478 125456 8774
rect 125416 7472 125468 7478
rect 125416 7414 125468 7420
rect 125416 7336 125468 7342
rect 125416 7278 125468 7284
rect 125428 6798 125456 7278
rect 125506 7168 125562 7177
rect 125506 7103 125562 7112
rect 125416 6792 125468 6798
rect 125416 6734 125468 6740
rect 125416 6656 125468 6662
rect 125416 6598 125468 6604
rect 125428 5642 125456 6598
rect 125416 5636 125468 5642
rect 125416 5578 125468 5584
rect 125520 5370 125548 7103
rect 125690 5808 125746 5817
rect 125690 5743 125746 5752
rect 125704 5574 125732 5743
rect 125796 5710 125824 11018
rect 125888 7750 125916 14282
rect 126072 13462 126100 15200
rect 126900 13530 126928 15286
rect 127162 15200 127218 16000
rect 127714 15314 127770 16000
rect 127714 15286 128032 15314
rect 127714 15200 127770 15286
rect 126888 13524 126940 13530
rect 126888 13466 126940 13472
rect 126060 13456 126112 13462
rect 126060 13398 126112 13404
rect 126334 13016 126390 13025
rect 126334 12951 126390 12960
rect 126888 12980 126940 12986
rect 125968 12912 126020 12918
rect 125968 12854 126020 12860
rect 125980 12646 126008 12854
rect 125968 12640 126020 12646
rect 125968 12582 126020 12588
rect 126060 12436 126112 12442
rect 126060 12378 126112 12384
rect 125968 11756 126020 11762
rect 125968 11698 126020 11704
rect 125980 9518 126008 11698
rect 125968 9512 126020 9518
rect 125968 9454 126020 9460
rect 125876 7744 125928 7750
rect 125876 7686 125928 7692
rect 125784 5704 125836 5710
rect 125784 5646 125836 5652
rect 125692 5568 125744 5574
rect 125888 5545 125916 7686
rect 125968 6656 126020 6662
rect 125968 6598 126020 6604
rect 125980 6497 126008 6598
rect 125966 6488 126022 6497
rect 125966 6423 126022 6432
rect 126072 5710 126100 12378
rect 126348 12102 126376 12951
rect 126888 12922 126940 12928
rect 126900 12782 126928 12922
rect 126980 12912 127032 12918
rect 126980 12854 127032 12860
rect 126888 12776 126940 12782
rect 126888 12718 126940 12724
rect 126704 12640 126756 12646
rect 126704 12582 126756 12588
rect 126520 12232 126572 12238
rect 126520 12174 126572 12180
rect 126336 12096 126388 12102
rect 126336 12038 126388 12044
rect 126244 11144 126296 11150
rect 126244 11086 126296 11092
rect 126150 10840 126206 10849
rect 126150 10775 126206 10784
rect 126164 10674 126192 10775
rect 126152 10668 126204 10674
rect 126152 10610 126204 10616
rect 126152 10464 126204 10470
rect 126152 10406 126204 10412
rect 126164 10266 126192 10406
rect 126152 10260 126204 10266
rect 126152 10202 126204 10208
rect 126150 10024 126206 10033
rect 126150 9959 126206 9968
rect 126164 9761 126192 9959
rect 126150 9752 126206 9761
rect 126150 9687 126206 9696
rect 126256 9382 126284 11086
rect 126348 10033 126376 12038
rect 126334 10024 126390 10033
rect 126334 9959 126390 9968
rect 126428 9920 126480 9926
rect 126428 9862 126480 9868
rect 126152 9376 126204 9382
rect 126152 9318 126204 9324
rect 126244 9376 126296 9382
rect 126244 9318 126296 9324
rect 126164 8430 126192 9318
rect 126256 8838 126284 9318
rect 126244 8832 126296 8838
rect 126244 8774 126296 8780
rect 126152 8424 126204 8430
rect 126152 8366 126204 8372
rect 126256 7750 126284 8774
rect 126440 8537 126468 9862
rect 126426 8528 126482 8537
rect 126426 8463 126482 8472
rect 126244 7744 126296 7750
rect 126244 7686 126296 7692
rect 126152 7200 126204 7206
rect 126152 7142 126204 7148
rect 126164 6662 126192 7142
rect 126152 6656 126204 6662
rect 126152 6598 126204 6604
rect 126164 6458 126192 6598
rect 126152 6452 126204 6458
rect 126152 6394 126204 6400
rect 126060 5704 126112 5710
rect 126060 5646 126112 5652
rect 126256 5574 126284 7686
rect 126336 7472 126388 7478
rect 126336 7414 126388 7420
rect 126348 7206 126376 7414
rect 126428 7336 126480 7342
rect 126428 7278 126480 7284
rect 126336 7200 126388 7206
rect 126336 7142 126388 7148
rect 126440 7002 126468 7278
rect 126532 7154 126560 12174
rect 126716 12102 126744 12582
rect 126992 12434 127020 12854
rect 127176 12442 127204 15200
rect 127348 13796 127400 13802
rect 127348 13738 127400 13744
rect 127360 13025 127388 13738
rect 127532 13728 127584 13734
rect 127532 13670 127584 13676
rect 127544 13394 127572 13670
rect 128004 13530 128032 15286
rect 128266 15200 128322 16000
rect 128818 15200 128874 16000
rect 129370 15200 129426 16000
rect 129922 15200 129978 16000
rect 130474 15200 130530 16000
rect 131026 15200 131082 16000
rect 131578 15314 131634 16000
rect 132130 15314 132186 16000
rect 131578 15286 131896 15314
rect 131578 15200 131634 15286
rect 127992 13524 128044 13530
rect 127992 13466 128044 13472
rect 127440 13388 127492 13394
rect 127440 13330 127492 13336
rect 127532 13388 127584 13394
rect 127532 13330 127584 13336
rect 127346 13016 127402 13025
rect 127346 12951 127402 12960
rect 127452 12918 127480 13330
rect 127716 13320 127768 13326
rect 127716 13262 127768 13268
rect 127900 13320 127952 13326
rect 127900 13262 127952 13268
rect 127348 12912 127400 12918
rect 127348 12854 127400 12860
rect 127440 12912 127492 12918
rect 127440 12854 127492 12860
rect 127164 12436 127216 12442
rect 126992 12406 127112 12434
rect 126796 12368 126848 12374
rect 126796 12310 126848 12316
rect 126704 12096 126756 12102
rect 126704 12038 126756 12044
rect 126808 10826 126836 12310
rect 126888 12096 126940 12102
rect 126888 12038 126940 12044
rect 126980 12096 127032 12102
rect 126980 12038 127032 12044
rect 126900 11082 126928 12038
rect 126992 11762 127020 12038
rect 126980 11756 127032 11762
rect 126980 11698 127032 11704
rect 126888 11076 126940 11082
rect 126888 11018 126940 11024
rect 126716 10798 126836 10826
rect 126612 9036 126664 9042
rect 126612 8978 126664 8984
rect 126624 8498 126652 8978
rect 126612 8492 126664 8498
rect 126612 8434 126664 8440
rect 126612 7336 126664 7342
rect 126610 7304 126612 7313
rect 126664 7304 126666 7313
rect 126610 7239 126666 7248
rect 126532 7126 126652 7154
rect 126428 6996 126480 7002
rect 126428 6938 126480 6944
rect 126336 6928 126388 6934
rect 126336 6870 126388 6876
rect 126244 5568 126296 5574
rect 125692 5510 125744 5516
rect 125874 5536 125930 5545
rect 126244 5510 126296 5516
rect 125874 5471 125930 5480
rect 125508 5364 125560 5370
rect 125508 5306 125560 5312
rect 125876 5092 125928 5098
rect 125876 5034 125928 5040
rect 125416 5024 125468 5030
rect 125416 4966 125468 4972
rect 125428 4758 125456 4966
rect 125324 4752 125376 4758
rect 125324 4694 125376 4700
rect 125416 4752 125468 4758
rect 125468 4712 125548 4740
rect 125416 4694 125468 4700
rect 125336 4570 125364 4694
rect 125336 4554 125456 4570
rect 125336 4548 125468 4554
rect 125336 4542 125416 4548
rect 125416 4490 125468 4496
rect 125244 4236 125364 4264
rect 125048 4218 125100 4224
rect 125336 4146 125364 4236
rect 125232 4140 125284 4146
rect 125232 4082 125284 4088
rect 125324 4140 125376 4146
rect 125324 4082 125376 4088
rect 125244 4049 125272 4082
rect 125230 4040 125286 4049
rect 125230 3975 125286 3984
rect 125244 2854 125272 3975
rect 125336 3534 125364 4082
rect 125520 4078 125548 4712
rect 125508 4072 125560 4078
rect 125508 4014 125560 4020
rect 125600 3664 125652 3670
rect 125600 3606 125652 3612
rect 125324 3528 125376 3534
rect 125324 3470 125376 3476
rect 125612 2990 125640 3606
rect 125600 2984 125652 2990
rect 125600 2926 125652 2932
rect 125888 2854 125916 5034
rect 125968 4752 126020 4758
rect 125968 4694 126020 4700
rect 125980 3534 126008 4694
rect 126152 4140 126204 4146
rect 126152 4082 126204 4088
rect 126060 4004 126112 4010
rect 126060 3946 126112 3952
rect 125968 3528 126020 3534
rect 125968 3470 126020 3476
rect 125968 3120 126020 3126
rect 125968 3062 126020 3068
rect 125980 2990 126008 3062
rect 125968 2984 126020 2990
rect 125968 2926 126020 2932
rect 126072 2854 126100 3946
rect 126164 3738 126192 4082
rect 126152 3732 126204 3738
rect 126152 3674 126204 3680
rect 125232 2848 125284 2854
rect 125232 2790 125284 2796
rect 125876 2848 125928 2854
rect 125876 2790 125928 2796
rect 126060 2848 126112 2854
rect 126060 2790 126112 2796
rect 124968 2746 125180 2774
rect 125152 2650 125180 2746
rect 126348 2650 126376 6870
rect 125140 2644 125192 2650
rect 125140 2586 125192 2592
rect 126336 2644 126388 2650
rect 126336 2586 126388 2592
rect 126348 2446 126376 2586
rect 126440 2582 126468 6938
rect 126520 6656 126572 6662
rect 126520 6598 126572 6604
rect 126532 6361 126560 6598
rect 126518 6352 126574 6361
rect 126518 6287 126574 6296
rect 126520 6180 126572 6186
rect 126520 6122 126572 6128
rect 126532 5846 126560 6122
rect 126520 5840 126572 5846
rect 126520 5782 126572 5788
rect 126520 5024 126572 5030
rect 126520 4966 126572 4972
rect 126532 4486 126560 4966
rect 126520 4480 126572 4486
rect 126520 4422 126572 4428
rect 126624 4321 126652 7126
rect 126716 6458 126744 10798
rect 126796 10736 126848 10742
rect 126796 10678 126848 10684
rect 126808 9926 126836 10678
rect 126888 10668 126940 10674
rect 126888 10610 126940 10616
rect 126980 10668 127032 10674
rect 127084 10656 127112 12406
rect 127164 12378 127216 12384
rect 127162 12336 127218 12345
rect 127162 12271 127218 12280
rect 127176 11762 127204 12271
rect 127360 11937 127388 12854
rect 127440 12232 127492 12238
rect 127728 12209 127756 13262
rect 127912 12238 127940 13262
rect 128280 12986 128308 15200
rect 128450 14376 128506 14385
rect 128450 14311 128506 14320
rect 128268 12980 128320 12986
rect 128268 12922 128320 12928
rect 127992 12776 128044 12782
rect 127992 12718 128044 12724
rect 128004 12374 128032 12718
rect 128464 12442 128492 14311
rect 128832 13462 128860 15200
rect 129096 14476 129148 14482
rect 129096 14418 129148 14424
rect 128912 14000 128964 14006
rect 128912 13942 128964 13948
rect 129004 14000 129056 14006
rect 129004 13942 129056 13948
rect 128820 13456 128872 13462
rect 128820 13398 128872 13404
rect 128728 13320 128780 13326
rect 128728 13262 128780 13268
rect 128636 13184 128688 13190
rect 128636 13126 128688 13132
rect 128648 12889 128676 13126
rect 128634 12880 128690 12889
rect 128634 12815 128690 12824
rect 128452 12436 128504 12442
rect 128452 12378 128504 12384
rect 127992 12368 128044 12374
rect 127992 12310 128044 12316
rect 128464 12306 128492 12378
rect 128452 12300 128504 12306
rect 128452 12242 128504 12248
rect 128544 12300 128596 12306
rect 128544 12242 128596 12248
rect 127900 12232 127952 12238
rect 127440 12174 127492 12180
rect 127714 12200 127770 12209
rect 127346 11928 127402 11937
rect 127346 11863 127402 11872
rect 127164 11756 127216 11762
rect 127164 11698 127216 11704
rect 127348 11756 127400 11762
rect 127348 11698 127400 11704
rect 127256 11688 127308 11694
rect 127256 11630 127308 11636
rect 127084 10628 127204 10656
rect 126980 10610 127032 10616
rect 126796 9920 126848 9926
rect 126796 9862 126848 9868
rect 126796 8424 126848 8430
rect 126796 8366 126848 8372
rect 126704 6452 126756 6458
rect 126704 6394 126756 6400
rect 126704 5568 126756 5574
rect 126704 5510 126756 5516
rect 126716 5234 126744 5510
rect 126808 5370 126836 8366
rect 126796 5364 126848 5370
rect 126796 5306 126848 5312
rect 126704 5228 126756 5234
rect 126704 5170 126756 5176
rect 126796 5092 126848 5098
rect 126796 5034 126848 5040
rect 126610 4312 126666 4321
rect 126610 4247 126666 4256
rect 126808 3194 126836 5034
rect 126900 3738 126928 10610
rect 126992 9110 127020 10610
rect 127070 10568 127126 10577
rect 127070 10503 127072 10512
rect 127124 10503 127126 10512
rect 127072 10474 127124 10480
rect 127072 9376 127124 9382
rect 127072 9318 127124 9324
rect 126980 9104 127032 9110
rect 126980 9046 127032 9052
rect 127084 7954 127112 9318
rect 127176 8090 127204 10628
rect 127268 8498 127296 11630
rect 127360 8498 127388 11698
rect 127256 8492 127308 8498
rect 127256 8434 127308 8440
rect 127348 8492 127400 8498
rect 127348 8434 127400 8440
rect 127164 8084 127216 8090
rect 127164 8026 127216 8032
rect 127072 7948 127124 7954
rect 127072 7890 127124 7896
rect 127072 7744 127124 7750
rect 127072 7686 127124 7692
rect 127084 7478 127112 7686
rect 127072 7472 127124 7478
rect 127072 7414 127124 7420
rect 127268 7342 127296 8434
rect 127256 7336 127308 7342
rect 127256 7278 127308 7284
rect 127070 6624 127126 6633
rect 127070 6559 127126 6568
rect 127084 5846 127112 6559
rect 127072 5840 127124 5846
rect 127072 5782 127124 5788
rect 126978 5400 127034 5409
rect 126978 5335 127034 5344
rect 126992 4690 127020 5335
rect 127072 5296 127124 5302
rect 127072 5238 127124 5244
rect 127162 5264 127218 5273
rect 126980 4684 127032 4690
rect 126980 4626 127032 4632
rect 126888 3732 126940 3738
rect 126888 3674 126940 3680
rect 127084 3618 127112 5238
rect 127162 5199 127164 5208
rect 127216 5199 127218 5208
rect 127164 5170 127216 5176
rect 127452 4010 127480 12174
rect 127900 12174 127952 12180
rect 127714 12135 127770 12144
rect 128360 11688 128412 11694
rect 128360 11630 128412 11636
rect 127900 11552 127952 11558
rect 127900 11494 127952 11500
rect 127912 11257 127940 11494
rect 127898 11248 127954 11257
rect 127898 11183 127954 11192
rect 127808 11144 127860 11150
rect 128084 11144 128136 11150
rect 127808 11086 127860 11092
rect 128082 11112 128084 11121
rect 128268 11144 128320 11150
rect 128136 11112 128138 11121
rect 127532 10464 127584 10470
rect 127532 10406 127584 10412
rect 127544 9674 127572 10406
rect 127544 9646 127664 9674
rect 127532 9512 127584 9518
rect 127532 9454 127584 9460
rect 127544 9042 127572 9454
rect 127532 9036 127584 9042
rect 127532 8978 127584 8984
rect 127636 8430 127664 9646
rect 127716 8832 127768 8838
rect 127716 8774 127768 8780
rect 127624 8424 127676 8430
rect 127624 8366 127676 8372
rect 127728 8362 127756 8774
rect 127716 8356 127768 8362
rect 127716 8298 127768 8304
rect 127820 7546 127848 11086
rect 128268 11086 128320 11092
rect 128082 11047 128138 11056
rect 128084 10668 128136 10674
rect 128084 10610 128136 10616
rect 127990 10568 128046 10577
rect 127990 10503 128046 10512
rect 127900 9580 127952 9586
rect 127900 9522 127952 9528
rect 127808 7540 127860 7546
rect 127808 7482 127860 7488
rect 127808 7336 127860 7342
rect 127808 7278 127860 7284
rect 127820 6662 127848 7278
rect 127808 6656 127860 6662
rect 127808 6598 127860 6604
rect 127532 6316 127584 6322
rect 127532 6258 127584 6264
rect 127544 5914 127572 6258
rect 127624 6112 127676 6118
rect 127624 6054 127676 6060
rect 127532 5908 127584 5914
rect 127532 5850 127584 5856
rect 127636 5710 127664 6054
rect 127624 5704 127676 5710
rect 127624 5646 127676 5652
rect 127820 5370 127848 6598
rect 127912 5710 127940 9522
rect 128004 6458 128032 10503
rect 128096 10130 128124 10610
rect 128176 10464 128228 10470
rect 128176 10406 128228 10412
rect 128188 10198 128216 10406
rect 128176 10192 128228 10198
rect 128176 10134 128228 10140
rect 128084 10124 128136 10130
rect 128084 10066 128136 10072
rect 128280 9382 128308 11086
rect 128372 10674 128400 11630
rect 128452 11552 128504 11558
rect 128452 11494 128504 11500
rect 128464 10674 128492 11494
rect 128360 10668 128412 10674
rect 128360 10610 128412 10616
rect 128452 10668 128504 10674
rect 128452 10610 128504 10616
rect 128372 10198 128400 10610
rect 128360 10192 128412 10198
rect 128360 10134 128412 10140
rect 128268 9376 128320 9382
rect 128268 9318 128320 9324
rect 128268 9172 128320 9178
rect 128268 9114 128320 9120
rect 128280 9081 128308 9114
rect 128266 9072 128322 9081
rect 128266 9007 128322 9016
rect 128556 8838 128584 12242
rect 128636 11756 128688 11762
rect 128636 11698 128688 11704
rect 128648 10985 128676 11698
rect 128740 11558 128768 13262
rect 128820 13184 128872 13190
rect 128820 13126 128872 13132
rect 128832 12850 128860 13126
rect 128820 12844 128872 12850
rect 128820 12786 128872 12792
rect 128728 11552 128780 11558
rect 128728 11494 128780 11500
rect 128634 10976 128690 10985
rect 128634 10911 128690 10920
rect 128924 10674 128952 13942
rect 129016 12850 129044 13942
rect 129108 13190 129136 14418
rect 129384 14226 129412 15200
rect 129188 14204 129240 14210
rect 129384 14198 129688 14226
rect 129188 14146 129240 14152
rect 129096 13184 129148 13190
rect 129096 13126 129148 13132
rect 129004 12844 129056 12850
rect 129004 12786 129056 12792
rect 129108 12442 129136 13126
rect 129096 12436 129148 12442
rect 129096 12378 129148 12384
rect 129096 11348 129148 11354
rect 129200 11336 129228 14146
rect 129556 14136 129608 14142
rect 129556 14078 129608 14084
rect 129568 13297 129596 14078
rect 129554 13288 129610 13297
rect 129554 13223 129610 13232
rect 129568 12986 129596 13223
rect 129556 12980 129608 12986
rect 129660 12968 129688 14198
rect 129936 13530 129964 15200
rect 129924 13524 129976 13530
rect 129924 13466 129976 13472
rect 130384 13388 130436 13394
rect 130384 13330 130436 13336
rect 130108 13320 130160 13326
rect 130396 13297 130424 13330
rect 130108 13262 130160 13268
rect 130382 13288 130438 13297
rect 129740 12980 129792 12986
rect 129660 12940 129740 12968
rect 129556 12922 129608 12928
rect 129740 12922 129792 12928
rect 130016 12912 130068 12918
rect 130016 12854 130068 12860
rect 129924 12844 129976 12850
rect 129924 12786 129976 12792
rect 129936 12646 129964 12786
rect 129924 12640 129976 12646
rect 129924 12582 129976 12588
rect 130028 12238 130056 12854
rect 130120 12238 130148 13262
rect 130382 13223 130438 13232
rect 130488 12986 130516 15200
rect 130660 14612 130712 14618
rect 130660 14554 130712 14560
rect 130476 12980 130528 12986
rect 130476 12922 130528 12928
rect 130476 12844 130528 12850
rect 130476 12786 130528 12792
rect 130488 12442 130516 12786
rect 130568 12776 130620 12782
rect 130568 12718 130620 12724
rect 130476 12436 130528 12442
rect 130476 12378 130528 12384
rect 130198 12336 130254 12345
rect 130580 12322 130608 12718
rect 130672 12434 130700 14554
rect 131040 13512 131068 15200
rect 131120 13524 131172 13530
rect 131040 13484 131120 13512
rect 131120 13466 131172 13472
rect 131212 13184 131264 13190
rect 131212 13126 131264 13132
rect 131224 12986 131252 13126
rect 131302 13016 131358 13025
rect 131212 12980 131264 12986
rect 131868 12986 131896 15286
rect 132130 15286 132448 15314
rect 132130 15200 132186 15286
rect 132420 13512 132448 15286
rect 132682 15200 132738 16000
rect 133234 15200 133290 16000
rect 133786 15200 133842 16000
rect 134338 15200 134394 16000
rect 134890 15200 134946 16000
rect 135442 15314 135498 16000
rect 135994 15314 136050 16000
rect 135442 15286 135760 15314
rect 135442 15200 135498 15286
rect 132500 13524 132552 13530
rect 132420 13484 132500 13512
rect 132500 13466 132552 13472
rect 132696 13462 132724 15200
rect 132960 14408 133012 14414
rect 132960 14350 133012 14356
rect 132684 13456 132736 13462
rect 132684 13398 132736 13404
rect 131948 13320 132000 13326
rect 132408 13320 132460 13326
rect 132000 13280 132080 13308
rect 131948 13262 132000 13268
rect 131302 12951 131358 12960
rect 131856 12980 131908 12986
rect 131212 12922 131264 12928
rect 130672 12406 130884 12434
rect 130198 12271 130254 12280
rect 130488 12294 130608 12322
rect 130016 12232 130068 12238
rect 130016 12174 130068 12180
rect 130108 12232 130160 12238
rect 130108 12174 130160 12180
rect 130028 12073 130056 12174
rect 130014 12064 130070 12073
rect 130014 11999 130070 12008
rect 130212 11898 130240 12271
rect 130200 11892 130252 11898
rect 130200 11834 130252 11840
rect 129372 11824 129424 11830
rect 129372 11766 129424 11772
rect 129148 11308 129228 11336
rect 129280 11348 129332 11354
rect 129096 11290 129148 11296
rect 129280 11290 129332 11296
rect 128912 10668 128964 10674
rect 128912 10610 128964 10616
rect 129108 9353 129136 11290
rect 129094 9344 129150 9353
rect 129094 9279 129150 9288
rect 129292 9194 129320 11290
rect 129384 11150 129412 11766
rect 129372 11144 129424 11150
rect 129372 11086 129424 11092
rect 130200 11144 130252 11150
rect 130200 11086 130252 11092
rect 129372 11008 129424 11014
rect 129372 10950 129424 10956
rect 128924 9166 129320 9194
rect 128818 9072 128874 9081
rect 128818 9007 128874 9016
rect 128832 8974 128860 9007
rect 128820 8968 128872 8974
rect 128820 8910 128872 8916
rect 128544 8832 128596 8838
rect 128544 8774 128596 8780
rect 128082 8664 128138 8673
rect 128082 8599 128138 8608
rect 127992 6452 128044 6458
rect 127992 6394 128044 6400
rect 128096 6254 128124 8599
rect 128372 8486 128676 8514
rect 128372 8362 128400 8486
rect 128360 8356 128412 8362
rect 128360 8298 128412 8304
rect 128452 8356 128504 8362
rect 128452 8298 128504 8304
rect 128176 6792 128228 6798
rect 128176 6734 128228 6740
rect 128084 6248 128136 6254
rect 128084 6190 128136 6196
rect 128188 5953 128216 6734
rect 128360 6656 128412 6662
rect 128360 6598 128412 6604
rect 128268 6384 128320 6390
rect 128268 6326 128320 6332
rect 128280 6254 128308 6326
rect 128268 6248 128320 6254
rect 128268 6190 128320 6196
rect 128174 5944 128230 5953
rect 128372 5914 128400 6598
rect 128174 5879 128230 5888
rect 128360 5908 128412 5914
rect 128360 5850 128412 5856
rect 127900 5704 127952 5710
rect 127900 5646 127952 5652
rect 127808 5364 127860 5370
rect 127808 5306 127860 5312
rect 127820 4486 127848 5306
rect 127808 4480 127860 4486
rect 127808 4422 127860 4428
rect 127532 4276 127584 4282
rect 127532 4218 127584 4224
rect 127440 4004 127492 4010
rect 127440 3946 127492 3952
rect 127084 3590 127204 3618
rect 127072 3528 127124 3534
rect 127072 3470 127124 3476
rect 127084 3194 127112 3470
rect 126612 3188 126664 3194
rect 126612 3130 126664 3136
rect 126796 3188 126848 3194
rect 126796 3130 126848 3136
rect 127072 3188 127124 3194
rect 127072 3130 127124 3136
rect 126624 2990 126652 3130
rect 127084 3040 127112 3130
rect 126992 3012 127112 3040
rect 126612 2984 126664 2990
rect 126612 2926 126664 2932
rect 126428 2576 126480 2582
rect 126428 2518 126480 2524
rect 126336 2440 126388 2446
rect 126336 2382 126388 2388
rect 125324 2304 125376 2310
rect 125324 2246 125376 2252
rect 124864 1964 124916 1970
rect 124864 1906 124916 1912
rect 124404 1828 124456 1834
rect 124404 1770 124456 1776
rect 125336 1698 125364 2246
rect 125324 1692 125376 1698
rect 125324 1634 125376 1640
rect 125336 1494 125364 1634
rect 126992 1562 127020 3012
rect 127176 2774 127204 3590
rect 127544 3058 127572 4218
rect 127624 3936 127676 3942
rect 127624 3878 127676 3884
rect 127636 3398 127664 3878
rect 127716 3596 127768 3602
rect 127716 3538 127768 3544
rect 127728 3398 127756 3538
rect 127624 3392 127676 3398
rect 127624 3334 127676 3340
rect 127716 3392 127768 3398
rect 127716 3334 127768 3340
rect 127532 3052 127584 3058
rect 127532 2994 127584 3000
rect 127820 2990 127848 4422
rect 127912 3738 127940 5646
rect 128084 5364 128136 5370
rect 128084 5306 128136 5312
rect 128360 5364 128412 5370
rect 128360 5306 128412 5312
rect 128096 5234 128124 5306
rect 128084 5228 128136 5234
rect 128084 5170 128136 5176
rect 127992 5160 128044 5166
rect 127992 5102 128044 5108
rect 128004 4842 128032 5102
rect 128004 4814 128124 4842
rect 127992 4752 128044 4758
rect 127992 4694 128044 4700
rect 128004 4486 128032 4694
rect 127992 4480 128044 4486
rect 127992 4422 128044 4428
rect 127990 4312 128046 4321
rect 127990 4247 128046 4256
rect 128004 4146 128032 4247
rect 127992 4140 128044 4146
rect 127992 4082 128044 4088
rect 128096 4026 128124 4814
rect 128372 4706 128400 5306
rect 128188 4678 128400 4706
rect 128188 4214 128216 4678
rect 128176 4208 128228 4214
rect 128176 4150 128228 4156
rect 128268 4208 128320 4214
rect 128268 4150 128320 4156
rect 128280 4026 128308 4150
rect 128096 3998 128308 4026
rect 127992 3936 128044 3942
rect 127992 3878 128044 3884
rect 128004 3738 128032 3878
rect 128358 3768 128414 3777
rect 127900 3732 127952 3738
rect 127900 3674 127952 3680
rect 127992 3732 128044 3738
rect 128358 3703 128414 3712
rect 127992 3674 128044 3680
rect 128372 3534 128400 3703
rect 128360 3528 128412 3534
rect 128360 3470 128412 3476
rect 127900 3188 127952 3194
rect 127900 3130 127952 3136
rect 127808 2984 127860 2990
rect 127808 2926 127860 2932
rect 127912 2854 127940 3130
rect 127900 2848 127952 2854
rect 127900 2790 127952 2796
rect 127084 2746 127204 2774
rect 127084 2650 127112 2746
rect 127072 2644 127124 2650
rect 127072 2586 127124 2592
rect 126980 1556 127032 1562
rect 126980 1498 127032 1504
rect 125324 1488 125376 1494
rect 125324 1430 125376 1436
rect 123206 1320 123262 1329
rect 123206 1255 123262 1264
rect 121184 1216 121236 1222
rect 121184 1158 121236 1164
rect 119804 1148 119856 1154
rect 119804 1090 119856 1096
rect 128464 1086 128492 8298
rect 128542 7304 128598 7313
rect 128542 7239 128598 7248
rect 128556 6934 128584 7239
rect 128544 6928 128596 6934
rect 128544 6870 128596 6876
rect 128556 6458 128584 6870
rect 128544 6452 128596 6458
rect 128544 6394 128596 6400
rect 128544 6112 128596 6118
rect 128544 6054 128596 6060
rect 128556 5574 128584 6054
rect 128544 5568 128596 5574
rect 128544 5510 128596 5516
rect 128648 4049 128676 8486
rect 128924 8242 128952 9166
rect 129096 9104 129148 9110
rect 129096 9046 129148 9052
rect 128832 8214 128952 8242
rect 128728 6860 128780 6866
rect 128728 6802 128780 6808
rect 128740 6118 128768 6802
rect 128728 6112 128780 6118
rect 128728 6054 128780 6060
rect 128634 4040 128690 4049
rect 128634 3975 128690 3984
rect 128832 2854 128860 8214
rect 128910 8120 128966 8129
rect 128910 8055 128966 8064
rect 128924 7721 128952 8055
rect 128910 7712 128966 7721
rect 128910 7647 128966 7656
rect 128912 7540 128964 7546
rect 128912 7482 128964 7488
rect 128924 7410 128952 7482
rect 128912 7404 128964 7410
rect 128912 7346 128964 7352
rect 129108 6798 129136 9046
rect 129280 7812 129332 7818
rect 129280 7754 129332 7760
rect 129186 7712 129242 7721
rect 129186 7647 129242 7656
rect 129096 6792 129148 6798
rect 129096 6734 129148 6740
rect 129094 6352 129150 6361
rect 129094 6287 129150 6296
rect 129108 5846 129136 6287
rect 129096 5840 129148 5846
rect 129096 5782 129148 5788
rect 129200 5370 129228 7647
rect 129292 7478 129320 7754
rect 129384 7546 129412 10950
rect 130212 10810 130240 11086
rect 130384 11076 130436 11082
rect 130384 11018 130436 11024
rect 130200 10804 130252 10810
rect 130200 10746 130252 10752
rect 130200 10464 130252 10470
rect 130200 10406 130252 10412
rect 130292 10464 130344 10470
rect 130292 10406 130344 10412
rect 129646 10296 129702 10305
rect 129646 10231 129702 10240
rect 129660 9450 129688 10231
rect 130212 10130 130240 10406
rect 130200 10124 130252 10130
rect 130200 10066 130252 10072
rect 129740 10056 129792 10062
rect 129740 9998 129792 10004
rect 130016 10056 130068 10062
rect 130016 9998 130068 10004
rect 129648 9444 129700 9450
rect 129648 9386 129700 9392
rect 129556 8900 129608 8906
rect 129556 8842 129608 8848
rect 129372 7540 129424 7546
rect 129372 7482 129424 7488
rect 129280 7472 129332 7478
rect 129568 7426 129596 8842
rect 129648 8288 129700 8294
rect 129648 8230 129700 8236
rect 129660 8022 129688 8230
rect 129648 8016 129700 8022
rect 129648 7958 129700 7964
rect 129646 7576 129702 7585
rect 129646 7511 129702 7520
rect 129280 7414 129332 7420
rect 129476 7398 129596 7426
rect 129372 6724 129424 6730
rect 129372 6666 129424 6672
rect 129280 6656 129332 6662
rect 129280 6598 129332 6604
rect 129292 6322 129320 6598
rect 129384 6322 129412 6666
rect 129280 6316 129332 6322
rect 129280 6258 129332 6264
rect 129372 6316 129424 6322
rect 129372 6258 129424 6264
rect 129188 5364 129240 5370
rect 129188 5306 129240 5312
rect 128910 4720 128966 4729
rect 128910 4655 128966 4664
rect 129372 4684 129424 4690
rect 128924 4554 128952 4655
rect 129372 4626 129424 4632
rect 128912 4548 128964 4554
rect 128912 4490 128964 4496
rect 129004 3936 129056 3942
rect 129004 3878 129056 3884
rect 129016 3618 129044 3878
rect 129016 3590 129228 3618
rect 128820 2848 128872 2854
rect 128820 2790 128872 2796
rect 129016 2378 129044 3590
rect 129200 3534 129228 3590
rect 129188 3528 129240 3534
rect 129188 3470 129240 3476
rect 129096 3460 129148 3466
rect 129096 3402 129148 3408
rect 129108 3194 129136 3402
rect 129096 3188 129148 3194
rect 129096 3130 129148 3136
rect 129108 2774 129136 3130
rect 129384 3058 129412 4626
rect 129476 3670 129504 7398
rect 129556 7336 129608 7342
rect 129556 7278 129608 7284
rect 129568 6458 129596 7278
rect 129556 6452 129608 6458
rect 129556 6394 129608 6400
rect 129660 5914 129688 7511
rect 129752 6089 129780 9998
rect 129922 7984 129978 7993
rect 129922 7919 129978 7928
rect 129936 7886 129964 7919
rect 129924 7880 129976 7886
rect 129924 7822 129976 7828
rect 129832 7404 129884 7410
rect 129832 7346 129884 7352
rect 129844 6866 129872 7346
rect 129936 7002 129964 7822
rect 129924 6996 129976 7002
rect 129924 6938 129976 6944
rect 129832 6860 129884 6866
rect 129832 6802 129884 6808
rect 129738 6080 129794 6089
rect 129738 6015 129794 6024
rect 129922 6080 129978 6089
rect 129922 6015 129978 6024
rect 129648 5908 129700 5914
rect 129648 5850 129700 5856
rect 129738 5536 129794 5545
rect 129738 5471 129794 5480
rect 129752 5370 129780 5471
rect 129740 5364 129792 5370
rect 129740 5306 129792 5312
rect 129832 5364 129884 5370
rect 129832 5306 129884 5312
rect 129752 5166 129780 5306
rect 129740 5160 129792 5166
rect 129740 5102 129792 5108
rect 129844 4554 129872 5306
rect 129832 4548 129884 4554
rect 129832 4490 129884 4496
rect 129936 4078 129964 6015
rect 129924 4072 129976 4078
rect 129924 4014 129976 4020
rect 129464 3664 129516 3670
rect 129464 3606 129516 3612
rect 129476 3398 129504 3606
rect 129740 3596 129792 3602
rect 129740 3538 129792 3544
rect 129752 3466 129780 3538
rect 129740 3460 129792 3466
rect 129740 3402 129792 3408
rect 129464 3392 129516 3398
rect 129464 3334 129516 3340
rect 129924 3392 129976 3398
rect 129924 3334 129976 3340
rect 129372 3052 129424 3058
rect 129372 2994 129424 3000
rect 129936 2922 129964 3334
rect 129924 2916 129976 2922
rect 129924 2858 129976 2864
rect 130028 2774 130056 9998
rect 130304 9654 130332 10406
rect 130292 9648 130344 9654
rect 130292 9590 130344 9596
rect 130200 9512 130252 9518
rect 130200 9454 130252 9460
rect 130292 9512 130344 9518
rect 130292 9454 130344 9460
rect 130108 7880 130160 7886
rect 130108 7822 130160 7828
rect 130120 5710 130148 7822
rect 130212 7546 130240 9454
rect 130304 8906 130332 9454
rect 130292 8900 130344 8906
rect 130292 8842 130344 8848
rect 130292 8560 130344 8566
rect 130292 8502 130344 8508
rect 130304 8362 130332 8502
rect 130292 8356 130344 8362
rect 130292 8298 130344 8304
rect 130292 8084 130344 8090
rect 130292 8026 130344 8032
rect 130200 7540 130252 7546
rect 130200 7482 130252 7488
rect 130304 7313 130332 8026
rect 130396 8022 130424 11018
rect 130384 8016 130436 8022
rect 130384 7958 130436 7964
rect 130290 7304 130346 7313
rect 130290 7239 130346 7248
rect 130200 6792 130252 6798
rect 130200 6734 130252 6740
rect 130212 6458 130240 6734
rect 130200 6452 130252 6458
rect 130200 6394 130252 6400
rect 130108 5704 130160 5710
rect 130108 5646 130160 5652
rect 130200 5636 130252 5642
rect 130200 5578 130252 5584
rect 130212 4593 130240 5578
rect 130198 4584 130254 4593
rect 130198 4519 130254 4528
rect 130488 3466 130516 12294
rect 130658 12200 130714 12209
rect 130658 12135 130714 12144
rect 130672 12102 130700 12135
rect 130660 12096 130712 12102
rect 130660 12038 130712 12044
rect 130672 11121 130700 12038
rect 130658 11112 130714 11121
rect 130658 11047 130714 11056
rect 130752 11076 130804 11082
rect 130752 11018 130804 11024
rect 130568 11008 130620 11014
rect 130568 10950 130620 10956
rect 130580 10674 130608 10950
rect 130568 10668 130620 10674
rect 130568 10610 130620 10616
rect 130580 10062 130608 10610
rect 130568 10056 130620 10062
rect 130568 9998 130620 10004
rect 130660 8288 130712 8294
rect 130660 8230 130712 8236
rect 130672 7886 130700 8230
rect 130660 7880 130712 7886
rect 130660 7822 130712 7828
rect 130568 7812 130620 7818
rect 130568 7754 130620 7760
rect 130580 6390 130608 7754
rect 130568 6384 130620 6390
rect 130568 6326 130620 6332
rect 130764 3505 130792 11018
rect 130856 9217 130884 12406
rect 131212 12096 131264 12102
rect 131212 12038 131264 12044
rect 131224 11937 131252 12038
rect 131210 11928 131266 11937
rect 131210 11863 131266 11872
rect 130936 11144 130988 11150
rect 130936 11086 130988 11092
rect 130948 10062 130976 11086
rect 130936 10056 130988 10062
rect 130936 9998 130988 10004
rect 130948 9654 130976 9998
rect 130936 9648 130988 9654
rect 130936 9590 130988 9596
rect 130842 9208 130898 9217
rect 130948 9178 130976 9590
rect 131120 9444 131172 9450
rect 131120 9386 131172 9392
rect 130842 9143 130898 9152
rect 130936 9172 130988 9178
rect 130856 9110 130884 9143
rect 130936 9114 130988 9120
rect 131028 9172 131080 9178
rect 131028 9114 131080 9120
rect 130844 9104 130896 9110
rect 130844 9046 130896 9052
rect 130844 8832 130896 8838
rect 130844 8774 130896 8780
rect 130856 7546 130884 8774
rect 131040 7857 131068 9114
rect 131132 9110 131160 9386
rect 131120 9104 131172 9110
rect 131118 9072 131120 9081
rect 131172 9072 131174 9081
rect 131118 9007 131174 9016
rect 131316 8634 131344 12951
rect 131856 12922 131908 12928
rect 131948 12980 132000 12986
rect 131948 12922 132000 12928
rect 131764 12300 131816 12306
rect 131764 12242 131816 12248
rect 131776 12102 131804 12242
rect 131764 12096 131816 12102
rect 131764 12038 131816 12044
rect 131776 10305 131804 12038
rect 131856 11552 131908 11558
rect 131856 11494 131908 11500
rect 131762 10296 131818 10305
rect 131762 10231 131818 10240
rect 131672 8968 131724 8974
rect 131672 8910 131724 8916
rect 131684 8634 131712 8910
rect 131304 8628 131356 8634
rect 131304 8570 131356 8576
rect 131672 8628 131724 8634
rect 131672 8570 131724 8576
rect 131304 8288 131356 8294
rect 131304 8230 131356 8236
rect 131026 7848 131082 7857
rect 131026 7783 131082 7792
rect 130844 7540 130896 7546
rect 130844 7482 130896 7488
rect 131212 7540 131264 7546
rect 131212 7482 131264 7488
rect 130844 7404 130896 7410
rect 130844 7346 130896 7352
rect 130856 7313 130884 7346
rect 130842 7304 130898 7313
rect 130842 7239 130898 7248
rect 130856 7002 130884 7239
rect 130844 6996 130896 7002
rect 130844 6938 130896 6944
rect 130936 6996 130988 7002
rect 130936 6938 130988 6944
rect 130948 6866 130976 6938
rect 130936 6860 130988 6866
rect 130936 6802 130988 6808
rect 130844 6248 130896 6254
rect 130844 6190 130896 6196
rect 130856 5710 130884 6190
rect 131224 6118 131252 7482
rect 131316 7342 131344 8230
rect 131304 7336 131356 7342
rect 131304 7278 131356 7284
rect 131316 6882 131344 7278
rect 131762 7168 131818 7177
rect 131762 7103 131818 7112
rect 131316 6854 131436 6882
rect 131212 6112 131264 6118
rect 131212 6054 131264 6060
rect 131224 5778 131252 6054
rect 131302 5944 131358 5953
rect 131302 5879 131358 5888
rect 131212 5772 131264 5778
rect 131212 5714 131264 5720
rect 130844 5704 130896 5710
rect 130844 5646 130896 5652
rect 131316 5642 131344 5879
rect 131304 5636 131356 5642
rect 131304 5578 131356 5584
rect 131028 5568 131080 5574
rect 131028 5510 131080 5516
rect 130844 5024 130896 5030
rect 130844 4966 130896 4972
rect 130856 4321 130884 4966
rect 130842 4312 130898 4321
rect 130842 4247 130898 4256
rect 130750 3496 130806 3505
rect 130476 3460 130528 3466
rect 130750 3431 130806 3440
rect 130476 3402 130528 3408
rect 130200 3052 130252 3058
rect 130200 2994 130252 3000
rect 130212 2961 130240 2994
rect 130198 2952 130254 2961
rect 130198 2887 130200 2896
rect 130252 2887 130254 2896
rect 130200 2858 130252 2864
rect 129108 2746 129228 2774
rect 130028 2746 130240 2774
rect 129004 2372 129056 2378
rect 129004 2314 129056 2320
rect 128544 2304 128596 2310
rect 128544 2246 128596 2252
rect 128556 2106 128584 2246
rect 128544 2100 128596 2106
rect 128544 2042 128596 2048
rect 129200 1086 129228 2746
rect 130212 2650 130240 2746
rect 130200 2644 130252 2650
rect 130200 2586 130252 2592
rect 129554 2544 129610 2553
rect 129554 2479 129556 2488
rect 129608 2479 129610 2488
rect 129556 2450 129608 2456
rect 130856 1834 130884 4247
rect 131040 3670 131068 5510
rect 131120 4480 131172 4486
rect 131120 4422 131172 4428
rect 131132 4185 131160 4422
rect 131118 4176 131174 4185
rect 131118 4111 131174 4120
rect 131028 3664 131080 3670
rect 131028 3606 131080 3612
rect 131132 3505 131160 4111
rect 131212 3596 131264 3602
rect 131212 3538 131264 3544
rect 131118 3496 131174 3505
rect 131224 3466 131252 3538
rect 131118 3431 131174 3440
rect 131212 3460 131264 3466
rect 131212 3402 131264 3408
rect 131120 2848 131172 2854
rect 131120 2790 131172 2796
rect 131132 2514 131160 2790
rect 131316 2553 131344 5578
rect 131408 5234 131436 6854
rect 131580 6384 131632 6390
rect 131580 6326 131632 6332
rect 131592 6186 131620 6326
rect 131580 6180 131632 6186
rect 131580 6122 131632 6128
rect 131488 6112 131540 6118
rect 131488 6054 131540 6060
rect 131500 5234 131528 6054
rect 131396 5228 131448 5234
rect 131396 5170 131448 5176
rect 131488 5228 131540 5234
rect 131488 5170 131540 5176
rect 131500 4758 131528 5170
rect 131488 4752 131540 4758
rect 131488 4694 131540 4700
rect 131592 3126 131620 6122
rect 131672 5160 131724 5166
rect 131672 5102 131724 5108
rect 131684 4214 131712 5102
rect 131776 4758 131804 7103
rect 131764 4752 131816 4758
rect 131764 4694 131816 4700
rect 131672 4208 131724 4214
rect 131672 4150 131724 4156
rect 131764 4140 131816 4146
rect 131764 4082 131816 4088
rect 131776 4010 131804 4082
rect 131764 4004 131816 4010
rect 131764 3946 131816 3952
rect 131868 3126 131896 11494
rect 131960 9178 131988 12922
rect 131948 9172 132000 9178
rect 131948 9114 132000 9120
rect 131948 8356 132000 8362
rect 131948 8298 132000 8304
rect 131960 7478 131988 8298
rect 132052 7546 132080 13280
rect 132408 13262 132460 13268
rect 132132 12232 132184 12238
rect 132132 12174 132184 12180
rect 132144 11558 132172 12174
rect 132420 12102 132448 13262
rect 132776 12776 132828 12782
rect 132776 12718 132828 12724
rect 132408 12096 132460 12102
rect 132408 12038 132460 12044
rect 132316 11892 132368 11898
rect 132316 11834 132368 11840
rect 132132 11552 132184 11558
rect 132132 11494 132184 11500
rect 132224 9444 132276 9450
rect 132224 9386 132276 9392
rect 132130 8936 132186 8945
rect 132130 8871 132132 8880
rect 132184 8871 132186 8880
rect 132132 8842 132184 8848
rect 132040 7540 132092 7546
rect 132040 7482 132092 7488
rect 131948 7472 132000 7478
rect 131948 7414 132000 7420
rect 132040 7200 132092 7206
rect 132040 7142 132092 7148
rect 131948 5636 132000 5642
rect 131948 5578 132000 5584
rect 131960 3194 131988 5578
rect 132052 5302 132080 7142
rect 132236 6254 132264 9386
rect 132328 8634 132356 11834
rect 132500 11688 132552 11694
rect 132500 11630 132552 11636
rect 132408 11552 132460 11558
rect 132408 11494 132460 11500
rect 132420 10674 132448 11494
rect 132512 11218 132540 11630
rect 132788 11354 132816 12718
rect 132776 11348 132828 11354
rect 132776 11290 132828 11296
rect 132500 11212 132552 11218
rect 132500 11154 132552 11160
rect 132408 10668 132460 10674
rect 132408 10610 132460 10616
rect 132684 10056 132736 10062
rect 132684 9998 132736 10004
rect 132592 9580 132644 9586
rect 132592 9522 132644 9528
rect 132500 9376 132552 9382
rect 132500 9318 132552 9324
rect 132512 9110 132540 9318
rect 132500 9104 132552 9110
rect 132500 9046 132552 9052
rect 132316 8628 132368 8634
rect 132316 8570 132368 8576
rect 132224 6248 132276 6254
rect 132224 6190 132276 6196
rect 132328 6118 132356 8570
rect 132604 8514 132632 9522
rect 132420 8498 132632 8514
rect 132408 8492 132632 8498
rect 132460 8486 132632 8492
rect 132408 8434 132460 8440
rect 132500 7336 132552 7342
rect 132500 7278 132552 7284
rect 132512 7206 132540 7278
rect 132500 7200 132552 7206
rect 132500 7142 132552 7148
rect 132316 6112 132368 6118
rect 132316 6054 132368 6060
rect 132316 5772 132368 5778
rect 132316 5714 132368 5720
rect 132040 5296 132092 5302
rect 132040 5238 132092 5244
rect 132328 5030 132356 5714
rect 132500 5160 132552 5166
rect 132500 5102 132552 5108
rect 132316 5024 132368 5030
rect 132316 4966 132368 4972
rect 132328 4690 132356 4966
rect 132316 4684 132368 4690
rect 132316 4626 132368 4632
rect 132512 4486 132540 5102
rect 132500 4480 132552 4486
rect 132500 4422 132552 4428
rect 132038 4176 132094 4185
rect 132038 4111 132094 4120
rect 132052 4078 132080 4111
rect 132040 4072 132092 4078
rect 132040 4014 132092 4020
rect 132512 3534 132540 4422
rect 132696 3534 132724 9998
rect 132776 9988 132828 9994
rect 132776 9930 132828 9936
rect 132788 8634 132816 9930
rect 132868 8832 132920 8838
rect 132868 8774 132920 8780
rect 132776 8628 132828 8634
rect 132776 8570 132828 8576
rect 132788 6866 132816 8570
rect 132880 7954 132908 8774
rect 132972 7954 133000 14350
rect 133052 13932 133104 13938
rect 133052 13874 133104 13880
rect 133064 12782 133092 13874
rect 133248 13530 133276 15200
rect 133236 13524 133288 13530
rect 133236 13466 133288 13472
rect 133142 13288 133198 13297
rect 133142 13223 133198 13232
rect 133604 13252 133656 13258
rect 133156 13190 133184 13223
rect 133604 13194 133656 13200
rect 133144 13184 133196 13190
rect 133144 13126 133196 13132
rect 133616 12986 133644 13194
rect 133800 12986 133828 15200
rect 134352 13530 134380 15200
rect 134616 14544 134668 14550
rect 134616 14486 134668 14492
rect 134524 14408 134576 14414
rect 134524 14350 134576 14356
rect 134340 13524 134392 13530
rect 134340 13466 134392 13472
rect 133880 13320 133932 13326
rect 133880 13262 133932 13268
rect 133604 12980 133656 12986
rect 133604 12922 133656 12928
rect 133788 12980 133840 12986
rect 133788 12922 133840 12928
rect 133144 12912 133196 12918
rect 133144 12854 133196 12860
rect 133052 12776 133104 12782
rect 133156 12753 133184 12854
rect 133052 12718 133104 12724
rect 133142 12744 133198 12753
rect 133142 12679 133198 12688
rect 133892 12374 133920 13262
rect 134156 12844 134208 12850
rect 134156 12786 134208 12792
rect 134340 12844 134392 12850
rect 134340 12786 134392 12792
rect 133880 12368 133932 12374
rect 133880 12310 133932 12316
rect 133144 12232 133196 12238
rect 133144 12174 133196 12180
rect 133970 12200 134026 12209
rect 133052 11552 133104 11558
rect 133050 11520 133052 11529
rect 133104 11520 133106 11529
rect 133050 11455 133106 11464
rect 133064 11354 133092 11455
rect 133052 11348 133104 11354
rect 133052 11290 133104 11296
rect 133156 11218 133184 12174
rect 133970 12135 134026 12144
rect 133328 12096 133380 12102
rect 133328 12038 133380 12044
rect 133236 11620 133288 11626
rect 133236 11562 133288 11568
rect 133144 11212 133196 11218
rect 133144 11154 133196 11160
rect 133052 10464 133104 10470
rect 133052 10406 133104 10412
rect 132868 7948 132920 7954
rect 132868 7890 132920 7896
rect 132960 7948 133012 7954
rect 132960 7890 133012 7896
rect 132960 7744 133012 7750
rect 132960 7686 133012 7692
rect 132868 6928 132920 6934
rect 132868 6870 132920 6876
rect 132776 6860 132828 6866
rect 132776 6802 132828 6808
rect 132776 6248 132828 6254
rect 132776 6190 132828 6196
rect 132788 3777 132816 6190
rect 132880 5914 132908 6870
rect 132972 6254 133000 7686
rect 133064 6798 133092 10406
rect 133156 9518 133184 11154
rect 133248 11150 133276 11562
rect 133236 11144 133288 11150
rect 133236 11086 133288 11092
rect 133144 9512 133196 9518
rect 133144 9454 133196 9460
rect 133144 8424 133196 8430
rect 133144 8366 133196 8372
rect 133156 7954 133184 8366
rect 133144 7948 133196 7954
rect 133144 7890 133196 7896
rect 133052 6792 133104 6798
rect 133052 6734 133104 6740
rect 133340 6730 133368 12038
rect 133420 11688 133472 11694
rect 133420 11630 133472 11636
rect 133432 9466 133460 11630
rect 133696 11076 133748 11082
rect 133696 11018 133748 11024
rect 133708 10470 133736 11018
rect 133696 10464 133748 10470
rect 133696 10406 133748 10412
rect 133708 10266 133736 10406
rect 133696 10260 133748 10266
rect 133696 10202 133748 10208
rect 133788 10260 133840 10266
rect 133788 10202 133840 10208
rect 133512 9920 133564 9926
rect 133512 9862 133564 9868
rect 133524 9586 133552 9862
rect 133800 9722 133828 10202
rect 133984 9926 134012 12135
rect 134168 10062 134196 12786
rect 134352 12753 134380 12786
rect 134338 12744 134394 12753
rect 134338 12679 134394 12688
rect 134432 11688 134484 11694
rect 134432 11630 134484 11636
rect 134444 11014 134472 11630
rect 134536 11354 134564 14350
rect 134524 11348 134576 11354
rect 134524 11290 134576 11296
rect 134432 11008 134484 11014
rect 134432 10950 134484 10956
rect 134536 10441 134564 11290
rect 134522 10432 134578 10441
rect 134522 10367 134578 10376
rect 134156 10056 134208 10062
rect 134156 9998 134208 10004
rect 134064 9988 134116 9994
rect 134064 9930 134116 9936
rect 133972 9920 134024 9926
rect 133972 9862 134024 9868
rect 133878 9752 133934 9761
rect 133788 9716 133840 9722
rect 133878 9687 133934 9696
rect 133788 9658 133840 9664
rect 133512 9580 133564 9586
rect 133512 9522 133564 9528
rect 133432 9438 133552 9466
rect 133524 8974 133552 9438
rect 133512 8968 133564 8974
rect 133512 8910 133564 8916
rect 133696 8968 133748 8974
rect 133696 8910 133748 8916
rect 133524 8838 133552 8910
rect 133512 8832 133564 8838
rect 133512 8774 133564 8780
rect 133524 7886 133552 8774
rect 133604 7948 133656 7954
rect 133604 7890 133656 7896
rect 133512 7880 133564 7886
rect 133512 7822 133564 7828
rect 133418 6896 133474 6905
rect 133418 6831 133474 6840
rect 133236 6724 133288 6730
rect 133236 6666 133288 6672
rect 133328 6724 133380 6730
rect 133328 6666 133380 6672
rect 132960 6248 133012 6254
rect 132960 6190 133012 6196
rect 133052 6248 133104 6254
rect 133052 6190 133104 6196
rect 132960 6112 133012 6118
rect 132960 6054 133012 6060
rect 132868 5908 132920 5914
rect 132868 5850 132920 5856
rect 132972 5778 133000 6054
rect 132960 5772 133012 5778
rect 132960 5714 133012 5720
rect 133064 5574 133092 6190
rect 133052 5568 133104 5574
rect 133052 5510 133104 5516
rect 133064 5030 133092 5510
rect 133052 5024 133104 5030
rect 133052 4966 133104 4972
rect 133064 4622 133092 4966
rect 133052 4616 133104 4622
rect 133052 4558 133104 4564
rect 133248 4282 133276 6666
rect 133432 6662 133460 6831
rect 133420 6656 133472 6662
rect 133420 6598 133472 6604
rect 133236 4276 133288 4282
rect 133236 4218 133288 4224
rect 133142 4176 133198 4185
rect 133142 4111 133198 4120
rect 132774 3768 132830 3777
rect 132774 3703 132830 3712
rect 132958 3632 133014 3641
rect 132958 3567 133014 3576
rect 132972 3534 133000 3567
rect 132500 3528 132552 3534
rect 132500 3470 132552 3476
rect 132684 3528 132736 3534
rect 132684 3470 132736 3476
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 132512 3194 132540 3470
rect 131948 3188 132000 3194
rect 131948 3130 132000 3136
rect 132500 3188 132552 3194
rect 132500 3130 132552 3136
rect 131580 3120 131632 3126
rect 131580 3062 131632 3068
rect 131856 3120 131908 3126
rect 131856 3062 131908 3068
rect 131592 2650 131620 3062
rect 133156 2854 133184 4111
rect 133524 3534 133552 7822
rect 133616 7002 133644 7890
rect 133708 7750 133736 8910
rect 133788 8832 133840 8838
rect 133788 8774 133840 8780
rect 133800 8294 133828 8774
rect 133788 8288 133840 8294
rect 133788 8230 133840 8236
rect 133800 7886 133828 8230
rect 133788 7880 133840 7886
rect 133788 7822 133840 7828
rect 133696 7744 133748 7750
rect 133696 7686 133748 7692
rect 133800 7274 133828 7822
rect 133892 7585 133920 9687
rect 133878 7576 133934 7585
rect 133878 7511 133934 7520
rect 133984 7426 134012 9862
rect 134076 9586 134104 9930
rect 134064 9580 134116 9586
rect 134064 9522 134116 9528
rect 134064 8288 134116 8294
rect 134064 8230 134116 8236
rect 133892 7398 134012 7426
rect 133788 7268 133840 7274
rect 133788 7210 133840 7216
rect 133800 7002 133828 7210
rect 133604 6996 133656 7002
rect 133604 6938 133656 6944
rect 133788 6996 133840 7002
rect 133788 6938 133840 6944
rect 133616 4622 133644 6938
rect 133788 6792 133840 6798
rect 133788 6734 133840 6740
rect 133696 6656 133748 6662
rect 133696 6598 133748 6604
rect 133604 4616 133656 4622
rect 133604 4558 133656 4564
rect 133616 4185 133644 4558
rect 133602 4176 133658 4185
rect 133602 4111 133658 4120
rect 133616 4078 133644 4111
rect 133604 4072 133656 4078
rect 133604 4014 133656 4020
rect 133708 3913 133736 6598
rect 133800 5574 133828 6734
rect 133892 6225 133920 7398
rect 133878 6216 133934 6225
rect 133878 6151 133934 6160
rect 133972 5908 134024 5914
rect 133972 5850 134024 5856
rect 133984 5710 134012 5850
rect 133972 5704 134024 5710
rect 133972 5646 134024 5652
rect 133788 5568 133840 5574
rect 133788 5510 133840 5516
rect 133970 4312 134026 4321
rect 133970 4247 134026 4256
rect 133984 4078 134012 4247
rect 133972 4072 134024 4078
rect 133972 4014 134024 4020
rect 133694 3904 133750 3913
rect 133694 3839 133750 3848
rect 133236 3528 133288 3534
rect 133236 3470 133288 3476
rect 133512 3528 133564 3534
rect 133512 3470 133564 3476
rect 133144 2848 133196 2854
rect 133144 2790 133196 2796
rect 131580 2644 131632 2650
rect 131580 2586 131632 2592
rect 131302 2544 131358 2553
rect 131120 2508 131172 2514
rect 133156 2514 133184 2790
rect 131302 2479 131358 2488
rect 133144 2508 133196 2514
rect 131120 2450 131172 2456
rect 133144 2450 133196 2456
rect 133248 2394 133276 3470
rect 133156 2378 133276 2394
rect 133144 2372 133276 2378
rect 133196 2366 133276 2372
rect 133144 2314 133196 2320
rect 134076 2281 134104 8230
rect 134340 8016 134392 8022
rect 134340 7958 134392 7964
rect 134352 7002 134380 7958
rect 134432 7744 134484 7750
rect 134432 7686 134484 7692
rect 134340 6996 134392 7002
rect 134340 6938 134392 6944
rect 134156 6724 134208 6730
rect 134156 6666 134208 6672
rect 134168 3233 134196 6666
rect 134248 6384 134300 6390
rect 134248 6326 134300 6332
rect 134260 4078 134288 6326
rect 134444 6225 134472 7686
rect 134430 6216 134486 6225
rect 134430 6151 134486 6160
rect 134524 5704 134576 5710
rect 134522 5672 134524 5681
rect 134576 5672 134578 5681
rect 134522 5607 134578 5616
rect 134628 4826 134656 14486
rect 134904 12986 134932 15200
rect 135732 13530 135760 15286
rect 135994 15286 136404 15314
rect 135994 15200 136050 15286
rect 136376 13530 136404 15286
rect 136546 15200 136602 16000
rect 137098 15200 137154 16000
rect 137650 15314 137706 16000
rect 137650 15286 137968 15314
rect 137650 15200 137706 15286
rect 135720 13524 135772 13530
rect 135720 13466 135772 13472
rect 136364 13524 136416 13530
rect 136364 13466 136416 13472
rect 135352 13388 135404 13394
rect 135352 13330 135404 13336
rect 135168 13184 135220 13190
rect 135168 13126 135220 13132
rect 134892 12980 134944 12986
rect 134892 12922 134944 12928
rect 134890 12880 134946 12889
rect 134890 12815 134946 12824
rect 134708 11348 134760 11354
rect 134708 11290 134760 11296
rect 134720 11082 134748 11290
rect 134708 11076 134760 11082
rect 134708 11018 134760 11024
rect 134708 9920 134760 9926
rect 134708 9862 134760 9868
rect 134720 8514 134748 9862
rect 134800 9376 134852 9382
rect 134904 9364 134932 12815
rect 135180 12594 135208 13126
rect 135364 12646 135392 13330
rect 135628 13320 135680 13326
rect 135628 13262 135680 13268
rect 136088 13320 136140 13326
rect 136088 13262 136140 13268
rect 135536 13184 135588 13190
rect 135536 13126 135588 13132
rect 135352 12640 135404 12646
rect 135180 12566 135300 12594
rect 135352 12582 135404 12588
rect 135076 12436 135128 12442
rect 135076 12378 135128 12384
rect 134984 11892 135036 11898
rect 134984 11834 135036 11840
rect 134996 11694 135024 11834
rect 134984 11688 135036 11694
rect 134984 11630 135036 11636
rect 135088 11014 135116 12378
rect 135272 11898 135300 12566
rect 135548 12442 135576 13126
rect 135536 12436 135588 12442
rect 135536 12378 135588 12384
rect 135352 12164 135404 12170
rect 135352 12106 135404 12112
rect 135260 11892 135312 11898
rect 135260 11834 135312 11840
rect 134984 11008 135036 11014
rect 134984 10950 135036 10956
rect 135076 11008 135128 11014
rect 135076 10950 135128 10956
rect 135166 10976 135222 10985
rect 134996 10470 135024 10950
rect 135166 10911 135222 10920
rect 134984 10464 135036 10470
rect 134984 10406 135036 10412
rect 134984 9580 135036 9586
rect 134984 9522 135036 9528
rect 134852 9336 134932 9364
rect 134800 9318 134852 9324
rect 134812 9178 134840 9318
rect 134800 9172 134852 9178
rect 134800 9114 134852 9120
rect 134720 8486 134840 8514
rect 134708 8424 134760 8430
rect 134708 8366 134760 8372
rect 134616 4820 134668 4826
rect 134616 4762 134668 4768
rect 134720 4706 134748 8366
rect 134812 7954 134840 8486
rect 134800 7948 134852 7954
rect 134800 7890 134852 7896
rect 134812 7410 134840 7890
rect 134800 7404 134852 7410
rect 134800 7346 134852 7352
rect 134800 5228 134852 5234
rect 134800 5170 134852 5176
rect 134812 5030 134840 5170
rect 134800 5024 134852 5030
rect 134800 4966 134852 4972
rect 134628 4678 134748 4706
rect 134248 4072 134300 4078
rect 134248 4014 134300 4020
rect 134154 3224 134210 3233
rect 134154 3159 134210 3168
rect 134628 2650 134656 4678
rect 134996 4078 135024 9522
rect 135180 9489 135208 10911
rect 135166 9480 135222 9489
rect 135166 9415 135222 9424
rect 135076 9172 135128 9178
rect 135076 9114 135128 9120
rect 135088 8974 135116 9114
rect 135076 8968 135128 8974
rect 135076 8910 135128 8916
rect 135076 6724 135128 6730
rect 135076 6666 135128 6672
rect 135088 6458 135116 6666
rect 135180 6662 135208 9415
rect 135260 8968 135312 8974
rect 135260 8910 135312 8916
rect 135272 8838 135300 8910
rect 135260 8832 135312 8838
rect 135260 8774 135312 8780
rect 135168 6656 135220 6662
rect 135168 6598 135220 6604
rect 135076 6452 135128 6458
rect 135076 6394 135128 6400
rect 135272 6118 135300 8774
rect 135364 8498 135392 12106
rect 135640 11336 135668 13262
rect 135720 12776 135772 12782
rect 135718 12744 135720 12753
rect 135772 12744 135774 12753
rect 135718 12679 135774 12688
rect 135904 12232 135956 12238
rect 135904 12174 135956 12180
rect 135720 11620 135772 11626
rect 135720 11562 135772 11568
rect 135548 11308 135668 11336
rect 135548 11082 135576 11308
rect 135536 11076 135588 11082
rect 135536 11018 135588 11024
rect 135548 10577 135576 11018
rect 135534 10568 135590 10577
rect 135534 10503 135590 10512
rect 135536 10464 135588 10470
rect 135536 10406 135588 10412
rect 135548 10062 135576 10406
rect 135444 10056 135496 10062
rect 135444 9998 135496 10004
rect 135536 10056 135588 10062
rect 135536 9998 135588 10004
rect 135352 8492 135404 8498
rect 135352 8434 135404 8440
rect 135352 7812 135404 7818
rect 135352 7754 135404 7760
rect 135364 7410 135392 7754
rect 135352 7404 135404 7410
rect 135352 7346 135404 7352
rect 135350 6352 135406 6361
rect 135350 6287 135406 6296
rect 135260 6112 135312 6118
rect 135260 6054 135312 6060
rect 135260 5908 135312 5914
rect 135364 5896 135392 6287
rect 135312 5868 135392 5896
rect 135260 5850 135312 5856
rect 135076 4820 135128 4826
rect 135076 4762 135128 4768
rect 134984 4072 135036 4078
rect 134984 4014 135036 4020
rect 134708 3392 134760 3398
rect 134708 3334 134760 3340
rect 134720 3194 134748 3334
rect 134708 3188 134760 3194
rect 134708 3130 134760 3136
rect 135088 2689 135116 4762
rect 135260 3936 135312 3942
rect 135260 3878 135312 3884
rect 135074 2680 135130 2689
rect 134616 2644 134668 2650
rect 135074 2615 135130 2624
rect 134616 2586 134668 2592
rect 135272 2310 135300 3878
rect 135352 3528 135404 3534
rect 135352 3470 135404 3476
rect 135364 3398 135392 3470
rect 135352 3392 135404 3398
rect 135352 3334 135404 3340
rect 135364 2514 135392 3334
rect 135456 3194 135484 9998
rect 135548 9450 135576 9998
rect 135628 9988 135680 9994
rect 135628 9930 135680 9936
rect 135640 9761 135668 9930
rect 135626 9752 135682 9761
rect 135626 9687 135682 9696
rect 135536 9444 135588 9450
rect 135536 9386 135588 9392
rect 135536 8832 135588 8838
rect 135536 8774 135588 8780
rect 135548 6934 135576 8774
rect 135732 8498 135760 11562
rect 135812 11076 135864 11082
rect 135812 11018 135864 11024
rect 135720 8492 135772 8498
rect 135720 8434 135772 8440
rect 135720 8356 135772 8362
rect 135720 8298 135772 8304
rect 135732 7886 135760 8298
rect 135720 7880 135772 7886
rect 135720 7822 135772 7828
rect 135628 7200 135680 7206
rect 135628 7142 135680 7148
rect 135536 6928 135588 6934
rect 135536 6870 135588 6876
rect 135548 5642 135576 6870
rect 135536 5636 135588 5642
rect 135536 5578 135588 5584
rect 135444 3188 135496 3194
rect 135444 3130 135496 3136
rect 135352 2508 135404 2514
rect 135352 2450 135404 2456
rect 135640 2446 135668 7142
rect 135732 5914 135760 7822
rect 135824 6798 135852 11018
rect 135812 6792 135864 6798
rect 135812 6734 135864 6740
rect 135916 6390 135944 12174
rect 136100 11082 136128 13262
rect 136560 12986 136588 15200
rect 136914 14104 136970 14113
rect 136914 14039 136970 14048
rect 136732 13388 136784 13394
rect 136732 13330 136784 13336
rect 136548 12980 136600 12986
rect 136548 12922 136600 12928
rect 136640 12844 136692 12850
rect 136640 12786 136692 12792
rect 136180 12776 136232 12782
rect 136180 12718 136232 12724
rect 136088 11076 136140 11082
rect 136088 11018 136140 11024
rect 136192 10810 136220 12718
rect 136652 12481 136680 12786
rect 136744 12617 136772 13330
rect 136730 12608 136786 12617
rect 136730 12543 136786 12552
rect 136638 12472 136694 12481
rect 136638 12407 136694 12416
rect 136928 12345 136956 14039
rect 137112 13530 137140 15200
rect 137100 13524 137152 13530
rect 137100 13466 137152 13472
rect 137940 12986 137968 15286
rect 138202 15200 138258 16000
rect 138754 15314 138810 16000
rect 138754 15286 138888 15314
rect 138754 15200 138810 15286
rect 138020 13932 138072 13938
rect 138020 13874 138072 13880
rect 137928 12980 137980 12986
rect 137928 12922 137980 12928
rect 137744 12844 137796 12850
rect 137744 12786 137796 12792
rect 137192 12436 137244 12442
rect 137192 12378 137244 12384
rect 136914 12336 136970 12345
rect 136914 12271 136970 12280
rect 136456 11756 136508 11762
rect 136376 11716 136456 11744
rect 136180 10804 136232 10810
rect 136180 10746 136232 10752
rect 136272 9988 136324 9994
rect 136192 9948 136272 9976
rect 135996 8968 136048 8974
rect 135996 8910 136048 8916
rect 136008 8838 136036 8910
rect 135996 8832 136048 8838
rect 135996 8774 136048 8780
rect 135994 8120 136050 8129
rect 135994 8055 136050 8064
rect 135904 6384 135956 6390
rect 135904 6326 135956 6332
rect 135720 5908 135772 5914
rect 135720 5850 135772 5856
rect 135720 5092 135772 5098
rect 135720 5034 135772 5040
rect 135732 4622 135760 5034
rect 135916 4826 135944 6326
rect 135904 4820 135956 4826
rect 135904 4762 135956 4768
rect 135720 4616 135772 4622
rect 135720 4558 135772 4564
rect 135732 4078 135760 4558
rect 135720 4072 135772 4078
rect 135720 4014 135772 4020
rect 136008 2961 136036 8055
rect 136088 6112 136140 6118
rect 136088 6054 136140 6060
rect 136100 4078 136128 6054
rect 136088 4072 136140 4078
rect 136088 4014 136140 4020
rect 135994 2952 136050 2961
rect 135994 2887 136050 2896
rect 136192 2774 136220 9948
rect 136272 9930 136324 9936
rect 136376 8673 136404 11716
rect 136456 11698 136508 11704
rect 136732 11688 136784 11694
rect 136732 11630 136784 11636
rect 136744 10690 136772 11630
rect 136928 10810 136956 12271
rect 137204 11830 137232 12378
rect 137192 11824 137244 11830
rect 137192 11766 137244 11772
rect 137008 11756 137060 11762
rect 137008 11698 137060 11704
rect 137020 11354 137048 11698
rect 137008 11348 137060 11354
rect 137008 11290 137060 11296
rect 137284 11212 137336 11218
rect 137284 11154 137336 11160
rect 136916 10804 136968 10810
rect 136916 10746 136968 10752
rect 136652 10662 136772 10690
rect 136652 10656 136680 10662
rect 136468 10628 136680 10656
rect 136468 9926 136496 10628
rect 136732 10600 136784 10606
rect 136638 10568 136694 10577
rect 136732 10542 136784 10548
rect 136638 10503 136694 10512
rect 136652 10470 136680 10503
rect 136548 10464 136600 10470
rect 136548 10406 136600 10412
rect 136640 10464 136692 10470
rect 136640 10406 136692 10412
rect 136456 9920 136508 9926
rect 136456 9862 136508 9868
rect 136560 9178 136588 10406
rect 136456 9172 136508 9178
rect 136456 9114 136508 9120
rect 136548 9172 136600 9178
rect 136548 9114 136600 9120
rect 136468 8974 136496 9114
rect 136456 8968 136508 8974
rect 136456 8910 136508 8916
rect 136456 8832 136508 8838
rect 136456 8774 136508 8780
rect 136362 8664 136418 8673
rect 136362 8599 136418 8608
rect 136468 8090 136496 8774
rect 136456 8084 136508 8090
rect 136456 8026 136508 8032
rect 136362 7848 136418 7857
rect 136362 7783 136364 7792
rect 136416 7783 136418 7792
rect 136364 7754 136416 7760
rect 136652 7449 136680 10406
rect 136744 9994 136772 10542
rect 137190 10296 137246 10305
rect 137190 10231 137246 10240
rect 136732 9988 136784 9994
rect 136732 9930 136784 9936
rect 136916 9716 136968 9722
rect 136916 9658 136968 9664
rect 136928 9450 136956 9658
rect 136916 9444 136968 9450
rect 136916 9386 136968 9392
rect 136928 8838 136956 9386
rect 136916 8832 136968 8838
rect 136916 8774 136968 8780
rect 136928 8430 136956 8774
rect 137204 8430 137232 10231
rect 136916 8424 136968 8430
rect 136916 8366 136968 8372
rect 137192 8424 137244 8430
rect 137192 8366 137244 8372
rect 136638 7440 136694 7449
rect 136638 7375 136694 7384
rect 136824 7268 136876 7274
rect 136824 7210 136876 7216
rect 136640 7200 136692 7206
rect 136640 7142 136692 7148
rect 136652 6798 136680 7142
rect 136640 6792 136692 6798
rect 136640 6734 136692 6740
rect 136652 6118 136680 6734
rect 136640 6112 136692 6118
rect 136640 6054 136692 6060
rect 136272 5908 136324 5914
rect 136272 5850 136324 5856
rect 136284 5574 136312 5850
rect 136652 5710 136680 6054
rect 136640 5704 136692 5710
rect 136640 5646 136692 5652
rect 136272 5568 136324 5574
rect 136272 5510 136324 5516
rect 136836 5234 136864 7210
rect 136928 6458 136956 8366
rect 137296 7478 137324 11154
rect 137652 10804 137704 10810
rect 137652 10746 137704 10752
rect 137664 10606 137692 10746
rect 137652 10600 137704 10606
rect 137652 10542 137704 10548
rect 137756 10266 137784 12786
rect 138032 12238 138060 13874
rect 138216 13530 138244 15200
rect 138480 14068 138532 14074
rect 138480 14010 138532 14016
rect 138204 13524 138256 13530
rect 138204 13466 138256 13472
rect 138388 13456 138440 13462
rect 138388 13398 138440 13404
rect 138112 13320 138164 13326
rect 138112 13262 138164 13268
rect 138020 12232 138072 12238
rect 138020 12174 138072 12180
rect 138124 12102 138152 13262
rect 138112 12096 138164 12102
rect 138112 12038 138164 12044
rect 138018 10840 138074 10849
rect 138018 10775 138074 10784
rect 138032 10674 138060 10775
rect 138020 10668 138072 10674
rect 138020 10610 138072 10616
rect 137744 10260 137796 10266
rect 137744 10202 137796 10208
rect 137560 10124 137612 10130
rect 137560 10066 137612 10072
rect 137572 9654 137600 10066
rect 137560 9648 137612 9654
rect 137560 9590 137612 9596
rect 137468 9580 137520 9586
rect 137468 9522 137520 9528
rect 137376 9376 137428 9382
rect 137480 9353 137508 9522
rect 138018 9480 138074 9489
rect 138018 9415 138074 9424
rect 137836 9376 137888 9382
rect 137376 9318 137428 9324
rect 137466 9344 137522 9353
rect 137388 9042 137416 9318
rect 137836 9318 137888 9324
rect 137466 9279 137522 9288
rect 137848 9178 137876 9318
rect 137926 9208 137982 9217
rect 137836 9172 137888 9178
rect 137926 9143 137982 9152
rect 137836 9114 137888 9120
rect 137376 9036 137428 9042
rect 137376 8978 137428 8984
rect 137560 9036 137612 9042
rect 137560 8978 137612 8984
rect 137374 8936 137430 8945
rect 137374 8871 137376 8880
rect 137428 8871 137430 8880
rect 137376 8842 137428 8848
rect 137468 8832 137520 8838
rect 137468 8774 137520 8780
rect 137480 8294 137508 8774
rect 137468 8288 137520 8294
rect 137468 8230 137520 8236
rect 137376 7744 137428 7750
rect 137376 7686 137428 7692
rect 137284 7472 137336 7478
rect 137098 7440 137154 7449
rect 137284 7414 137336 7420
rect 137098 7375 137154 7384
rect 137112 7177 137140 7375
rect 137098 7168 137154 7177
rect 137098 7103 137154 7112
rect 137282 7032 137338 7041
rect 137282 6967 137338 6976
rect 136916 6452 136968 6458
rect 136916 6394 136968 6400
rect 137008 5908 137060 5914
rect 137008 5850 137060 5856
rect 137020 5778 137048 5850
rect 137296 5846 137324 6967
rect 137284 5840 137336 5846
rect 137284 5782 137336 5788
rect 137008 5772 137060 5778
rect 137008 5714 137060 5720
rect 136916 5636 136968 5642
rect 136916 5578 136968 5584
rect 136928 5234 136956 5578
rect 137296 5302 137324 5782
rect 137388 5370 137416 7686
rect 137572 7546 137600 8978
rect 137848 8498 137876 9114
rect 137940 9110 137968 9143
rect 137928 9104 137980 9110
rect 137928 9046 137980 9052
rect 137836 8492 137888 8498
rect 137836 8434 137888 8440
rect 137836 8084 137888 8090
rect 137836 8026 137888 8032
rect 137744 7812 137796 7818
rect 137744 7754 137796 7760
rect 137560 7540 137612 7546
rect 137560 7482 137612 7488
rect 137756 5817 137784 7754
rect 137742 5808 137798 5817
rect 137742 5743 137798 5752
rect 137376 5364 137428 5370
rect 137376 5306 137428 5312
rect 137192 5296 137244 5302
rect 137192 5238 137244 5244
rect 137284 5296 137336 5302
rect 137284 5238 137336 5244
rect 136824 5228 136876 5234
rect 136824 5170 136876 5176
rect 136916 5228 136968 5234
rect 136916 5170 136968 5176
rect 136928 5030 136956 5170
rect 136916 5024 136968 5030
rect 136916 4966 136968 4972
rect 137204 3398 137232 5238
rect 137560 5024 137612 5030
rect 137560 4966 137612 4972
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136916 3392 136968 3398
rect 136916 3334 136968 3340
rect 137192 3392 137244 3398
rect 137192 3334 137244 3340
rect 136468 3194 136496 3334
rect 136364 3188 136416 3194
rect 136364 3130 136416 3136
rect 136456 3188 136508 3194
rect 136456 3130 136508 3136
rect 136376 2938 136404 3130
rect 136928 3058 136956 3334
rect 137296 3058 137324 3470
rect 137572 3126 137600 4966
rect 137652 4004 137704 4010
rect 137652 3946 137704 3952
rect 137664 3534 137692 3946
rect 137652 3528 137704 3534
rect 137652 3470 137704 3476
rect 137560 3120 137612 3126
rect 137756 3097 137784 5743
rect 137848 5370 137876 8026
rect 138032 7410 138060 9415
rect 138020 7404 138072 7410
rect 138020 7346 138072 7352
rect 137928 6996 137980 7002
rect 137928 6938 137980 6944
rect 137940 6905 137968 6938
rect 137926 6896 137982 6905
rect 137926 6831 137982 6840
rect 137928 6112 137980 6118
rect 137928 6054 137980 6060
rect 137940 5710 137968 6054
rect 137928 5704 137980 5710
rect 137928 5646 137980 5652
rect 137836 5364 137888 5370
rect 137836 5306 137888 5312
rect 137834 4584 137890 4593
rect 137834 4519 137890 4528
rect 137848 4078 137876 4519
rect 137926 4312 137982 4321
rect 137926 4247 137982 4256
rect 137940 4214 137968 4247
rect 137928 4208 137980 4214
rect 137928 4150 137980 4156
rect 137836 4072 137888 4078
rect 137836 4014 137888 4020
rect 138032 3670 138060 7346
rect 137928 3664 137980 3670
rect 137926 3632 137928 3641
rect 138020 3664 138072 3670
rect 137980 3632 137982 3641
rect 138020 3606 138072 3612
rect 137926 3567 137982 3576
rect 137560 3062 137612 3068
rect 137742 3088 137798 3097
rect 136916 3052 136968 3058
rect 136916 2994 136968 3000
rect 137284 3052 137336 3058
rect 137742 3023 137798 3032
rect 137284 2994 137336 3000
rect 136376 2910 136956 2938
rect 136928 2854 136956 2910
rect 136916 2848 136968 2854
rect 136916 2790 136968 2796
rect 136100 2746 136220 2774
rect 135628 2440 135680 2446
rect 135628 2382 135680 2388
rect 135260 2304 135312 2310
rect 134062 2272 134118 2281
rect 135260 2246 135312 2252
rect 134062 2207 134118 2216
rect 134076 2038 134104 2207
rect 134064 2032 134116 2038
rect 134064 1974 134116 1980
rect 130844 1828 130896 1834
rect 130844 1770 130896 1776
rect 136100 1630 136128 2746
rect 136638 2680 136694 2689
rect 137296 2650 137324 2994
rect 136638 2615 136694 2624
rect 137284 2644 137336 2650
rect 136652 2038 136680 2615
rect 137284 2586 137336 2592
rect 138018 2408 138074 2417
rect 138018 2343 138020 2352
rect 138072 2343 138074 2352
rect 138020 2314 138072 2320
rect 136640 2032 136692 2038
rect 136640 1974 136692 1980
rect 136088 1624 136140 1630
rect 136088 1566 136140 1572
rect 128452 1080 128504 1086
rect 128452 1022 128504 1028
rect 129188 1080 129240 1086
rect 129188 1022 129240 1028
rect 138124 1018 138152 12038
rect 138204 11688 138256 11694
rect 138204 11630 138256 11636
rect 138216 11558 138244 11630
rect 138204 11552 138256 11558
rect 138204 11494 138256 11500
rect 138216 9926 138244 11494
rect 138296 11144 138348 11150
rect 138296 11086 138348 11092
rect 138204 9920 138256 9926
rect 138204 9862 138256 9868
rect 138202 9208 138258 9217
rect 138202 9143 138204 9152
rect 138256 9143 138258 9152
rect 138204 9114 138256 9120
rect 138204 8492 138256 8498
rect 138204 8434 138256 8440
rect 138216 8090 138244 8434
rect 138204 8084 138256 8090
rect 138204 8026 138256 8032
rect 138204 6860 138256 6866
rect 138204 6802 138256 6808
rect 138216 6390 138244 6802
rect 138204 6384 138256 6390
rect 138204 6326 138256 6332
rect 138308 5846 138336 11086
rect 138400 6633 138428 13398
rect 138492 12434 138520 14010
rect 138756 14000 138808 14006
rect 138756 13942 138808 13948
rect 138662 13696 138718 13705
rect 138662 13631 138718 13640
rect 138572 13456 138624 13462
rect 138572 13398 138624 13404
rect 138584 12918 138612 13398
rect 138572 12912 138624 12918
rect 138572 12854 138624 12860
rect 138492 12406 138612 12434
rect 138480 11892 138532 11898
rect 138480 11834 138532 11840
rect 138492 11354 138520 11834
rect 138480 11348 138532 11354
rect 138480 11290 138532 11296
rect 138584 9625 138612 12406
rect 138676 11898 138704 13631
rect 138664 11892 138716 11898
rect 138664 11834 138716 11840
rect 138664 11756 138716 11762
rect 138664 11698 138716 11704
rect 138676 11286 138704 11698
rect 138664 11280 138716 11286
rect 138664 11222 138716 11228
rect 138768 10849 138796 13942
rect 138860 13530 138888 15286
rect 139306 15200 139362 16000
rect 139858 15200 139914 16000
rect 140410 15314 140466 16000
rect 140962 15314 141018 16000
rect 141514 15314 141570 16000
rect 140410 15286 140728 15314
rect 140410 15200 140466 15286
rect 139320 13818 139348 15200
rect 139320 13790 139440 13818
rect 139007 13628 139315 13637
rect 139007 13626 139013 13628
rect 139069 13626 139093 13628
rect 139149 13626 139173 13628
rect 139229 13626 139253 13628
rect 139309 13626 139315 13628
rect 139069 13574 139071 13626
rect 139251 13574 139253 13626
rect 139007 13572 139013 13574
rect 139069 13572 139093 13574
rect 139149 13572 139173 13574
rect 139229 13572 139253 13574
rect 139309 13572 139315 13574
rect 139007 13563 139315 13572
rect 138848 13524 138900 13530
rect 138848 13466 138900 13472
rect 139412 13410 139440 13790
rect 139584 13728 139636 13734
rect 139584 13670 139636 13676
rect 139412 13382 139532 13410
rect 139400 13320 139452 13326
rect 139400 13262 139452 13268
rect 139007 12540 139315 12549
rect 139007 12538 139013 12540
rect 139069 12538 139093 12540
rect 139149 12538 139173 12540
rect 139229 12538 139253 12540
rect 139309 12538 139315 12540
rect 139069 12486 139071 12538
rect 139251 12486 139253 12538
rect 139007 12484 139013 12486
rect 139069 12484 139093 12486
rect 139149 12484 139173 12486
rect 139229 12484 139253 12486
rect 139309 12484 139315 12486
rect 139007 12475 139315 12484
rect 139124 12096 139176 12102
rect 139124 12038 139176 12044
rect 139136 11762 139164 12038
rect 139124 11756 139176 11762
rect 139124 11698 139176 11704
rect 139007 11452 139315 11461
rect 139007 11450 139013 11452
rect 139069 11450 139093 11452
rect 139149 11450 139173 11452
rect 139229 11450 139253 11452
rect 139309 11450 139315 11452
rect 139069 11398 139071 11450
rect 139251 11398 139253 11450
rect 139007 11396 139013 11398
rect 139069 11396 139093 11398
rect 139149 11396 139173 11398
rect 139229 11396 139253 11398
rect 139309 11396 139315 11398
rect 139007 11387 139315 11396
rect 138754 10840 138810 10849
rect 138664 10804 138716 10810
rect 138754 10775 138756 10784
rect 138664 10746 138716 10752
rect 138808 10775 138810 10784
rect 138756 10746 138808 10752
rect 138676 10538 138704 10746
rect 138768 10715 138796 10746
rect 138664 10532 138716 10538
rect 138664 10474 138716 10480
rect 139007 10364 139315 10373
rect 139007 10362 139013 10364
rect 139069 10362 139093 10364
rect 139149 10362 139173 10364
rect 139229 10362 139253 10364
rect 139309 10362 139315 10364
rect 139069 10310 139071 10362
rect 139251 10310 139253 10362
rect 139007 10308 139013 10310
rect 139069 10308 139093 10310
rect 139149 10308 139173 10310
rect 139229 10308 139253 10310
rect 139309 10308 139315 10310
rect 139007 10299 139315 10308
rect 138664 9920 138716 9926
rect 138664 9862 138716 9868
rect 138570 9616 138626 9625
rect 138570 9551 138626 9560
rect 138676 9110 138704 9862
rect 139306 9616 139362 9625
rect 139306 9551 139362 9560
rect 138940 9512 138992 9518
rect 138860 9472 138940 9500
rect 138860 9353 138888 9472
rect 138940 9454 138992 9460
rect 139320 9450 139348 9551
rect 139308 9444 139360 9450
rect 139308 9386 139360 9392
rect 138846 9344 138902 9353
rect 138846 9279 138902 9288
rect 139007 9276 139315 9285
rect 139007 9274 139013 9276
rect 139069 9274 139093 9276
rect 139149 9274 139173 9276
rect 139229 9274 139253 9276
rect 139309 9274 139315 9276
rect 139069 9222 139071 9274
rect 139251 9222 139253 9274
rect 139007 9220 139013 9222
rect 139069 9220 139093 9222
rect 139149 9220 139173 9222
rect 139229 9220 139253 9222
rect 139309 9220 139315 9222
rect 139007 9211 139315 9220
rect 138664 9104 138716 9110
rect 138664 9046 138716 9052
rect 138676 8974 138704 9046
rect 138664 8968 138716 8974
rect 138664 8910 138716 8916
rect 138572 8356 138624 8362
rect 138572 8298 138624 8304
rect 138584 8090 138612 8298
rect 138664 8288 138716 8294
rect 138664 8230 138716 8236
rect 138572 8084 138624 8090
rect 138572 8026 138624 8032
rect 138480 7200 138532 7206
rect 138480 7142 138532 7148
rect 138386 6624 138442 6633
rect 138386 6559 138442 6568
rect 138296 5840 138348 5846
rect 138296 5782 138348 5788
rect 138308 4758 138336 5782
rect 138388 5364 138440 5370
rect 138388 5306 138440 5312
rect 138296 4752 138348 4758
rect 138296 4694 138348 4700
rect 138400 4622 138428 5306
rect 138388 4616 138440 4622
rect 138388 4558 138440 4564
rect 138294 4176 138350 4185
rect 138294 4111 138296 4120
rect 138348 4111 138350 4120
rect 138296 4082 138348 4088
rect 138308 3466 138336 4082
rect 138296 3460 138348 3466
rect 138296 3402 138348 3408
rect 138492 2514 138520 7142
rect 138584 7002 138612 8026
rect 138676 7954 138704 8230
rect 139007 8188 139315 8197
rect 139007 8186 139013 8188
rect 139069 8186 139093 8188
rect 139149 8186 139173 8188
rect 139229 8186 139253 8188
rect 139309 8186 139315 8188
rect 139069 8134 139071 8186
rect 139251 8134 139253 8186
rect 139007 8132 139013 8134
rect 139069 8132 139093 8134
rect 139149 8132 139173 8134
rect 139229 8132 139253 8134
rect 139309 8132 139315 8134
rect 139007 8123 139315 8132
rect 138664 7948 138716 7954
rect 138664 7890 138716 7896
rect 139216 7540 139268 7546
rect 139216 7482 139268 7488
rect 139228 7410 139256 7482
rect 139216 7404 139268 7410
rect 139216 7346 139268 7352
rect 138940 7200 138992 7206
rect 139228 7188 139256 7346
rect 138992 7160 139256 7188
rect 138940 7142 138992 7148
rect 139007 7100 139315 7109
rect 139007 7098 139013 7100
rect 139069 7098 139093 7100
rect 139149 7098 139173 7100
rect 139229 7098 139253 7100
rect 139309 7098 139315 7100
rect 139069 7046 139071 7098
rect 139251 7046 139253 7098
rect 139007 7044 139013 7046
rect 139069 7044 139093 7046
rect 139149 7044 139173 7046
rect 139229 7044 139253 7046
rect 139309 7044 139315 7046
rect 139007 7035 139315 7044
rect 138572 6996 138624 7002
rect 138572 6938 138624 6944
rect 138664 6316 138716 6322
rect 138664 6258 138716 6264
rect 138676 5574 138704 6258
rect 138940 6180 138992 6186
rect 138860 6140 138940 6168
rect 138860 5778 138888 6140
rect 138940 6122 138992 6128
rect 139007 6012 139315 6021
rect 139007 6010 139013 6012
rect 139069 6010 139093 6012
rect 139149 6010 139173 6012
rect 139229 6010 139253 6012
rect 139309 6010 139315 6012
rect 139069 5958 139071 6010
rect 139251 5958 139253 6010
rect 139007 5956 139013 5958
rect 139069 5956 139093 5958
rect 139149 5956 139173 5958
rect 139229 5956 139253 5958
rect 139309 5956 139315 5958
rect 139007 5947 139315 5956
rect 138848 5772 138900 5778
rect 138848 5714 138900 5720
rect 139308 5704 139360 5710
rect 139308 5646 139360 5652
rect 138664 5568 138716 5574
rect 138664 5510 138716 5516
rect 139320 5370 139348 5646
rect 139308 5364 139360 5370
rect 139308 5306 139360 5312
rect 138572 5228 138624 5234
rect 138572 5170 138624 5176
rect 138584 4826 138612 5170
rect 139007 4924 139315 4933
rect 139007 4922 139013 4924
rect 139069 4922 139093 4924
rect 139149 4922 139173 4924
rect 139229 4922 139253 4924
rect 139309 4922 139315 4924
rect 139069 4870 139071 4922
rect 139251 4870 139253 4922
rect 139007 4868 139013 4870
rect 139069 4868 139093 4870
rect 139149 4868 139173 4870
rect 139229 4868 139253 4870
rect 139309 4868 139315 4870
rect 139007 4859 139315 4868
rect 138572 4820 138624 4826
rect 138572 4762 138624 4768
rect 139032 4752 139084 4758
rect 139032 4694 139084 4700
rect 139044 4554 139072 4694
rect 139032 4548 139084 4554
rect 139032 4490 139084 4496
rect 139412 4010 139440 13262
rect 139504 12986 139532 13382
rect 139596 13258 139624 13670
rect 139872 13530 139900 15200
rect 140596 13796 140648 13802
rect 140596 13738 140648 13744
rect 139860 13524 139912 13530
rect 139860 13466 139912 13472
rect 139584 13252 139636 13258
rect 139584 13194 139636 13200
rect 139676 13252 139728 13258
rect 139676 13194 139728 13200
rect 139492 12980 139544 12986
rect 139492 12922 139544 12928
rect 139584 12844 139636 12850
rect 139584 12786 139636 12792
rect 139490 11384 139546 11393
rect 139490 11319 139546 11328
rect 139504 11150 139532 11319
rect 139492 11144 139544 11150
rect 139492 11086 139544 11092
rect 139492 10600 139544 10606
rect 139492 10542 139544 10548
rect 139504 9654 139532 10542
rect 139492 9648 139544 9654
rect 139492 9590 139544 9596
rect 139492 9512 139544 9518
rect 139492 9454 139544 9460
rect 139504 9110 139532 9454
rect 139492 9104 139544 9110
rect 139492 9046 139544 9052
rect 139504 8945 139532 9046
rect 139596 9042 139624 12786
rect 139584 9036 139636 9042
rect 139584 8978 139636 8984
rect 139490 8936 139546 8945
rect 139490 8871 139546 8880
rect 139688 8838 139716 13194
rect 140608 12986 140636 13738
rect 140700 13530 140728 15286
rect 140962 15286 141280 15314
rect 140962 15200 141018 15286
rect 141148 13796 141200 13802
rect 141148 13738 141200 13744
rect 140688 13524 140740 13530
rect 140688 13466 140740 13472
rect 141160 13462 141188 13738
rect 141252 13462 141280 15286
rect 141344 15286 141570 15314
rect 141148 13456 141200 13462
rect 141148 13398 141200 13404
rect 141240 13456 141292 13462
rect 141240 13398 141292 13404
rect 140780 13320 140832 13326
rect 140780 13262 140832 13268
rect 140872 13320 140924 13326
rect 140872 13262 140924 13268
rect 140596 12980 140648 12986
rect 140596 12922 140648 12928
rect 139950 12472 140006 12481
rect 139950 12407 140006 12416
rect 139964 11626 139992 12407
rect 140594 12336 140650 12345
rect 140594 12271 140650 12280
rect 140608 12238 140636 12271
rect 140504 12232 140556 12238
rect 140504 12174 140556 12180
rect 140596 12232 140648 12238
rect 140596 12174 140648 12180
rect 140044 12096 140096 12102
rect 140044 12038 140096 12044
rect 139952 11620 140004 11626
rect 139952 11562 140004 11568
rect 139768 11348 139820 11354
rect 139768 11290 139820 11296
rect 139780 10441 139808 11290
rect 139860 10804 139912 10810
rect 139860 10746 139912 10752
rect 139872 10470 139900 10746
rect 139860 10464 139912 10470
rect 139766 10432 139822 10441
rect 139860 10406 139912 10412
rect 139952 10464 140004 10470
rect 139952 10406 140004 10412
rect 139766 10367 139822 10376
rect 139858 10296 139914 10305
rect 139858 10231 139914 10240
rect 139768 9988 139820 9994
rect 139768 9930 139820 9936
rect 139780 9761 139808 9930
rect 139872 9926 139900 10231
rect 139860 9920 139912 9926
rect 139860 9862 139912 9868
rect 139766 9752 139822 9761
rect 139766 9687 139822 9696
rect 139860 9376 139912 9382
rect 139858 9344 139860 9353
rect 139912 9344 139914 9353
rect 139858 9279 139914 9288
rect 139768 9104 139820 9110
rect 139768 9046 139820 9052
rect 139676 8832 139728 8838
rect 139676 8774 139728 8780
rect 139780 8294 139808 9046
rect 139860 8424 139912 8430
rect 139860 8366 139912 8372
rect 139768 8288 139820 8294
rect 139768 8230 139820 8236
rect 139872 7818 139900 8366
rect 139860 7812 139912 7818
rect 139860 7754 139912 7760
rect 139768 7744 139820 7750
rect 139768 7686 139820 7692
rect 139492 7200 139544 7206
rect 139492 7142 139544 7148
rect 139674 7168 139730 7177
rect 139504 7002 139532 7142
rect 139674 7103 139730 7112
rect 139492 6996 139544 7002
rect 139492 6938 139544 6944
rect 139504 6662 139532 6938
rect 139688 6798 139716 7103
rect 139676 6792 139728 6798
rect 139676 6734 139728 6740
rect 139584 6724 139636 6730
rect 139584 6666 139636 6672
rect 139492 6656 139544 6662
rect 139492 6598 139544 6604
rect 139596 6089 139624 6666
rect 139676 6452 139728 6458
rect 139676 6394 139728 6400
rect 139688 6254 139716 6394
rect 139676 6248 139728 6254
rect 139676 6190 139728 6196
rect 139582 6080 139638 6089
rect 139582 6015 139638 6024
rect 139490 5264 139546 5273
rect 139490 5199 139546 5208
rect 139400 4004 139452 4010
rect 139400 3946 139452 3952
rect 139007 3836 139315 3845
rect 139007 3834 139013 3836
rect 139069 3834 139093 3836
rect 139149 3834 139173 3836
rect 139229 3834 139253 3836
rect 139309 3834 139315 3836
rect 139069 3782 139071 3834
rect 139251 3782 139253 3834
rect 139007 3780 139013 3782
rect 139069 3780 139093 3782
rect 139149 3780 139173 3782
rect 139229 3780 139253 3782
rect 139309 3780 139315 3782
rect 139007 3771 139315 3780
rect 138756 3732 138808 3738
rect 138756 3674 138808 3680
rect 138768 3466 138796 3674
rect 139504 3466 139532 5199
rect 139584 5024 139636 5030
rect 139582 4992 139584 5001
rect 139636 4992 139638 5001
rect 139582 4927 139638 4936
rect 138756 3460 138808 3466
rect 138756 3402 138808 3408
rect 139492 3460 139544 3466
rect 139492 3402 139544 3408
rect 139596 2774 139624 4927
rect 139688 3194 139716 6190
rect 139780 5234 139808 7686
rect 139872 7002 139900 7754
rect 139860 6996 139912 7002
rect 139860 6938 139912 6944
rect 139860 6656 139912 6662
rect 139860 6598 139912 6604
rect 139872 6458 139900 6598
rect 139860 6452 139912 6458
rect 139860 6394 139912 6400
rect 139860 6112 139912 6118
rect 139860 6054 139912 6060
rect 139872 5234 139900 6054
rect 139768 5228 139820 5234
rect 139768 5170 139820 5176
rect 139860 5228 139912 5234
rect 139860 5170 139912 5176
rect 139768 5024 139820 5030
rect 139768 4966 139820 4972
rect 139780 3942 139808 4966
rect 139964 4622 139992 10406
rect 140056 10062 140084 12038
rect 140228 11688 140280 11694
rect 140228 11630 140280 11636
rect 140044 10056 140096 10062
rect 140044 9998 140096 10004
rect 140240 9908 140268 11630
rect 140410 11112 140466 11121
rect 140410 11047 140466 11056
rect 140320 10668 140372 10674
rect 140320 10610 140372 10616
rect 140332 10266 140360 10610
rect 140320 10260 140372 10266
rect 140320 10202 140372 10208
rect 140320 9920 140372 9926
rect 140240 9880 140320 9908
rect 140320 9862 140372 9868
rect 140042 9616 140098 9625
rect 140042 9551 140044 9560
rect 140096 9551 140098 9560
rect 140044 9522 140096 9528
rect 140228 8016 140280 8022
rect 140056 7964 140228 7970
rect 140056 7958 140280 7964
rect 140056 7942 140268 7958
rect 140056 7206 140084 7942
rect 140332 7460 140360 9862
rect 140424 7818 140452 11047
rect 140516 10606 140544 12174
rect 140596 11144 140648 11150
rect 140596 11086 140648 11092
rect 140504 10600 140556 10606
rect 140504 10542 140556 10548
rect 140516 10266 140544 10542
rect 140504 10260 140556 10266
rect 140504 10202 140556 10208
rect 140608 10146 140636 11086
rect 140688 11076 140740 11082
rect 140688 11018 140740 11024
rect 140516 10118 140636 10146
rect 140412 7812 140464 7818
rect 140412 7754 140464 7760
rect 140240 7432 140360 7460
rect 140044 7200 140096 7206
rect 140044 7142 140096 7148
rect 140136 7200 140188 7206
rect 140136 7142 140188 7148
rect 140056 6118 140084 7142
rect 140148 6798 140176 7142
rect 140136 6792 140188 6798
rect 140136 6734 140188 6740
rect 140044 6112 140096 6118
rect 140044 6054 140096 6060
rect 140044 5840 140096 5846
rect 140044 5782 140096 5788
rect 140056 5642 140084 5782
rect 140044 5636 140096 5642
rect 140044 5578 140096 5584
rect 140240 5302 140268 7432
rect 140516 7392 140544 10118
rect 140700 9674 140728 11018
rect 140792 10810 140820 13262
rect 140780 10804 140832 10810
rect 140780 10746 140832 10752
rect 140792 9994 140820 10746
rect 140884 10198 140912 13262
rect 141344 12442 141372 15286
rect 141514 15200 141570 15286
rect 142066 15200 142122 16000
rect 142618 15200 142674 16000
rect 143170 15200 143226 16000
rect 143722 15200 143778 16000
rect 144274 15200 144330 16000
rect 144826 15200 144882 16000
rect 145378 15200 145434 16000
rect 145930 15200 145986 16000
rect 146482 15200 146538 16000
rect 147034 15200 147090 16000
rect 147586 15200 147642 16000
rect 148138 15314 148194 16000
rect 148138 15286 148456 15314
rect 148138 15200 148194 15286
rect 141884 14816 141936 14822
rect 141884 14758 141936 14764
rect 141516 13524 141568 13530
rect 141516 13466 141568 13472
rect 141528 12850 141556 13466
rect 141516 12844 141568 12850
rect 141516 12786 141568 12792
rect 141332 12436 141384 12442
rect 141332 12378 141384 12384
rect 141896 12374 141924 14758
rect 142080 12968 142108 15200
rect 142528 13524 142580 13530
rect 142528 13466 142580 13472
rect 142160 12980 142212 12986
rect 142080 12940 142160 12968
rect 142160 12922 142212 12928
rect 142540 12850 142568 13466
rect 142528 12844 142580 12850
rect 142528 12786 142580 12792
rect 142344 12708 142396 12714
rect 142344 12650 142396 12656
rect 141884 12368 141936 12374
rect 141884 12310 141936 12316
rect 141240 12232 141292 12238
rect 141240 12174 141292 12180
rect 141148 11552 141200 11558
rect 141148 11494 141200 11500
rect 141056 11076 141108 11082
rect 141056 11018 141108 11024
rect 140872 10192 140924 10198
rect 140872 10134 140924 10140
rect 140780 9988 140832 9994
rect 140780 9930 140832 9936
rect 140596 9648 140648 9654
rect 140700 9646 141004 9674
rect 140596 9590 140648 9596
rect 140608 9110 140636 9590
rect 140780 9376 140832 9382
rect 140780 9318 140832 9324
rect 140596 9104 140648 9110
rect 140596 9046 140648 9052
rect 140688 9104 140740 9110
rect 140688 9046 140740 9052
rect 140608 8838 140636 9046
rect 140596 8832 140648 8838
rect 140596 8774 140648 8780
rect 140700 8362 140728 9046
rect 140688 8356 140740 8362
rect 140688 8298 140740 8304
rect 140596 8288 140648 8294
rect 140596 8230 140648 8236
rect 140332 7364 140544 7392
rect 140228 5296 140280 5302
rect 140228 5238 140280 5244
rect 140044 5228 140096 5234
rect 140044 5170 140096 5176
rect 139952 4616 140004 4622
rect 140056 4593 140084 5170
rect 139952 4558 140004 4564
rect 140042 4584 140098 4593
rect 140042 4519 140098 4528
rect 139950 4176 140006 4185
rect 139860 4140 139912 4146
rect 139950 4111 140006 4120
rect 139860 4082 139912 4088
rect 139768 3936 139820 3942
rect 139768 3878 139820 3884
rect 139872 3398 139900 4082
rect 139964 4010 139992 4111
rect 139952 4004 140004 4010
rect 139952 3946 140004 3952
rect 140056 3942 140084 4519
rect 140136 4276 140188 4282
rect 140136 4218 140188 4224
rect 140148 4185 140176 4218
rect 140134 4176 140190 4185
rect 140332 4146 140360 7364
rect 140504 7268 140556 7274
rect 140504 7210 140556 7216
rect 140412 6112 140464 6118
rect 140412 6054 140464 6060
rect 140424 4978 140452 6054
rect 140516 5710 140544 7210
rect 140608 6118 140636 8230
rect 140688 7880 140740 7886
rect 140688 7822 140740 7828
rect 140700 6254 140728 7822
rect 140792 7177 140820 9318
rect 140976 8974 141004 9646
rect 140964 8968 141016 8974
rect 140964 8910 141016 8916
rect 140976 8430 141004 8910
rect 140964 8424 141016 8430
rect 140964 8366 141016 8372
rect 140976 7800 141004 8366
rect 141068 7954 141096 11018
rect 141160 10674 141188 11494
rect 141252 10985 141280 12174
rect 141424 12164 141476 12170
rect 141424 12106 141476 12112
rect 141884 12164 141936 12170
rect 141884 12106 141936 12112
rect 141330 11384 141386 11393
rect 141330 11319 141386 11328
rect 141344 11150 141372 11319
rect 141332 11144 141384 11150
rect 141332 11086 141384 11092
rect 141332 11008 141384 11014
rect 141238 10976 141294 10985
rect 141332 10950 141384 10956
rect 141238 10911 141294 10920
rect 141344 10810 141372 10950
rect 141332 10804 141384 10810
rect 141332 10746 141384 10752
rect 141240 10736 141292 10742
rect 141240 10678 141292 10684
rect 141148 10668 141200 10674
rect 141148 10610 141200 10616
rect 141148 9920 141200 9926
rect 141148 9862 141200 9868
rect 141056 7948 141108 7954
rect 141056 7890 141108 7896
rect 141056 7812 141108 7818
rect 140976 7772 141056 7800
rect 141056 7754 141108 7760
rect 141160 7721 141188 9862
rect 141146 7712 141202 7721
rect 141146 7647 141202 7656
rect 140872 7404 140924 7410
rect 140872 7346 140924 7352
rect 140778 7168 140834 7177
rect 140778 7103 140834 7112
rect 140780 6656 140832 6662
rect 140778 6624 140780 6633
rect 140832 6624 140834 6633
rect 140778 6559 140834 6568
rect 140688 6248 140740 6254
rect 140688 6190 140740 6196
rect 140596 6112 140648 6118
rect 140596 6054 140648 6060
rect 140504 5704 140556 5710
rect 140504 5646 140556 5652
rect 140780 5636 140832 5642
rect 140780 5578 140832 5584
rect 140594 5128 140650 5137
rect 140594 5063 140596 5072
rect 140648 5063 140650 5072
rect 140596 5034 140648 5040
rect 140424 4950 140636 4978
rect 140608 4622 140636 4950
rect 140792 4758 140820 5578
rect 140780 4752 140832 4758
rect 140780 4694 140832 4700
rect 140596 4616 140648 4622
rect 140596 4558 140648 4564
rect 140134 4111 140190 4120
rect 140320 4140 140372 4146
rect 140320 4082 140372 4088
rect 140044 3936 140096 3942
rect 140044 3878 140096 3884
rect 140504 3936 140556 3942
rect 140504 3878 140556 3884
rect 140516 3738 140544 3878
rect 140504 3732 140556 3738
rect 140504 3674 140556 3680
rect 139952 3528 140004 3534
rect 139952 3470 140004 3476
rect 139860 3392 139912 3398
rect 139860 3334 139912 3340
rect 139872 3194 139900 3334
rect 139964 3194 139992 3470
rect 140608 3398 140636 4558
rect 140686 4448 140742 4457
rect 140686 4383 140742 4392
rect 140700 3777 140728 4383
rect 140686 3768 140742 3777
rect 140686 3703 140742 3712
rect 140688 3460 140740 3466
rect 140688 3402 140740 3408
rect 140596 3392 140648 3398
rect 140596 3334 140648 3340
rect 139676 3188 139728 3194
rect 139676 3130 139728 3136
rect 139860 3188 139912 3194
rect 139860 3130 139912 3136
rect 139952 3188 140004 3194
rect 139952 3130 140004 3136
rect 140700 2854 140728 3402
rect 140688 2848 140740 2854
rect 140688 2790 140740 2796
rect 139007 2748 139315 2757
rect 139007 2746 139013 2748
rect 139069 2746 139093 2748
rect 139149 2746 139173 2748
rect 139229 2746 139253 2748
rect 139309 2746 139315 2748
rect 139596 2746 139808 2774
rect 139069 2694 139071 2746
rect 139251 2694 139253 2746
rect 139007 2692 139013 2694
rect 139069 2692 139093 2694
rect 139149 2692 139173 2694
rect 139229 2692 139253 2694
rect 139309 2692 139315 2694
rect 139007 2683 139315 2692
rect 139780 2650 139808 2746
rect 138664 2644 138716 2650
rect 138664 2586 138716 2592
rect 139768 2644 139820 2650
rect 139768 2586 139820 2592
rect 138480 2508 138532 2514
rect 138480 2450 138532 2456
rect 138676 2446 138704 2586
rect 138664 2440 138716 2446
rect 138664 2382 138716 2388
rect 140594 2408 140650 2417
rect 140884 2378 140912 7346
rect 141148 6928 141200 6934
rect 141148 6870 141200 6876
rect 141160 6361 141188 6870
rect 141252 6390 141280 10678
rect 141332 10668 141384 10674
rect 141332 10610 141384 10616
rect 141344 10470 141372 10610
rect 141332 10464 141384 10470
rect 141332 10406 141384 10412
rect 141332 8900 141384 8906
rect 141332 8842 141384 8848
rect 141344 8498 141372 8842
rect 141332 8492 141384 8498
rect 141332 8434 141384 8440
rect 141436 8022 141464 12106
rect 141516 11688 141568 11694
rect 141568 11648 141648 11676
rect 141516 11630 141568 11636
rect 141516 11552 141568 11558
rect 141516 11494 141568 11500
rect 141528 11354 141556 11494
rect 141516 11348 141568 11354
rect 141516 11290 141568 11296
rect 141528 11257 141556 11290
rect 141514 11248 141570 11257
rect 141620 11218 141648 11648
rect 141514 11183 141570 11192
rect 141608 11212 141660 11218
rect 141608 11154 141660 11160
rect 141608 11076 141660 11082
rect 141608 11018 141660 11024
rect 141620 9058 141648 11018
rect 141700 9512 141752 9518
rect 141752 9472 141832 9500
rect 141700 9454 141752 9460
rect 141528 9030 141648 9058
rect 141528 8974 141556 9030
rect 141516 8968 141568 8974
rect 141516 8910 141568 8916
rect 141804 8673 141832 9472
rect 141790 8664 141846 8673
rect 141790 8599 141846 8608
rect 141516 8492 141568 8498
rect 141516 8434 141568 8440
rect 141424 8016 141476 8022
rect 141424 7958 141476 7964
rect 141332 7948 141384 7954
rect 141332 7890 141384 7896
rect 141344 7449 141372 7890
rect 141330 7440 141386 7449
rect 141330 7375 141386 7384
rect 141422 6896 141478 6905
rect 141422 6831 141478 6840
rect 141240 6384 141292 6390
rect 141146 6352 141202 6361
rect 141240 6326 141292 6332
rect 141332 6384 141384 6390
rect 141332 6326 141384 6332
rect 141146 6287 141202 6296
rect 141344 5914 141372 6326
rect 141332 5908 141384 5914
rect 141332 5850 141384 5856
rect 141148 5228 141200 5234
rect 141148 5170 141200 5176
rect 140964 5160 141016 5166
rect 141016 5120 141096 5148
rect 140964 5102 141016 5108
rect 141068 4593 141096 5120
rect 141054 4584 141110 4593
rect 141054 4519 141110 4528
rect 141068 4486 141096 4519
rect 141056 4480 141108 4486
rect 141056 4422 141108 4428
rect 141160 4282 141188 5170
rect 141436 4486 141464 6831
rect 141528 5370 141556 8434
rect 141608 8424 141660 8430
rect 141608 8366 141660 8372
rect 141516 5364 141568 5370
rect 141516 5306 141568 5312
rect 141424 4480 141476 4486
rect 141424 4422 141476 4428
rect 141148 4276 141200 4282
rect 141148 4218 141200 4224
rect 141056 4004 141108 4010
rect 141056 3946 141108 3952
rect 141068 3466 141096 3946
rect 141056 3460 141108 3466
rect 141056 3402 141108 3408
rect 141160 2774 141188 4218
rect 141424 3936 141476 3942
rect 141424 3878 141476 3884
rect 141436 3194 141464 3878
rect 141424 3188 141476 3194
rect 141424 3130 141476 3136
rect 141068 2746 141188 2774
rect 141068 2689 141096 2746
rect 141054 2680 141110 2689
rect 141620 2650 141648 8366
rect 141792 8356 141844 8362
rect 141792 8298 141844 8304
rect 141804 7546 141832 8298
rect 141792 7540 141844 7546
rect 141792 7482 141844 7488
rect 141790 4040 141846 4049
rect 141790 3975 141792 3984
rect 141844 3975 141846 3984
rect 141792 3946 141844 3952
rect 141700 3120 141752 3126
rect 141700 3062 141752 3068
rect 141054 2615 141110 2624
rect 141608 2644 141660 2650
rect 140594 2343 140650 2352
rect 140872 2372 140924 2378
rect 140608 2310 140636 2343
rect 140872 2314 140924 2320
rect 140596 2304 140648 2310
rect 141068 2281 141096 2615
rect 141608 2586 141660 2592
rect 141712 2378 141740 3062
rect 141896 2774 141924 12106
rect 142356 12102 142384 12650
rect 142632 12646 142660 15200
rect 142712 13184 142764 13190
rect 142712 13126 142764 13132
rect 142724 12850 142752 13126
rect 142712 12844 142764 12850
rect 142712 12786 142764 12792
rect 142620 12640 142672 12646
rect 142620 12582 142672 12588
rect 143184 12442 143212 15200
rect 143356 13320 143408 13326
rect 143356 13262 143408 13268
rect 143368 12918 143396 13262
rect 143356 12912 143408 12918
rect 143356 12854 143408 12860
rect 143172 12436 143224 12442
rect 143172 12378 143224 12384
rect 143264 12300 143316 12306
rect 143264 12242 143316 12248
rect 142344 12096 142396 12102
rect 143172 12096 143224 12102
rect 142344 12038 142396 12044
rect 143078 12064 143134 12073
rect 143172 12038 143224 12044
rect 143078 11999 143134 12008
rect 142618 11928 142674 11937
rect 142618 11863 142674 11872
rect 142160 10260 142212 10266
rect 142160 10202 142212 10208
rect 142172 9994 142200 10202
rect 142160 9988 142212 9994
rect 142160 9930 142212 9936
rect 142160 9376 142212 9382
rect 142160 9318 142212 9324
rect 142342 9344 142398 9353
rect 141976 8968 142028 8974
rect 141976 8910 142028 8916
rect 141988 8430 142016 8910
rect 141976 8424 142028 8430
rect 141976 8366 142028 8372
rect 142068 8288 142120 8294
rect 142068 8230 142120 8236
rect 142080 7993 142108 8230
rect 142066 7984 142122 7993
rect 142066 7919 142122 7928
rect 142066 7712 142122 7721
rect 142066 7647 142122 7656
rect 141976 7540 142028 7546
rect 141976 7482 142028 7488
rect 141988 7449 142016 7482
rect 141974 7440 142030 7449
rect 141974 7375 142030 7384
rect 141988 5545 142016 7375
rect 142080 7177 142108 7647
rect 142066 7168 142122 7177
rect 142066 7103 142122 7112
rect 142172 5953 142200 9318
rect 142342 9279 142398 9288
rect 142252 7744 142304 7750
rect 142252 7686 142304 7692
rect 142264 6633 142292 7686
rect 142356 7041 142384 9279
rect 142436 7744 142488 7750
rect 142436 7686 142488 7692
rect 142448 7546 142476 7686
rect 142436 7540 142488 7546
rect 142436 7482 142488 7488
rect 142342 7032 142398 7041
rect 142342 6967 142398 6976
rect 142356 6866 142384 6967
rect 142632 6866 142660 11863
rect 142988 11756 143040 11762
rect 142988 11698 143040 11704
rect 142896 11688 142948 11694
rect 142896 11630 142948 11636
rect 142908 10470 142936 11630
rect 143000 11150 143028 11698
rect 142988 11144 143040 11150
rect 142988 11086 143040 11092
rect 142896 10464 142948 10470
rect 142896 10406 142948 10412
rect 142908 10062 142936 10406
rect 142896 10056 142948 10062
rect 142896 9998 142948 10004
rect 142802 9888 142858 9897
rect 142802 9823 142858 9832
rect 142816 9217 142844 9823
rect 142802 9208 142858 9217
rect 142802 9143 142858 9152
rect 143092 8838 143120 11999
rect 143184 11665 143212 12038
rect 143170 11656 143226 11665
rect 143170 11591 143226 11600
rect 143276 11558 143304 12242
rect 143264 11552 143316 11558
rect 143262 11520 143264 11529
rect 143316 11520 143318 11529
rect 143262 11455 143318 11464
rect 143172 11008 143224 11014
rect 143172 10950 143224 10956
rect 142896 8832 142948 8838
rect 142896 8774 142948 8780
rect 143080 8832 143132 8838
rect 143080 8774 143132 8780
rect 142344 6860 142396 6866
rect 142344 6802 142396 6808
rect 142620 6860 142672 6866
rect 142620 6802 142672 6808
rect 142250 6624 142306 6633
rect 142250 6559 142306 6568
rect 142158 5944 142214 5953
rect 142158 5879 142214 5888
rect 141974 5536 142030 5545
rect 141974 5471 142030 5480
rect 142356 5234 142384 6802
rect 142436 5704 142488 5710
rect 142436 5646 142488 5652
rect 142344 5228 142396 5234
rect 142344 5170 142396 5176
rect 142356 3738 142384 5170
rect 142448 4808 142476 5646
rect 142632 5574 142660 6802
rect 142804 6792 142856 6798
rect 142804 6734 142856 6740
rect 142816 6322 142844 6734
rect 142908 6322 142936 8774
rect 143080 8492 143132 8498
rect 143080 8434 143132 8440
rect 143092 8106 143120 8434
rect 143000 8090 143120 8106
rect 142988 8084 143120 8090
rect 143040 8078 143120 8084
rect 142988 8026 143040 8032
rect 142988 7880 143040 7886
rect 142988 7822 143040 7828
rect 143080 7880 143132 7886
rect 143080 7822 143132 7828
rect 143000 7750 143028 7822
rect 142988 7744 143040 7750
rect 142988 7686 143040 7692
rect 143092 6798 143120 7822
rect 143080 6792 143132 6798
rect 143080 6734 143132 6740
rect 143080 6656 143132 6662
rect 143080 6598 143132 6604
rect 142804 6316 142856 6322
rect 142804 6258 142856 6264
rect 142896 6316 142948 6322
rect 142896 6258 142948 6264
rect 142816 5710 142844 6258
rect 142804 5704 142856 5710
rect 142804 5646 142856 5652
rect 142620 5568 142672 5574
rect 142620 5510 142672 5516
rect 142712 5364 142764 5370
rect 142712 5306 142764 5312
rect 142724 5030 142752 5306
rect 142816 5302 142844 5646
rect 143092 5574 143120 6598
rect 143080 5568 143132 5574
rect 143080 5510 143132 5516
rect 142804 5296 142856 5302
rect 142804 5238 142856 5244
rect 142712 5024 142764 5030
rect 142712 4966 142764 4972
rect 142448 4780 142660 4808
rect 142448 4690 142476 4780
rect 142436 4684 142488 4690
rect 142436 4626 142488 4632
rect 142632 3738 142660 4780
rect 143080 4616 143132 4622
rect 143080 4558 143132 4564
rect 143092 4321 143120 4558
rect 143078 4312 143134 4321
rect 143078 4247 143134 4256
rect 142896 4140 142948 4146
rect 142896 4082 142948 4088
rect 142344 3732 142396 3738
rect 142344 3674 142396 3680
rect 142620 3732 142672 3738
rect 142620 3674 142672 3680
rect 142632 3194 142660 3674
rect 142908 3194 142936 4082
rect 142988 3392 143040 3398
rect 142988 3334 143040 3340
rect 141976 3188 142028 3194
rect 141976 3130 142028 3136
rect 142620 3188 142672 3194
rect 142620 3130 142672 3136
rect 142896 3188 142948 3194
rect 142896 3130 142948 3136
rect 141804 2746 141924 2774
rect 141804 2428 141832 2746
rect 141988 2514 142016 3130
rect 142632 2774 142660 3130
rect 143000 3126 143028 3334
rect 142988 3120 143040 3126
rect 142988 3062 143040 3068
rect 143184 2774 143212 10950
rect 143368 8634 143396 12854
rect 143736 11778 143764 15200
rect 143998 14240 144054 14249
rect 143998 14175 144054 14184
rect 143906 14104 143962 14113
rect 143906 14039 143962 14048
rect 143816 13184 143868 13190
rect 143816 13126 143868 13132
rect 143828 11898 143856 13126
rect 143920 12714 143948 14039
rect 144012 13258 144040 14175
rect 144000 13252 144052 13258
rect 144000 13194 144052 13200
rect 144288 13025 144316 15200
rect 144274 13016 144330 13025
rect 144274 12951 144330 12960
rect 143908 12708 143960 12714
rect 143908 12650 143960 12656
rect 144736 12640 144788 12646
rect 144736 12582 144788 12588
rect 144182 12336 144238 12345
rect 144182 12271 144238 12280
rect 143816 11892 143868 11898
rect 143816 11834 143868 11840
rect 143908 11892 143960 11898
rect 143908 11834 143960 11840
rect 143920 11778 143948 11834
rect 143736 11750 143948 11778
rect 144196 11762 144224 12271
rect 144748 12238 144776 12582
rect 144840 12238 144868 15200
rect 145392 13802 145420 15200
rect 145944 15026 145972 15200
rect 146496 15094 146524 15200
rect 146484 15088 146536 15094
rect 146484 15030 146536 15036
rect 145932 15020 145984 15026
rect 145932 14962 145984 14968
rect 146024 14816 146076 14822
rect 146024 14758 146076 14764
rect 145380 13796 145432 13802
rect 145380 13738 145432 13744
rect 145654 13288 145710 13297
rect 145654 13223 145710 13232
rect 145840 13252 145892 13258
rect 145104 13184 145156 13190
rect 145104 13126 145156 13132
rect 145116 12617 145144 13126
rect 145564 12640 145616 12646
rect 145102 12608 145158 12617
rect 145564 12582 145616 12588
rect 145102 12543 145158 12552
rect 144736 12232 144788 12238
rect 144736 12174 144788 12180
rect 144828 12232 144880 12238
rect 144828 12174 144880 12180
rect 144276 12164 144328 12170
rect 144276 12106 144328 12112
rect 144184 11756 144236 11762
rect 144184 11698 144236 11704
rect 143816 11280 143868 11286
rect 143816 11222 143868 11228
rect 143446 11112 143502 11121
rect 143446 11047 143502 11056
rect 143460 11014 143488 11047
rect 143448 11008 143500 11014
rect 143448 10950 143500 10956
rect 143540 10532 143592 10538
rect 143540 10474 143592 10480
rect 143448 10056 143500 10062
rect 143448 9998 143500 10004
rect 143460 9586 143488 9998
rect 143552 9722 143580 10474
rect 143540 9716 143592 9722
rect 143540 9658 143592 9664
rect 143448 9580 143500 9586
rect 143448 9522 143500 9528
rect 143540 9580 143592 9586
rect 143540 9522 143592 9528
rect 143448 9104 143500 9110
rect 143552 9058 143580 9522
rect 143724 9376 143776 9382
rect 143722 9344 143724 9353
rect 143776 9344 143778 9353
rect 143722 9279 143778 9288
rect 143500 9052 143580 9058
rect 143448 9046 143580 9052
rect 143460 9030 143580 9046
rect 143632 8968 143684 8974
rect 143632 8910 143684 8916
rect 143356 8628 143408 8634
rect 143356 8570 143408 8576
rect 143264 8492 143316 8498
rect 143264 8434 143316 8440
rect 143276 7342 143304 8434
rect 143264 7336 143316 7342
rect 143264 7278 143316 7284
rect 143448 7336 143500 7342
rect 143448 7278 143500 7284
rect 143460 6798 143488 7278
rect 143448 6792 143500 6798
rect 143448 6734 143500 6740
rect 143356 6452 143408 6458
rect 143356 6394 143408 6400
rect 143368 5642 143396 6394
rect 143356 5636 143408 5642
rect 143356 5578 143408 5584
rect 143356 4616 143408 4622
rect 143356 4558 143408 4564
rect 143368 4214 143396 4558
rect 143644 4321 143672 8910
rect 143736 8809 143764 9279
rect 143722 8800 143778 8809
rect 143722 8735 143778 8744
rect 143828 7993 143856 11222
rect 144000 11076 144052 11082
rect 144000 11018 144052 11024
rect 144012 9761 144040 11018
rect 144184 10668 144236 10674
rect 144184 10610 144236 10616
rect 144092 9920 144144 9926
rect 144092 9862 144144 9868
rect 143998 9752 144054 9761
rect 143908 9716 143960 9722
rect 143998 9687 144054 9696
rect 143908 9658 143960 9664
rect 143920 8498 143948 9658
rect 144104 8809 144132 9862
rect 144090 8800 144146 8809
rect 144090 8735 144146 8744
rect 143908 8492 143960 8498
rect 143908 8434 143960 8440
rect 143814 7984 143870 7993
rect 143814 7919 143870 7928
rect 144000 7472 144052 7478
rect 144000 7414 144052 7420
rect 143736 6458 143948 6474
rect 143736 6452 143960 6458
rect 143736 6446 143908 6452
rect 143736 6390 143764 6446
rect 143908 6394 143960 6400
rect 143724 6384 143776 6390
rect 143816 6384 143868 6390
rect 143724 6326 143776 6332
rect 143814 6352 143816 6361
rect 143868 6352 143870 6361
rect 143814 6287 143870 6296
rect 143816 4820 143868 4826
rect 143816 4762 143868 4768
rect 143630 4312 143686 4321
rect 143630 4247 143686 4256
rect 143356 4208 143408 4214
rect 143356 4150 143408 4156
rect 143632 3936 143684 3942
rect 143632 3878 143684 3884
rect 143644 3641 143672 3878
rect 143630 3632 143686 3641
rect 143630 3567 143686 3576
rect 143632 3528 143684 3534
rect 143632 3470 143684 3476
rect 143724 3528 143776 3534
rect 143724 3470 143776 3476
rect 142540 2746 142660 2774
rect 142816 2746 143212 2774
rect 142540 2650 142568 2746
rect 142528 2644 142580 2650
rect 142528 2586 142580 2592
rect 141976 2508 142028 2514
rect 141976 2450 142028 2456
rect 141884 2440 141936 2446
rect 141804 2400 141884 2428
rect 141884 2382 141936 2388
rect 141700 2372 141752 2378
rect 141700 2314 141752 2320
rect 141976 2372 142028 2378
rect 141976 2314 142028 2320
rect 140596 2246 140648 2252
rect 141054 2272 141110 2281
rect 140608 1766 140636 2246
rect 141054 2207 141110 2216
rect 141988 1834 142016 2314
rect 141976 1828 142028 1834
rect 141976 1770 142028 1776
rect 140596 1760 140648 1766
rect 140596 1702 140648 1708
rect 142816 1698 142844 2746
rect 143644 1766 143672 3470
rect 143736 3398 143764 3470
rect 143724 3392 143776 3398
rect 143724 3334 143776 3340
rect 143828 2990 143856 4762
rect 143816 2984 143868 2990
rect 143816 2926 143868 2932
rect 143724 2576 143776 2582
rect 143722 2544 143724 2553
rect 143776 2544 143778 2553
rect 143722 2479 143778 2488
rect 143736 1873 143764 2479
rect 143722 1864 143778 1873
rect 143722 1799 143778 1808
rect 143632 1760 143684 1766
rect 143632 1702 143684 1708
rect 142804 1692 142856 1698
rect 142804 1634 142856 1640
rect 144012 1630 144040 7414
rect 144196 6905 144224 10610
rect 144288 9926 144316 12106
rect 144460 11756 144512 11762
rect 144460 11698 144512 11704
rect 144368 10192 144420 10198
rect 144368 10134 144420 10140
rect 144276 9920 144328 9926
rect 144276 9862 144328 9868
rect 144380 9586 144408 10134
rect 144368 9580 144420 9586
rect 144368 9522 144420 9528
rect 144472 8294 144500 11698
rect 144642 11248 144698 11257
rect 144642 11183 144698 11192
rect 144552 11076 144604 11082
rect 144552 11018 144604 11024
rect 144564 8838 144592 11018
rect 144656 9994 144684 11183
rect 144748 11098 144776 12174
rect 145012 12096 145064 12102
rect 145012 12038 145064 12044
rect 145024 11937 145052 12038
rect 145010 11928 145066 11937
rect 145010 11863 145066 11872
rect 144828 11756 144880 11762
rect 144828 11698 144880 11704
rect 144840 11218 144868 11698
rect 144920 11552 144972 11558
rect 144920 11494 144972 11500
rect 144932 11218 144960 11494
rect 145286 11384 145342 11393
rect 145286 11319 145342 11328
rect 144828 11212 144880 11218
rect 144828 11154 144880 11160
rect 144920 11212 144972 11218
rect 144920 11154 144972 11160
rect 144748 11070 144868 11098
rect 144734 10840 144790 10849
rect 144734 10775 144790 10784
rect 144748 10674 144776 10775
rect 144736 10668 144788 10674
rect 144736 10610 144788 10616
rect 144644 9988 144696 9994
rect 144644 9930 144696 9936
rect 144840 9926 144868 11070
rect 145300 11014 145328 11319
rect 145288 11008 145340 11014
rect 145288 10950 145340 10956
rect 145380 11008 145432 11014
rect 145380 10950 145432 10956
rect 144920 10736 144972 10742
rect 144920 10678 144972 10684
rect 144932 10198 144960 10678
rect 145196 10668 145248 10674
rect 145196 10610 145248 10616
rect 144920 10192 144972 10198
rect 144920 10134 144972 10140
rect 145208 10130 145236 10610
rect 145196 10124 145248 10130
rect 145196 10066 145248 10072
rect 144920 10056 144972 10062
rect 144920 9998 144972 10004
rect 144736 9920 144788 9926
rect 144736 9862 144788 9868
rect 144828 9920 144880 9926
rect 144828 9862 144880 9868
rect 144642 9752 144698 9761
rect 144642 9687 144698 9696
rect 144656 9110 144684 9687
rect 144644 9104 144696 9110
rect 144644 9046 144696 9052
rect 144644 8968 144696 8974
rect 144644 8910 144696 8916
rect 144552 8832 144604 8838
rect 144552 8774 144604 8780
rect 144472 8266 144592 8294
rect 144368 7880 144420 7886
rect 144368 7822 144420 7828
rect 144380 7410 144408 7822
rect 144368 7404 144420 7410
rect 144368 7346 144420 7352
rect 144182 6896 144238 6905
rect 144182 6831 144238 6840
rect 144092 6316 144144 6322
rect 144092 6258 144144 6264
rect 144104 5778 144132 6258
rect 144196 5846 144224 6831
rect 144564 6361 144592 8266
rect 144656 7834 144684 8910
rect 144748 8090 144776 9862
rect 144840 8974 144868 9862
rect 144932 9761 144960 9998
rect 144918 9752 144974 9761
rect 144918 9687 144974 9696
rect 145012 9580 145064 9586
rect 145012 9522 145064 9528
rect 145024 8974 145052 9522
rect 145208 9518 145236 10066
rect 145196 9512 145248 9518
rect 145196 9454 145248 9460
rect 145104 9104 145156 9110
rect 145104 9046 145156 9052
rect 144828 8968 144880 8974
rect 144828 8910 144880 8916
rect 145012 8968 145064 8974
rect 145012 8910 145064 8916
rect 144826 8664 144882 8673
rect 144826 8599 144882 8608
rect 144920 8628 144972 8634
rect 144840 8514 144868 8599
rect 144972 8588 145052 8616
rect 144920 8570 144972 8576
rect 144840 8486 144960 8514
rect 144932 8430 144960 8486
rect 144920 8424 144972 8430
rect 144920 8366 144972 8372
rect 144920 8288 144972 8294
rect 144920 8230 144972 8236
rect 144736 8084 144788 8090
rect 144736 8026 144788 8032
rect 144656 7806 144868 7834
rect 144644 7744 144696 7750
rect 144644 7686 144696 7692
rect 144550 6352 144606 6361
rect 144550 6287 144606 6296
rect 144184 5840 144236 5846
rect 144184 5782 144236 5788
rect 144092 5772 144144 5778
rect 144092 5714 144144 5720
rect 144656 5370 144684 7686
rect 144840 7041 144868 7806
rect 144932 7721 144960 8230
rect 144918 7712 144974 7721
rect 144918 7647 144974 7656
rect 145024 7342 145052 8588
rect 145012 7336 145064 7342
rect 145012 7278 145064 7284
rect 144826 7032 144882 7041
rect 144826 6967 144882 6976
rect 145010 7032 145066 7041
rect 145010 6967 145066 6976
rect 144840 6338 144868 6967
rect 145024 6458 145052 6967
rect 145012 6452 145064 6458
rect 145012 6394 145064 6400
rect 144840 6322 144960 6338
rect 144736 6316 144788 6322
rect 144840 6316 144972 6322
rect 144840 6310 144920 6316
rect 144736 6258 144788 6264
rect 144920 6258 144972 6264
rect 144748 6202 144776 6258
rect 144748 6174 145052 6202
rect 144920 5908 144972 5914
rect 145024 5896 145052 6174
rect 144972 5868 145052 5896
rect 144920 5850 144972 5856
rect 144644 5364 144696 5370
rect 144644 5306 144696 5312
rect 144184 5296 144236 5302
rect 144184 5238 144236 5244
rect 144196 4622 144224 5238
rect 144184 4616 144236 4622
rect 144184 4558 144236 4564
rect 144276 4616 144328 4622
rect 144276 4558 144328 4564
rect 144184 4140 144236 4146
rect 144288 4128 144316 4558
rect 144236 4100 144316 4128
rect 144734 4176 144790 4185
rect 144918 4176 144974 4185
rect 144790 4134 144918 4162
rect 144734 4111 144790 4120
rect 144918 4111 144974 4120
rect 144184 4082 144236 4088
rect 144196 3602 144224 4082
rect 144184 3596 144236 3602
rect 144184 3538 144236 3544
rect 144196 2650 144224 3538
rect 145024 3466 145052 5868
rect 145012 3460 145064 3466
rect 145012 3402 145064 3408
rect 145116 2774 145144 9046
rect 145300 8945 145328 10950
rect 145286 8936 145342 8945
rect 145286 8871 145342 8880
rect 145196 8016 145248 8022
rect 145196 7958 145248 7964
rect 145208 6882 145236 7958
rect 145288 7472 145340 7478
rect 145288 7414 145340 7420
rect 145300 7041 145328 7414
rect 145392 7274 145420 10950
rect 145472 9920 145524 9926
rect 145472 9862 145524 9868
rect 145484 9654 145512 9862
rect 145472 9648 145524 9654
rect 145576 9625 145604 12582
rect 145668 11558 145696 13223
rect 145840 13194 145892 13200
rect 145852 13161 145880 13194
rect 145838 13152 145894 13161
rect 145838 13087 145894 13096
rect 145840 12776 145892 12782
rect 145840 12718 145892 12724
rect 145852 11665 145880 12718
rect 145838 11656 145894 11665
rect 145838 11591 145894 11600
rect 145656 11552 145708 11558
rect 145656 11494 145708 11500
rect 146036 10062 146064 14758
rect 146206 13968 146262 13977
rect 146206 13903 146262 13912
rect 146220 13734 146248 13903
rect 146944 13864 146996 13870
rect 146944 13806 146996 13812
rect 146208 13728 146260 13734
rect 146208 13670 146260 13676
rect 146220 13258 146248 13670
rect 146956 13394 146984 13806
rect 147048 13705 147076 15200
rect 147034 13696 147090 13705
rect 147034 13631 147090 13640
rect 147600 13569 147628 15200
rect 148428 13938 148456 15286
rect 148690 15200 148746 16000
rect 149242 15200 149298 16000
rect 149794 15314 149850 16000
rect 150346 15314 150402 16000
rect 149794 15286 150112 15314
rect 149794 15200 149850 15286
rect 148416 13932 148468 13938
rect 148416 13874 148468 13880
rect 147586 13560 147642 13569
rect 147586 13495 147642 13504
rect 148048 13524 148100 13530
rect 148048 13466 148100 13472
rect 148600 13524 148652 13530
rect 148600 13466 148652 13472
rect 147404 13456 147456 13462
rect 148060 13433 148088 13466
rect 148140 13456 148192 13462
rect 147404 13398 147456 13404
rect 148046 13424 148102 13433
rect 146944 13388 146996 13394
rect 146944 13330 146996 13336
rect 146208 13252 146260 13258
rect 146208 13194 146260 13200
rect 146484 13252 146536 13258
rect 146484 13194 146536 13200
rect 146300 12980 146352 12986
rect 146300 12922 146352 12928
rect 146312 12753 146340 12922
rect 146298 12744 146354 12753
rect 146298 12679 146354 12688
rect 146496 12434 146524 13194
rect 147036 12640 147088 12646
rect 147036 12582 147088 12588
rect 146312 12406 146524 12434
rect 146116 12164 146168 12170
rect 146116 12106 146168 12112
rect 146024 10056 146076 10062
rect 146024 9998 146076 10004
rect 146128 9994 146156 12106
rect 146208 10124 146260 10130
rect 146208 10066 146260 10072
rect 146116 9988 146168 9994
rect 146116 9930 146168 9936
rect 145472 9590 145524 9596
rect 145562 9616 145618 9625
rect 145562 9551 145618 9560
rect 145656 9512 145708 9518
rect 145656 9454 145708 9460
rect 145564 9376 145616 9382
rect 145564 9318 145616 9324
rect 145472 9104 145524 9110
rect 145472 9046 145524 9052
rect 145380 7268 145432 7274
rect 145380 7210 145432 7216
rect 145286 7032 145342 7041
rect 145286 6967 145342 6976
rect 145208 6854 145420 6882
rect 145288 6724 145340 6730
rect 145288 6666 145340 6672
rect 145194 5944 145250 5953
rect 145300 5914 145328 6666
rect 145194 5879 145250 5888
rect 145288 5908 145340 5914
rect 145208 4146 145236 5879
rect 145288 5850 145340 5856
rect 145286 5536 145342 5545
rect 145286 5471 145342 5480
rect 145300 5234 145328 5471
rect 145288 5228 145340 5234
rect 145288 5170 145340 5176
rect 145300 5030 145328 5170
rect 145288 5024 145340 5030
rect 145288 4966 145340 4972
rect 145288 4752 145340 4758
rect 145288 4694 145340 4700
rect 145196 4140 145248 4146
rect 145196 4082 145248 4088
rect 145300 2990 145328 4694
rect 145392 3670 145420 6854
rect 145380 3664 145432 3670
rect 145380 3606 145432 3612
rect 145484 3126 145512 9046
rect 145576 8945 145604 9318
rect 145562 8936 145618 8945
rect 145562 8871 145618 8880
rect 145668 8498 145696 9454
rect 145748 9376 145800 9382
rect 145748 9318 145800 9324
rect 145760 9178 145788 9318
rect 145748 9172 145800 9178
rect 145748 9114 145800 9120
rect 146024 9172 146076 9178
rect 146024 9114 146076 9120
rect 145840 9036 145892 9042
rect 145840 8978 145892 8984
rect 145656 8492 145708 8498
rect 145656 8434 145708 8440
rect 145564 8424 145616 8430
rect 145564 8366 145616 8372
rect 145576 5370 145604 8366
rect 145852 8129 145880 8978
rect 145932 8832 145984 8838
rect 145932 8774 145984 8780
rect 145838 8120 145894 8129
rect 145838 8055 145894 8064
rect 145748 7812 145800 7818
rect 145748 7754 145800 7760
rect 145654 7576 145710 7585
rect 145654 7511 145710 7520
rect 145668 6458 145696 7511
rect 145656 6452 145708 6458
rect 145656 6394 145708 6400
rect 145656 6316 145708 6322
rect 145656 6258 145708 6264
rect 145668 5953 145696 6258
rect 145654 5944 145710 5953
rect 145654 5879 145710 5888
rect 145564 5364 145616 5370
rect 145564 5306 145616 5312
rect 145668 5250 145696 5879
rect 145576 5222 145696 5250
rect 145576 4758 145604 5222
rect 145656 5024 145708 5030
rect 145656 4966 145708 4972
rect 145564 4752 145616 4758
rect 145564 4694 145616 4700
rect 145564 4480 145616 4486
rect 145562 4448 145564 4457
rect 145616 4448 145618 4457
rect 145562 4383 145618 4392
rect 145562 4312 145618 4321
rect 145562 4247 145618 4256
rect 145576 4214 145604 4247
rect 145564 4208 145616 4214
rect 145668 4185 145696 4966
rect 145564 4150 145616 4156
rect 145654 4176 145710 4185
rect 145654 4111 145710 4120
rect 145564 4004 145616 4010
rect 145564 3946 145616 3952
rect 145472 3120 145524 3126
rect 145470 3088 145472 3097
rect 145524 3088 145526 3097
rect 145576 3058 145604 3946
rect 145470 3023 145526 3032
rect 145564 3052 145616 3058
rect 145564 2994 145616 3000
rect 145288 2984 145340 2990
rect 145288 2926 145340 2932
rect 145656 2984 145708 2990
rect 145656 2926 145708 2932
rect 145024 2746 145144 2774
rect 144184 2644 144236 2650
rect 144184 2586 144236 2592
rect 145024 2009 145052 2746
rect 145668 2514 145696 2926
rect 145656 2508 145708 2514
rect 145656 2450 145708 2456
rect 145010 2000 145066 2009
rect 145010 1935 145066 1944
rect 144000 1624 144052 1630
rect 144000 1566 144052 1572
rect 145760 1057 145788 7754
rect 145838 7576 145894 7585
rect 145838 7511 145894 7520
rect 145852 7177 145880 7511
rect 145944 7274 145972 8774
rect 146036 8634 146064 9114
rect 146220 9081 146248 10066
rect 146206 9072 146262 9081
rect 146206 9007 146262 9016
rect 146024 8628 146076 8634
rect 146024 8570 146076 8576
rect 146024 8288 146076 8294
rect 146024 8230 146076 8236
rect 145932 7268 145984 7274
rect 145932 7210 145984 7216
rect 146036 7206 146064 8230
rect 146312 7750 146340 12406
rect 146392 12232 146444 12238
rect 146392 12174 146444 12180
rect 146404 11830 146432 12174
rect 146392 11824 146444 11830
rect 146392 11766 146444 11772
rect 146404 11234 146432 11766
rect 146944 11756 146996 11762
rect 146944 11698 146996 11704
rect 146404 11206 146616 11234
rect 146588 11150 146616 11206
rect 146576 11144 146628 11150
rect 146576 11086 146628 11092
rect 146852 11144 146904 11150
rect 146852 11086 146904 11092
rect 146588 10588 146616 11086
rect 146668 10600 146720 10606
rect 146588 10560 146668 10588
rect 146668 10542 146720 10548
rect 146864 10554 146892 11086
rect 146956 10674 146984 11698
rect 146944 10668 146996 10674
rect 146944 10610 146996 10616
rect 146680 10266 146708 10542
rect 146864 10526 146984 10554
rect 146852 10464 146904 10470
rect 146852 10406 146904 10412
rect 146668 10260 146720 10266
rect 146668 10202 146720 10208
rect 146760 7948 146812 7954
rect 146760 7890 146812 7896
rect 146392 7880 146444 7886
rect 146392 7822 146444 7828
rect 146300 7744 146352 7750
rect 146300 7686 146352 7692
rect 146208 7540 146260 7546
rect 146208 7482 146260 7488
rect 146024 7200 146076 7206
rect 145838 7168 145894 7177
rect 146024 7142 146076 7148
rect 146116 7200 146168 7206
rect 146116 7142 146168 7148
rect 145838 7103 145894 7112
rect 145932 6316 145984 6322
rect 145932 6258 145984 6264
rect 145944 6186 145972 6258
rect 145932 6180 145984 6186
rect 145932 6122 145984 6128
rect 145932 5160 145984 5166
rect 145932 5102 145984 5108
rect 145840 4752 145892 4758
rect 145840 4694 145892 4700
rect 145852 4622 145880 4694
rect 145840 4616 145892 4622
rect 145840 4558 145892 4564
rect 145944 4321 145972 5102
rect 146022 4856 146078 4865
rect 146022 4791 146024 4800
rect 146076 4791 146078 4800
rect 146024 4762 146076 4768
rect 145930 4312 145986 4321
rect 145930 4247 145986 4256
rect 145932 2372 145984 2378
rect 145932 2314 145984 2320
rect 145944 2281 145972 2314
rect 145930 2272 145986 2281
rect 145930 2207 145986 2216
rect 145944 2106 145972 2207
rect 145932 2100 145984 2106
rect 145932 2042 145984 2048
rect 146128 1902 146156 7142
rect 146220 5794 146248 7482
rect 146404 7410 146432 7822
rect 146392 7404 146444 7410
rect 146392 7346 146444 7352
rect 146404 6798 146432 7346
rect 146576 7336 146628 7342
rect 146576 7278 146628 7284
rect 146484 6928 146536 6934
rect 146484 6870 146536 6876
rect 146392 6792 146444 6798
rect 146392 6734 146444 6740
rect 146300 6724 146352 6730
rect 146300 6666 146352 6672
rect 146312 6458 146340 6666
rect 146300 6452 146352 6458
rect 146300 6394 146352 6400
rect 146404 6118 146432 6734
rect 146496 6633 146524 6870
rect 146588 6798 146616 7278
rect 146576 6792 146628 6798
rect 146576 6734 146628 6740
rect 146772 6633 146800 7890
rect 146482 6624 146538 6633
rect 146482 6559 146538 6568
rect 146758 6624 146814 6633
rect 146758 6559 146814 6568
rect 146392 6112 146444 6118
rect 146392 6054 146444 6060
rect 146220 5766 146616 5794
rect 146392 5704 146444 5710
rect 146312 5664 146392 5692
rect 146208 5636 146260 5642
rect 146208 5578 146260 5584
rect 146220 3913 146248 5578
rect 146312 5001 146340 5664
rect 146392 5646 146444 5652
rect 146298 4992 146354 5001
rect 146298 4927 146354 4936
rect 146482 4992 146538 5001
rect 146482 4927 146538 4936
rect 146206 3904 146262 3913
rect 146206 3839 146262 3848
rect 146298 3768 146354 3777
rect 146298 3703 146300 3712
rect 146352 3703 146354 3712
rect 146300 3674 146352 3680
rect 146208 3392 146260 3398
rect 146208 3334 146260 3340
rect 146116 1896 146168 1902
rect 146116 1838 146168 1844
rect 146220 1698 146248 3334
rect 146496 3194 146524 4927
rect 146588 3398 146616 5766
rect 146772 5710 146800 6559
rect 146864 5794 146892 10406
rect 146956 7478 146984 10526
rect 147048 10470 147076 12582
rect 147310 12336 147366 12345
rect 147310 12271 147366 12280
rect 147128 11688 147180 11694
rect 147128 11630 147180 11636
rect 147140 11354 147168 11630
rect 147324 11354 147352 12271
rect 147416 11540 147444 13398
rect 148140 13398 148192 13404
rect 148046 13359 148102 13368
rect 147496 13320 147548 13326
rect 147496 13262 147548 13268
rect 147508 12850 147536 13262
rect 147496 12844 147548 12850
rect 147496 12786 147548 12792
rect 148152 12442 148180 13398
rect 148612 13258 148640 13466
rect 148600 13252 148652 13258
rect 148600 13194 148652 13200
rect 148508 12912 148560 12918
rect 148508 12854 148560 12860
rect 148140 12436 148192 12442
rect 148140 12378 148192 12384
rect 148416 12300 148468 12306
rect 148416 12242 148468 12248
rect 148048 12232 148100 12238
rect 148048 12174 148100 12180
rect 148232 12232 148284 12238
rect 148232 12174 148284 12180
rect 147680 12164 147732 12170
rect 147680 12106 147732 12112
rect 147588 12096 147640 12102
rect 147588 12038 147640 12044
rect 147600 11830 147628 12038
rect 147588 11824 147640 11830
rect 147588 11766 147640 11772
rect 147496 11688 147548 11694
rect 147548 11636 147628 11642
rect 147496 11630 147628 11636
rect 147508 11614 147628 11630
rect 147600 11558 147628 11614
rect 147496 11552 147548 11558
rect 147416 11512 147496 11540
rect 147496 11494 147548 11500
rect 147588 11552 147640 11558
rect 147588 11494 147640 11500
rect 147508 11354 147536 11494
rect 147692 11393 147720 12106
rect 148060 11393 148088 12174
rect 148244 11642 148272 12174
rect 148428 12102 148456 12242
rect 148324 12096 148376 12102
rect 148324 12038 148376 12044
rect 148416 12096 148468 12102
rect 148416 12038 148468 12044
rect 148336 11898 148364 12038
rect 148520 11937 148548 12854
rect 148600 12232 148652 12238
rect 148600 12174 148652 12180
rect 148506 11928 148562 11937
rect 148324 11892 148376 11898
rect 148506 11863 148562 11872
rect 148324 11834 148376 11840
rect 148324 11756 148376 11762
rect 148376 11716 148456 11744
rect 148324 11698 148376 11704
rect 148244 11614 148364 11642
rect 148140 11552 148192 11558
rect 148140 11494 148192 11500
rect 147678 11384 147734 11393
rect 147128 11348 147180 11354
rect 147312 11348 147364 11354
rect 147128 11290 147180 11296
rect 147232 11308 147312 11336
rect 147036 10464 147088 10470
rect 147036 10406 147088 10412
rect 147036 10260 147088 10266
rect 147088 10220 147168 10248
rect 147036 10202 147088 10208
rect 147036 10056 147088 10062
rect 147036 9998 147088 10004
rect 147048 7954 147076 9998
rect 147140 9518 147168 10220
rect 147232 10062 147260 11308
rect 147312 11290 147364 11296
rect 147496 11348 147548 11354
rect 148046 11384 148102 11393
rect 147678 11319 147734 11328
rect 147772 11348 147824 11354
rect 147496 11290 147548 11296
rect 148046 11319 148102 11328
rect 147772 11290 147824 11296
rect 147784 11121 147812 11290
rect 147770 11112 147826 11121
rect 147770 11047 147826 11056
rect 147312 10804 147364 10810
rect 147312 10746 147364 10752
rect 147324 10198 147352 10746
rect 147416 10390 147904 10418
rect 147312 10192 147364 10198
rect 147312 10134 147364 10140
rect 147220 10056 147272 10062
rect 147220 9998 147272 10004
rect 147416 9722 147444 10390
rect 147876 10266 147904 10390
rect 147772 10260 147824 10266
rect 147772 10202 147824 10208
rect 147864 10260 147916 10266
rect 147864 10202 147916 10208
rect 147784 10146 147812 10202
rect 147784 10118 147904 10146
rect 147876 9926 147904 10118
rect 148048 10056 148100 10062
rect 148048 9998 148100 10004
rect 147864 9920 147916 9926
rect 147864 9862 147916 9868
rect 147404 9716 147456 9722
rect 147404 9658 147456 9664
rect 147956 9716 148008 9722
rect 147956 9658 148008 9664
rect 147312 9580 147364 9586
rect 147312 9522 147364 9528
rect 147128 9512 147180 9518
rect 147128 9454 147180 9460
rect 147140 9042 147168 9454
rect 147220 9104 147272 9110
rect 147220 9046 147272 9052
rect 147128 9036 147180 9042
rect 147128 8978 147180 8984
rect 147128 8900 147180 8906
rect 147128 8842 147180 8848
rect 147140 8430 147168 8842
rect 147128 8424 147180 8430
rect 147128 8366 147180 8372
rect 147232 8362 147260 9046
rect 147220 8356 147272 8362
rect 147220 8298 147272 8304
rect 147218 8120 147274 8129
rect 147218 8055 147274 8064
rect 147232 8022 147260 8055
rect 147220 8016 147272 8022
rect 147220 7958 147272 7964
rect 147324 7970 147352 9522
rect 147496 9036 147548 9042
rect 147496 8978 147548 8984
rect 147404 8968 147456 8974
rect 147402 8936 147404 8945
rect 147456 8936 147458 8945
rect 147402 8871 147458 8880
rect 147508 8838 147536 8978
rect 147770 8936 147826 8945
rect 147770 8871 147826 8880
rect 147496 8832 147548 8838
rect 147496 8774 147548 8780
rect 147784 8634 147812 8871
rect 147772 8628 147824 8634
rect 147772 8570 147824 8576
rect 147404 8492 147456 8498
rect 147456 8452 147536 8480
rect 147404 8434 147456 8440
rect 147508 8378 147536 8452
rect 147404 8356 147456 8362
rect 147508 8350 147904 8378
rect 147404 8298 147456 8304
rect 147416 8072 147444 8298
rect 147416 8044 147812 8072
rect 147036 7948 147088 7954
rect 147324 7942 147628 7970
rect 147036 7890 147088 7896
rect 147312 7880 147364 7886
rect 147364 7840 147536 7868
rect 147312 7822 147364 7828
rect 147128 7812 147180 7818
rect 147128 7754 147180 7760
rect 146944 7472 146996 7478
rect 146944 7414 146996 7420
rect 147140 7256 147168 7754
rect 147048 7228 147168 7256
rect 147048 7002 147076 7228
rect 147126 7168 147182 7177
rect 147126 7103 147182 7112
rect 147036 6996 147088 7002
rect 147036 6938 147088 6944
rect 146942 6488 146998 6497
rect 146942 6423 146998 6432
rect 146956 6322 146984 6423
rect 147140 6322 147168 7103
rect 147312 6656 147364 6662
rect 147312 6598 147364 6604
rect 147324 6474 147352 6598
rect 147232 6446 147352 6474
rect 146944 6316 146996 6322
rect 146944 6258 146996 6264
rect 147128 6316 147180 6322
rect 147128 6258 147180 6264
rect 147036 6248 147088 6254
rect 147036 6190 147088 6196
rect 147048 5953 147076 6190
rect 147034 5944 147090 5953
rect 147034 5879 147090 5888
rect 146864 5766 147168 5794
rect 146760 5704 146812 5710
rect 146944 5704 146996 5710
rect 146760 5646 146812 5652
rect 146942 5672 146944 5681
rect 147036 5704 147088 5710
rect 146996 5672 146998 5681
rect 147036 5646 147088 5652
rect 146942 5607 146998 5616
rect 146668 5568 146720 5574
rect 146668 5510 146720 5516
rect 146680 4214 146708 5510
rect 146760 5364 146812 5370
rect 146760 5306 146812 5312
rect 146772 4486 146800 5306
rect 147048 5234 147076 5646
rect 146944 5228 146996 5234
rect 146944 5170 146996 5176
rect 147036 5228 147088 5234
rect 147036 5170 147088 5176
rect 146956 5137 146984 5170
rect 146942 5128 146998 5137
rect 147140 5098 147168 5766
rect 146942 5063 146998 5072
rect 147128 5092 147180 5098
rect 147128 5034 147180 5040
rect 146760 4480 146812 4486
rect 146944 4480 146996 4486
rect 146760 4422 146812 4428
rect 146942 4448 146944 4457
rect 146996 4448 146998 4457
rect 146942 4383 146998 4392
rect 146668 4208 146720 4214
rect 146668 4150 146720 4156
rect 147034 4176 147090 4185
rect 146680 3942 146708 4150
rect 147232 4146 147260 6446
rect 147404 6112 147456 6118
rect 147508 6100 147536 7840
rect 147600 6662 147628 7942
rect 147678 6896 147734 6905
rect 147678 6831 147734 6840
rect 147692 6798 147720 6831
rect 147680 6792 147732 6798
rect 147680 6734 147732 6740
rect 147784 6662 147812 8044
rect 147876 7274 147904 8350
rect 147968 7886 147996 9658
rect 148060 8265 148088 9998
rect 148152 9081 148180 11494
rect 148232 11076 148284 11082
rect 148232 11018 148284 11024
rect 148138 9072 148194 9081
rect 148244 9042 148272 11018
rect 148336 10849 148364 11614
rect 148428 11150 148456 11716
rect 148508 11552 148560 11558
rect 148508 11494 148560 11500
rect 148416 11144 148468 11150
rect 148416 11086 148468 11092
rect 148322 10840 148378 10849
rect 148322 10775 148378 10784
rect 148138 9007 148194 9016
rect 148232 9036 148284 9042
rect 148232 8978 148284 8984
rect 148336 8922 148364 10775
rect 148152 8894 148364 8922
rect 148152 8650 148180 8894
rect 148428 8888 148456 11086
rect 148520 8956 148548 11494
rect 148612 10130 148640 12174
rect 148704 11898 148732 15200
rect 149256 13734 149284 15200
rect 149336 14952 149388 14958
rect 149336 14894 149388 14900
rect 149244 13728 149296 13734
rect 149244 13670 149296 13676
rect 149244 13388 149296 13394
rect 149244 13330 149296 13336
rect 149256 13258 149284 13330
rect 149244 13252 149296 13258
rect 149244 13194 149296 13200
rect 149152 13184 149204 13190
rect 149152 13126 149204 13132
rect 148782 13016 148838 13025
rect 148782 12951 148838 12960
rect 148796 12918 148824 12951
rect 148784 12912 148836 12918
rect 148784 12854 148836 12860
rect 148876 12844 148928 12850
rect 148876 12786 148928 12792
rect 148888 12084 148916 12786
rect 149164 12714 149192 13126
rect 149152 12708 149204 12714
rect 149152 12650 149204 12656
rect 149244 12096 149296 12102
rect 148888 12056 149244 12084
rect 149244 12038 149296 12044
rect 148692 11892 148744 11898
rect 148692 11834 148744 11840
rect 149242 11656 149298 11665
rect 149242 11591 149298 11600
rect 148782 10840 148838 10849
rect 148782 10775 148784 10784
rect 148836 10775 148838 10784
rect 148784 10746 148836 10752
rect 148600 10124 148652 10130
rect 148600 10066 148652 10072
rect 148598 9888 148654 9897
rect 148598 9823 148654 9832
rect 148612 9110 148640 9823
rect 148796 9674 148824 10746
rect 149060 10464 149112 10470
rect 149060 10406 149112 10412
rect 148796 9646 148916 9674
rect 148888 9568 148916 9646
rect 148888 9540 149008 9568
rect 148690 9480 148746 9489
rect 148690 9415 148746 9424
rect 148874 9480 148930 9489
rect 148874 9415 148930 9424
rect 148600 9104 148652 9110
rect 148600 9046 148652 9052
rect 148520 8928 148640 8956
rect 148704 8945 148732 9415
rect 148888 9382 148916 9415
rect 148876 9376 148928 9382
rect 148876 9318 148928 9324
rect 148782 9208 148838 9217
rect 148782 9143 148784 9152
rect 148836 9143 148838 9152
rect 148784 9114 148836 9120
rect 148876 9104 148928 9110
rect 148876 9046 148928 9052
rect 148612 8888 148640 8928
rect 148690 8936 148746 8945
rect 148428 8860 148517 8888
rect 148612 8860 148649 8888
rect 148690 8871 148746 8880
rect 148324 8832 148376 8838
rect 148376 8792 148456 8820
rect 148324 8774 148376 8780
rect 148152 8622 148364 8650
rect 148336 8566 148364 8622
rect 148232 8560 148284 8566
rect 148232 8502 148284 8508
rect 148324 8560 148376 8566
rect 148324 8502 148376 8508
rect 148046 8256 148102 8265
rect 148046 8191 148102 8200
rect 148140 8016 148192 8022
rect 148140 7958 148192 7964
rect 147956 7880 148008 7886
rect 147956 7822 148008 7828
rect 148152 7750 148180 7958
rect 148244 7886 148272 8502
rect 148232 7880 148284 7886
rect 148232 7822 148284 7828
rect 148324 7812 148376 7818
rect 148324 7754 148376 7760
rect 148140 7744 148192 7750
rect 148140 7686 148192 7692
rect 148336 7546 148364 7754
rect 148324 7540 148376 7546
rect 148324 7482 148376 7488
rect 148140 7472 148192 7478
rect 148192 7432 148272 7460
rect 148140 7414 148192 7420
rect 147864 7268 147916 7274
rect 147864 7210 147916 7216
rect 148140 7200 148192 7206
rect 148046 7168 148102 7177
rect 148140 7142 148192 7148
rect 148046 7103 148102 7112
rect 147588 6656 147640 6662
rect 147588 6598 147640 6604
rect 147772 6656 147824 6662
rect 147772 6598 147824 6604
rect 147588 6452 147640 6458
rect 147588 6394 147640 6400
rect 147600 6202 147628 6394
rect 147864 6384 147916 6390
rect 147864 6326 147916 6332
rect 147876 6225 147904 6326
rect 147862 6216 147918 6225
rect 147600 6174 147812 6202
rect 147784 6118 147812 6174
rect 147862 6151 147918 6160
rect 147772 6112 147824 6118
rect 147508 6072 147628 6100
rect 147404 6054 147456 6060
rect 147416 5710 147444 6054
rect 147404 5704 147456 5710
rect 147310 5672 147366 5681
rect 147456 5664 147536 5692
rect 147404 5646 147456 5652
rect 147310 5607 147366 5616
rect 147324 5302 147352 5607
rect 147404 5568 147456 5574
rect 147404 5510 147456 5516
rect 147312 5296 147364 5302
rect 147312 5238 147364 5244
rect 147310 5128 147366 5137
rect 147310 5063 147366 5072
rect 147324 5030 147352 5063
rect 147312 5024 147364 5030
rect 147312 4966 147364 4972
rect 147034 4111 147090 4120
rect 147220 4140 147272 4146
rect 146944 4004 146996 4010
rect 146944 3946 146996 3952
rect 146668 3936 146720 3942
rect 146668 3878 146720 3884
rect 146956 3641 146984 3946
rect 146942 3632 146998 3641
rect 146942 3567 146998 3576
rect 146576 3392 146628 3398
rect 146576 3334 146628 3340
rect 147048 3194 147076 4111
rect 147220 4082 147272 4088
rect 147312 3460 147364 3466
rect 147312 3402 147364 3408
rect 147324 3369 147352 3402
rect 147310 3360 147366 3369
rect 147310 3295 147366 3304
rect 146484 3188 146536 3194
rect 146484 3130 146536 3136
rect 147036 3188 147088 3194
rect 147036 3130 147088 3136
rect 146944 2848 146996 2854
rect 146944 2790 146996 2796
rect 146956 2514 146984 2790
rect 146944 2508 146996 2514
rect 146944 2450 146996 2456
rect 147416 2428 147444 5510
rect 147508 4690 147536 5664
rect 147600 5370 147628 6072
rect 147772 6054 147824 6060
rect 147680 5908 147732 5914
rect 148060 5896 148088 7103
rect 148152 6934 148180 7142
rect 148140 6928 148192 6934
rect 148140 6870 148192 6876
rect 148244 6610 148272 7432
rect 147732 5868 148088 5896
rect 148152 6582 148272 6610
rect 147680 5850 147732 5856
rect 147588 5364 147640 5370
rect 147588 5306 147640 5312
rect 147680 5296 147732 5302
rect 147680 5238 147732 5244
rect 147496 4684 147548 4690
rect 147496 4626 147548 4632
rect 147692 4622 147720 5238
rect 147680 4616 147732 4622
rect 147680 4558 147732 4564
rect 147954 4312 148010 4321
rect 147692 4270 147954 4298
rect 147692 4162 147720 4270
rect 147954 4247 148010 4256
rect 147508 4134 147720 4162
rect 147508 3641 147536 4134
rect 148048 4072 148100 4078
rect 148048 4014 148100 4020
rect 147680 3936 147732 3942
rect 147680 3878 147732 3884
rect 147864 3936 147916 3942
rect 147864 3878 147916 3884
rect 147692 3641 147720 3878
rect 147494 3632 147550 3641
rect 147494 3567 147550 3576
rect 147678 3632 147734 3641
rect 147678 3567 147734 3576
rect 147680 3528 147732 3534
rect 147680 3470 147732 3476
rect 147588 3460 147640 3466
rect 147588 3402 147640 3408
rect 147600 3126 147628 3402
rect 147692 3194 147720 3470
rect 147876 3369 147904 3878
rect 148060 3534 148088 4014
rect 148048 3528 148100 3534
rect 148048 3470 148100 3476
rect 147862 3360 147918 3369
rect 147862 3295 147918 3304
rect 147680 3188 147732 3194
rect 147680 3130 147732 3136
rect 147588 3120 147640 3126
rect 147864 3120 147916 3126
rect 147588 3062 147640 3068
rect 147862 3088 147864 3097
rect 147916 3088 147918 3097
rect 147862 3023 147918 3032
rect 148060 2514 148088 3470
rect 148048 2508 148100 2514
rect 148048 2450 148100 2456
rect 147680 2440 147732 2446
rect 147416 2400 147680 2428
rect 147680 2382 147732 2388
rect 147496 2304 147548 2310
rect 147496 2246 147548 2252
rect 147864 2304 147916 2310
rect 147864 2246 147916 2252
rect 146668 2100 146720 2106
rect 146668 2042 146720 2048
rect 146680 1902 146708 2042
rect 147508 1970 147536 2246
rect 147496 1964 147548 1970
rect 147496 1906 147548 1912
rect 146668 1896 146720 1902
rect 146668 1838 146720 1844
rect 147876 1834 147904 2246
rect 148152 2009 148180 6582
rect 148232 6452 148284 6458
rect 148232 6394 148284 6400
rect 148244 5930 148272 6394
rect 148322 5944 148378 5953
rect 148244 5902 148322 5930
rect 148244 5273 148272 5902
rect 148322 5879 148378 5888
rect 148324 5568 148376 5574
rect 148428 5556 148456 8792
rect 148489 8650 148517 8860
rect 148621 8650 148649 8860
rect 148782 8800 148838 8809
rect 148782 8735 148838 8744
rect 148489 8622 148548 8650
rect 148520 7324 148548 8622
rect 148612 8622 148649 8650
rect 148612 7478 148640 8622
rect 148692 8560 148744 8566
rect 148692 8502 148744 8508
rect 148600 7472 148652 7478
rect 148600 7414 148652 7420
rect 148520 7296 148640 7324
rect 148508 6860 148560 6866
rect 148508 6802 148560 6808
rect 148520 6254 148548 6802
rect 148508 6248 148560 6254
rect 148508 6190 148560 6196
rect 148376 5528 148456 5556
rect 148324 5510 148376 5516
rect 148230 5264 148286 5273
rect 148230 5199 148286 5208
rect 148508 3936 148560 3942
rect 148508 3878 148560 3884
rect 148324 3664 148376 3670
rect 148324 3606 148376 3612
rect 148230 3496 148286 3505
rect 148230 3431 148232 3440
rect 148284 3431 148286 3440
rect 148232 3402 148284 3408
rect 148336 3210 148364 3606
rect 148336 3182 148456 3210
rect 148428 2802 148456 3182
rect 148520 2961 148548 3878
rect 148612 3210 148640 7296
rect 148704 3369 148732 8502
rect 148796 6186 148824 8735
rect 148888 7818 148916 9046
rect 148980 8430 149008 9540
rect 149072 8673 149100 10406
rect 149152 9648 149204 9654
rect 149152 9590 149204 9596
rect 149164 9450 149192 9590
rect 149152 9444 149204 9450
rect 149152 9386 149204 9392
rect 149256 9217 149284 11591
rect 149348 11354 149376 14894
rect 149520 14544 149572 14550
rect 149520 14486 149572 14492
rect 149980 14544 150032 14550
rect 149980 14486 150032 14492
rect 149532 12850 149560 14486
rect 149992 13870 150020 14486
rect 150084 13870 150112 15286
rect 150268 15286 150402 15314
rect 149980 13864 150032 13870
rect 149980 13806 150032 13812
rect 150072 13864 150124 13870
rect 150072 13806 150124 13812
rect 149888 13524 149940 13530
rect 149888 13466 149940 13472
rect 149520 12844 149572 12850
rect 149520 12786 149572 12792
rect 149704 12844 149756 12850
rect 149704 12786 149756 12792
rect 149426 11656 149482 11665
rect 149426 11591 149482 11600
rect 149336 11348 149388 11354
rect 149336 11290 149388 11296
rect 149440 11234 149468 11591
rect 149612 11552 149664 11558
rect 149612 11494 149664 11500
rect 149348 11206 149468 11234
rect 149348 11014 149376 11206
rect 149624 11150 149652 11494
rect 149612 11144 149664 11150
rect 149612 11086 149664 11092
rect 149520 11076 149572 11082
rect 149520 11018 149572 11024
rect 149336 11008 149388 11014
rect 149336 10950 149388 10956
rect 149348 10062 149376 10950
rect 149428 10668 149480 10674
rect 149428 10610 149480 10616
rect 149440 10305 149468 10610
rect 149426 10296 149482 10305
rect 149426 10231 149482 10240
rect 149336 10056 149388 10062
rect 149336 9998 149388 10004
rect 149532 9722 149560 11018
rect 149624 10130 149652 11086
rect 149612 10124 149664 10130
rect 149612 10066 149664 10072
rect 149520 9716 149572 9722
rect 149520 9658 149572 9664
rect 149532 9586 149560 9658
rect 149336 9580 149388 9586
rect 149336 9522 149388 9528
rect 149520 9580 149572 9586
rect 149520 9522 149572 9528
rect 149242 9208 149298 9217
rect 149242 9143 149298 9152
rect 149348 9160 149376 9522
rect 149520 9376 149572 9382
rect 149520 9318 149572 9324
rect 149348 9132 149385 9160
rect 149357 9092 149385 9132
rect 149256 9064 149385 9092
rect 149150 8800 149206 8809
rect 149150 8735 149206 8744
rect 149058 8664 149114 8673
rect 149058 8599 149114 8608
rect 148968 8424 149020 8430
rect 148968 8366 149020 8372
rect 149060 8356 149112 8362
rect 149060 8298 149112 8304
rect 149072 8265 149100 8298
rect 149058 8256 149114 8265
rect 149058 8191 149114 8200
rect 149164 8106 149192 8735
rect 149072 8078 149192 8106
rect 148968 7880 149020 7886
rect 148968 7822 149020 7828
rect 148876 7812 148928 7818
rect 148876 7754 148928 7760
rect 148980 7410 149008 7822
rect 148968 7404 149020 7410
rect 148968 7346 149020 7352
rect 148784 6180 148836 6186
rect 148784 6122 148836 6128
rect 148876 5704 148928 5710
rect 148876 5646 148928 5652
rect 148888 5234 148916 5646
rect 148876 5228 148928 5234
rect 148876 5170 148928 5176
rect 148784 4140 148836 4146
rect 148784 4082 148836 4088
rect 148690 3360 148746 3369
rect 148690 3295 148746 3304
rect 148612 3182 148732 3210
rect 148704 2972 148732 3182
rect 148796 3097 148824 4082
rect 148874 3496 148930 3505
rect 148874 3431 148930 3440
rect 148782 3088 148838 3097
rect 148782 3023 148838 3032
rect 148506 2952 148562 2961
rect 148704 2944 148824 2972
rect 148506 2887 148562 2896
rect 148600 2916 148652 2922
rect 148600 2858 148652 2864
rect 148612 2802 148640 2858
rect 148692 2848 148744 2854
rect 148428 2774 148640 2802
rect 148690 2816 148692 2825
rect 148744 2816 148746 2825
rect 148690 2751 148746 2760
rect 148796 2446 148824 2944
rect 148888 2650 148916 3431
rect 148980 2650 149008 7346
rect 149072 4049 149100 8078
rect 149256 8022 149284 9064
rect 149532 8498 149560 9318
rect 149624 8974 149652 10066
rect 149716 9568 149744 12786
rect 149900 10418 149928 13466
rect 150070 13152 150126 13161
rect 150070 13087 150126 13096
rect 150084 12714 150112 13087
rect 150072 12708 150124 12714
rect 150072 12650 150124 12656
rect 150268 12238 150296 15286
rect 150346 15200 150402 15286
rect 154396 15088 154448 15094
rect 154396 15030 154448 15036
rect 154304 15020 154356 15026
rect 154304 14962 154356 14968
rect 150716 14884 150768 14890
rect 150716 14826 150768 14832
rect 150348 12640 150400 12646
rect 150348 12582 150400 12588
rect 150256 12232 150308 12238
rect 150256 12174 150308 12180
rect 150164 11756 150216 11762
rect 150164 11698 150216 11704
rect 150176 11626 150204 11698
rect 150360 11694 150388 12582
rect 150532 12164 150584 12170
rect 150532 12106 150584 12112
rect 150440 11824 150492 11830
rect 150438 11792 150440 11801
rect 150492 11792 150494 11801
rect 150438 11727 150494 11736
rect 150348 11688 150400 11694
rect 150348 11630 150400 11636
rect 150164 11620 150216 11626
rect 150164 11562 150216 11568
rect 149980 11552 150032 11558
rect 149980 11494 150032 11500
rect 149992 11354 150020 11494
rect 149980 11348 150032 11354
rect 149980 11290 150032 11296
rect 150176 10674 150204 11562
rect 150440 11348 150492 11354
rect 150440 11290 150492 11296
rect 150256 10804 150308 10810
rect 150256 10746 150308 10752
rect 150164 10668 150216 10674
rect 150164 10610 150216 10616
rect 149980 10532 150032 10538
rect 150032 10492 150112 10520
rect 149980 10474 150032 10480
rect 149900 10390 150020 10418
rect 149716 9540 149928 9568
rect 149612 8968 149664 8974
rect 149612 8910 149664 8916
rect 149610 8664 149666 8673
rect 149900 8634 149928 9540
rect 149610 8599 149666 8608
rect 149888 8628 149940 8634
rect 149520 8492 149572 8498
rect 149520 8434 149572 8440
rect 149428 8288 149480 8294
rect 149428 8230 149480 8236
rect 149244 8016 149296 8022
rect 149244 7958 149296 7964
rect 149336 7812 149388 7818
rect 149336 7754 149388 7760
rect 149348 7478 149376 7754
rect 149336 7472 149388 7478
rect 149336 7414 149388 7420
rect 149244 7336 149296 7342
rect 149244 7278 149296 7284
rect 149152 6452 149204 6458
rect 149152 6394 149204 6400
rect 149164 6322 149192 6394
rect 149152 6316 149204 6322
rect 149152 6258 149204 6264
rect 149256 6118 149284 7278
rect 149348 6322 149376 7414
rect 149336 6316 149388 6322
rect 149336 6258 149388 6264
rect 149244 6112 149296 6118
rect 149244 6054 149296 6060
rect 149244 5772 149296 5778
rect 149244 5714 149296 5720
rect 149256 4214 149284 5714
rect 149348 5234 149376 6258
rect 149440 5846 149468 8230
rect 149532 7478 149560 8434
rect 149520 7472 149572 7478
rect 149520 7414 149572 7420
rect 149520 6112 149572 6118
rect 149520 6054 149572 6060
rect 149428 5840 149480 5846
rect 149428 5782 149480 5788
rect 149532 5710 149560 6054
rect 149520 5704 149572 5710
rect 149518 5672 149520 5681
rect 149572 5672 149574 5681
rect 149518 5607 149574 5616
rect 149532 5581 149560 5607
rect 149428 5568 149480 5574
rect 149428 5510 149480 5516
rect 149336 5228 149388 5234
rect 149336 5170 149388 5176
rect 149440 4486 149468 5510
rect 149624 4808 149652 8599
rect 149888 8570 149940 8576
rect 149888 8492 149940 8498
rect 149888 8434 149940 8440
rect 149900 8090 149928 8434
rect 149992 8294 150020 10390
rect 150084 10130 150112 10492
rect 150268 10470 150296 10746
rect 150452 10606 150480 11290
rect 150440 10600 150492 10606
rect 150440 10542 150492 10548
rect 150256 10464 150308 10470
rect 150256 10406 150308 10412
rect 150254 10296 150310 10305
rect 150310 10254 150388 10282
rect 150254 10231 150310 10240
rect 150256 10192 150308 10198
rect 150256 10134 150308 10140
rect 150072 10124 150124 10130
rect 150072 10066 150124 10072
rect 150070 10024 150126 10033
rect 150268 9994 150296 10134
rect 150070 9959 150126 9968
rect 150256 9988 150308 9994
rect 150084 9926 150112 9959
rect 150256 9930 150308 9936
rect 150072 9920 150124 9926
rect 150072 9862 150124 9868
rect 150360 9636 150388 10254
rect 150440 10124 150492 10130
rect 150440 10066 150492 10072
rect 150452 10033 150480 10066
rect 150438 10024 150494 10033
rect 150438 9959 150494 9968
rect 150360 9608 150397 9636
rect 150369 9500 150397 9608
rect 150360 9472 150397 9500
rect 150360 9024 150388 9472
rect 150544 9450 150572 12106
rect 150622 11928 150678 11937
rect 150622 11863 150678 11872
rect 150532 9444 150584 9450
rect 150532 9386 150584 9392
rect 150440 9104 150492 9110
rect 150440 9046 150492 9052
rect 150360 8996 150397 9024
rect 150256 8968 150308 8974
rect 150256 8910 150308 8916
rect 150268 8786 150296 8910
rect 150176 8758 150296 8786
rect 150176 8673 150204 8758
rect 150162 8664 150218 8673
rect 150369 8650 150397 8996
rect 150162 8599 150218 8608
rect 150268 8622 150397 8650
rect 150164 8424 150216 8430
rect 150164 8366 150216 8372
rect 149992 8266 150112 8294
rect 149888 8084 149940 8090
rect 149888 8026 149940 8032
rect 149796 7200 149848 7206
rect 149796 7142 149848 7148
rect 149704 6928 149756 6934
rect 149704 6870 149756 6876
rect 149716 6798 149744 6870
rect 149704 6792 149756 6798
rect 149704 6734 149756 6740
rect 149808 6458 149836 7142
rect 150084 7002 150112 8266
rect 150176 8265 150204 8366
rect 150162 8256 150218 8265
rect 150162 8191 150218 8200
rect 150164 8084 150216 8090
rect 150164 8026 150216 8032
rect 150176 7818 150204 8026
rect 150164 7812 150216 7818
rect 150164 7754 150216 7760
rect 150072 6996 150124 7002
rect 150072 6938 150124 6944
rect 150268 6798 150296 8622
rect 150452 7546 150480 9046
rect 150532 8832 150584 8838
rect 150532 8774 150584 8780
rect 150544 8673 150572 8774
rect 150530 8664 150586 8673
rect 150530 8599 150586 8608
rect 150532 7880 150584 7886
rect 150532 7822 150584 7828
rect 150440 7540 150492 7546
rect 150440 7482 150492 7488
rect 150440 6860 150492 6866
rect 150440 6802 150492 6808
rect 150256 6792 150308 6798
rect 150308 6752 150388 6780
rect 150256 6734 150308 6740
rect 150164 6656 150216 6662
rect 150164 6598 150216 6604
rect 149796 6452 149848 6458
rect 149796 6394 149848 6400
rect 149888 6452 149940 6458
rect 149888 6394 149940 6400
rect 149808 5930 149836 6394
rect 149900 6225 149928 6394
rect 149886 6216 149942 6225
rect 149886 6151 149942 6160
rect 150072 6180 150124 6186
rect 150072 6122 150124 6128
rect 149808 5902 150020 5930
rect 149888 5840 149940 5846
rect 149888 5782 149940 5788
rect 149702 5672 149758 5681
rect 149702 5607 149758 5616
rect 149716 5574 149744 5607
rect 149704 5568 149756 5574
rect 149704 5510 149756 5516
rect 149796 5228 149848 5234
rect 149796 5170 149848 5176
rect 149704 5024 149756 5030
rect 149704 4966 149756 4972
rect 149532 4780 149652 4808
rect 149428 4480 149480 4486
rect 149428 4422 149480 4428
rect 149244 4208 149296 4214
rect 149244 4150 149296 4156
rect 149058 4040 149114 4049
rect 149242 4040 149298 4049
rect 149058 3975 149114 3984
rect 149164 3998 149242 4026
rect 149060 3528 149112 3534
rect 149060 3470 149112 3476
rect 148876 2644 148928 2650
rect 148876 2586 148928 2592
rect 148968 2644 149020 2650
rect 148968 2586 149020 2592
rect 148784 2440 148836 2446
rect 148784 2382 148836 2388
rect 149072 2106 149100 3470
rect 149164 3398 149192 3998
rect 149242 3975 149298 3984
rect 149532 3890 149560 4780
rect 149532 3862 149652 3890
rect 149624 3738 149652 3862
rect 149520 3732 149572 3738
rect 149520 3674 149572 3680
rect 149612 3732 149664 3738
rect 149612 3674 149664 3680
rect 149152 3392 149204 3398
rect 149152 3334 149204 3340
rect 149244 3392 149296 3398
rect 149244 3334 149296 3340
rect 149164 2990 149192 3334
rect 149152 2984 149204 2990
rect 149152 2926 149204 2932
rect 149152 2372 149204 2378
rect 149152 2314 149204 2320
rect 149060 2100 149112 2106
rect 149060 2042 149112 2048
rect 148138 2000 148194 2009
rect 149164 1970 149192 2314
rect 148138 1935 148194 1944
rect 149152 1964 149204 1970
rect 149152 1906 149204 1912
rect 147772 1828 147824 1834
rect 147772 1770 147824 1776
rect 147864 1828 147916 1834
rect 147864 1770 147916 1776
rect 146208 1692 146260 1698
rect 146208 1634 146260 1640
rect 147784 1562 147812 1770
rect 149256 1737 149284 3334
rect 149532 3058 149560 3674
rect 149716 3641 149744 4966
rect 149808 4457 149836 5170
rect 149900 4486 149928 5782
rect 149888 4480 149940 4486
rect 149794 4448 149850 4457
rect 149888 4422 149940 4428
rect 149794 4383 149850 4392
rect 149888 4140 149940 4146
rect 149888 4082 149940 4088
rect 149702 3632 149758 3641
rect 149702 3567 149758 3576
rect 149428 3052 149480 3058
rect 149428 2994 149480 3000
rect 149520 3052 149572 3058
rect 149520 2994 149572 3000
rect 149440 2582 149468 2994
rect 149428 2576 149480 2582
rect 149428 2518 149480 2524
rect 149610 2544 149666 2553
rect 149716 2514 149744 3567
rect 149900 3466 149928 4082
rect 149992 3466 150020 5902
rect 150084 4758 150112 6122
rect 150176 5574 150204 6598
rect 150256 6316 150308 6322
rect 150256 6258 150308 6264
rect 150268 6225 150296 6258
rect 150254 6216 150310 6225
rect 150254 6151 150310 6160
rect 150256 6112 150308 6118
rect 150256 6054 150308 6060
rect 150164 5568 150216 5574
rect 150164 5510 150216 5516
rect 150268 5302 150296 6054
rect 150360 5302 150388 6752
rect 150452 6662 150480 6802
rect 150440 6656 150492 6662
rect 150440 6598 150492 6604
rect 150440 6452 150492 6458
rect 150440 6394 150492 6400
rect 150452 6361 150480 6394
rect 150438 6352 150494 6361
rect 150438 6287 150494 6296
rect 150256 5296 150308 5302
rect 150256 5238 150308 5244
rect 150348 5296 150400 5302
rect 150348 5238 150400 5244
rect 150348 5092 150400 5098
rect 150348 5034 150400 5040
rect 150072 4752 150124 4758
rect 150072 4694 150124 4700
rect 150072 4072 150124 4078
rect 150072 4014 150124 4020
rect 150084 3505 150112 4014
rect 150164 3732 150216 3738
rect 150164 3674 150216 3680
rect 150070 3496 150126 3505
rect 149888 3460 149940 3466
rect 149888 3402 149940 3408
rect 149980 3460 150032 3466
rect 150070 3431 150126 3440
rect 149980 3402 150032 3408
rect 150176 3194 150204 3674
rect 150164 3188 150216 3194
rect 150164 3130 150216 3136
rect 150256 2576 150308 2582
rect 150256 2518 150308 2524
rect 149610 2479 149666 2488
rect 149704 2508 149756 2514
rect 149624 2310 149652 2479
rect 149704 2450 149756 2456
rect 149612 2304 149664 2310
rect 149612 2246 149664 2252
rect 149624 2145 149652 2246
rect 149610 2136 149666 2145
rect 150268 2106 150296 2518
rect 150360 2446 150388 5034
rect 150438 3360 150494 3369
rect 150438 3295 150494 3304
rect 150452 2582 150480 3295
rect 150544 3058 150572 7822
rect 150636 5846 150664 11863
rect 150728 10810 150756 14826
rect 152464 14816 152516 14822
rect 152464 14758 152516 14764
rect 150808 14476 150860 14482
rect 150808 14418 150860 14424
rect 150820 13462 150848 14418
rect 150990 14376 151046 14385
rect 150990 14311 151046 14320
rect 150808 13456 150860 13462
rect 150808 13398 150860 13404
rect 150900 13320 150952 13326
rect 150900 13262 150952 13268
rect 150912 12986 150940 13262
rect 150900 12980 150952 12986
rect 150900 12922 150952 12928
rect 150806 12744 150862 12753
rect 150806 12679 150808 12688
rect 150860 12679 150862 12688
rect 150808 12650 150860 12656
rect 150808 11688 150860 11694
rect 150860 11648 150940 11676
rect 150808 11630 150860 11636
rect 150808 11348 150860 11354
rect 150808 11290 150860 11296
rect 150716 10804 150768 10810
rect 150716 10746 150768 10752
rect 150716 9920 150768 9926
rect 150716 9862 150768 9868
rect 150624 5840 150676 5846
rect 150624 5782 150676 5788
rect 150624 3460 150676 3466
rect 150624 3402 150676 3408
rect 150636 3058 150664 3402
rect 150728 3194 150756 9862
rect 150820 8634 150848 11290
rect 150912 10810 150940 11648
rect 151004 11354 151032 14311
rect 152476 13938 152504 14758
rect 152648 14680 152700 14686
rect 152648 14622 152700 14628
rect 152556 14272 152608 14278
rect 152556 14214 152608 14220
rect 152464 13932 152516 13938
rect 152464 13874 152516 13880
rect 152280 13864 152332 13870
rect 152280 13806 152332 13812
rect 151268 13524 151320 13530
rect 151268 13466 151320 13472
rect 151820 13524 151872 13530
rect 151820 13466 151872 13472
rect 151084 12164 151136 12170
rect 151084 12106 151136 12112
rect 150992 11348 151044 11354
rect 150992 11290 151044 11296
rect 150900 10804 150952 10810
rect 150900 10746 150952 10752
rect 150900 10532 150952 10538
rect 150900 10474 150952 10480
rect 150912 9926 150940 10474
rect 150900 9920 150952 9926
rect 150900 9862 150952 9868
rect 150992 9716 151044 9722
rect 150992 9658 151044 9664
rect 151004 9586 151032 9658
rect 150992 9580 151044 9586
rect 150992 9522 151044 9528
rect 150900 8900 150952 8906
rect 150900 8842 150952 8848
rect 150912 8809 150940 8842
rect 150992 8832 151044 8838
rect 150898 8800 150954 8809
rect 150992 8774 151044 8780
rect 150898 8735 150954 8744
rect 150808 8628 150860 8634
rect 150808 8570 150860 8576
rect 150900 8628 150952 8634
rect 150900 8570 150952 8576
rect 150912 8430 150940 8570
rect 150900 8424 150952 8430
rect 150900 8366 150952 8372
rect 150900 7948 150952 7954
rect 150900 7890 150952 7896
rect 150806 7576 150862 7585
rect 150806 7511 150808 7520
rect 150860 7511 150862 7520
rect 150808 7482 150860 7488
rect 150808 5024 150860 5030
rect 150808 4966 150860 4972
rect 150716 3188 150768 3194
rect 150716 3130 150768 3136
rect 150532 3052 150584 3058
rect 150532 2994 150584 3000
rect 150624 3052 150676 3058
rect 150624 2994 150676 3000
rect 150440 2576 150492 2582
rect 150440 2518 150492 2524
rect 150348 2440 150400 2446
rect 150348 2382 150400 2388
rect 150346 2136 150402 2145
rect 149610 2071 149666 2080
rect 150256 2100 150308 2106
rect 150346 2071 150402 2080
rect 150256 2042 150308 2048
rect 150360 2038 150388 2071
rect 150348 2032 150400 2038
rect 150348 1974 150400 1980
rect 149242 1728 149298 1737
rect 149242 1663 149298 1672
rect 147772 1556 147824 1562
rect 147772 1498 147824 1504
rect 150820 1154 150848 4966
rect 150912 4457 150940 7890
rect 151004 6304 151032 8774
rect 151096 8634 151124 12106
rect 151280 11150 151308 13466
rect 151832 13190 151860 13466
rect 152292 13410 152320 13806
rect 152292 13394 152412 13410
rect 152292 13388 152424 13394
rect 152292 13382 152372 13388
rect 152372 13330 152424 13336
rect 152464 13320 152516 13326
rect 152464 13262 152516 13268
rect 151820 13184 151872 13190
rect 151820 13126 151872 13132
rect 152372 13184 152424 13190
rect 152372 13126 152424 13132
rect 152004 12980 152056 12986
rect 152056 12940 152320 12968
rect 152004 12922 152056 12928
rect 151360 12912 151412 12918
rect 151360 12854 151412 12860
rect 151372 12238 151400 12854
rect 151360 12232 151412 12238
rect 151360 12174 151412 12180
rect 151372 11218 151400 12174
rect 151912 12096 151964 12102
rect 151912 12038 151964 12044
rect 151450 11656 151506 11665
rect 151450 11591 151506 11600
rect 151360 11212 151412 11218
rect 151360 11154 151412 11160
rect 151268 11144 151320 11150
rect 151268 11086 151320 11092
rect 151266 10024 151322 10033
rect 151266 9959 151322 9968
rect 151360 9988 151412 9994
rect 151280 9722 151308 9959
rect 151360 9930 151412 9936
rect 151268 9716 151320 9722
rect 151268 9658 151320 9664
rect 151174 8936 151230 8945
rect 151174 8871 151230 8880
rect 151084 8628 151136 8634
rect 151084 8570 151136 8576
rect 151188 8498 151216 8871
rect 151176 8492 151228 8498
rect 151176 8434 151228 8440
rect 151084 8288 151136 8294
rect 151084 8230 151136 8236
rect 151096 8129 151124 8230
rect 151082 8120 151138 8129
rect 151082 8055 151138 8064
rect 151266 8120 151322 8129
rect 151266 8055 151322 8064
rect 151176 7880 151228 7886
rect 151176 7822 151228 7828
rect 151084 7540 151136 7546
rect 151084 7482 151136 7488
rect 151096 7177 151124 7482
rect 151082 7168 151138 7177
rect 151082 7103 151138 7112
rect 151084 6316 151136 6322
rect 151004 6276 151084 6304
rect 151084 6258 151136 6264
rect 150990 6216 151046 6225
rect 150990 6151 151046 6160
rect 150898 4448 150954 4457
rect 150898 4383 150954 4392
rect 150900 3936 150952 3942
rect 150900 3878 150952 3884
rect 150912 1290 150940 3878
rect 151004 2530 151032 6151
rect 151084 5568 151136 5574
rect 151084 5510 151136 5516
rect 151096 5273 151124 5510
rect 151082 5264 151138 5273
rect 151082 5199 151138 5208
rect 151084 4548 151136 4554
rect 151084 4490 151136 4496
rect 151096 3369 151124 4490
rect 151082 3360 151138 3369
rect 151082 3295 151138 3304
rect 151004 2502 151124 2530
rect 151096 2378 151124 2502
rect 151084 2372 151136 2378
rect 151084 2314 151136 2320
rect 150900 1284 150952 1290
rect 150900 1226 150952 1232
rect 150808 1148 150860 1154
rect 150808 1090 150860 1096
rect 151188 1086 151216 7822
rect 151280 6798 151308 8055
rect 151268 6792 151320 6798
rect 151268 6734 151320 6740
rect 151372 5273 151400 9930
rect 151464 9926 151492 11591
rect 151544 11008 151596 11014
rect 151544 10950 151596 10956
rect 151452 9920 151504 9926
rect 151452 9862 151504 9868
rect 151452 9512 151504 9518
rect 151452 9454 151504 9460
rect 151464 6934 151492 9454
rect 151556 7750 151584 10950
rect 151636 10668 151688 10674
rect 151636 10610 151688 10616
rect 151648 10554 151676 10610
rect 151648 10526 151860 10554
rect 151726 10432 151782 10441
rect 151726 10367 151782 10376
rect 151740 9722 151768 10367
rect 151728 9716 151780 9722
rect 151728 9658 151780 9664
rect 151636 9444 151688 9450
rect 151636 9386 151688 9392
rect 151648 8974 151676 9386
rect 151832 9110 151860 10526
rect 151820 9104 151872 9110
rect 151820 9046 151872 9052
rect 151636 8968 151688 8974
rect 151636 8910 151688 8916
rect 151728 8900 151780 8906
rect 151728 8842 151780 8848
rect 151636 8560 151688 8566
rect 151636 8502 151688 8508
rect 151544 7744 151596 7750
rect 151544 7686 151596 7692
rect 151452 6928 151504 6934
rect 151452 6870 151504 6876
rect 151542 6624 151598 6633
rect 151542 6559 151598 6568
rect 151556 5794 151584 6559
rect 151648 6186 151676 8502
rect 151740 6798 151768 8842
rect 151820 8492 151872 8498
rect 151820 8434 151872 8440
rect 151832 8090 151860 8434
rect 151820 8084 151872 8090
rect 151820 8026 151872 8032
rect 151820 7744 151872 7750
rect 151820 7686 151872 7692
rect 151728 6792 151780 6798
rect 151728 6734 151780 6740
rect 151636 6180 151688 6186
rect 151636 6122 151688 6128
rect 151556 5766 151676 5794
rect 151544 5704 151596 5710
rect 151544 5646 151596 5652
rect 151452 5636 151504 5642
rect 151452 5578 151504 5584
rect 151358 5264 151414 5273
rect 151358 5199 151414 5208
rect 151464 4826 151492 5578
rect 151268 4820 151320 4826
rect 151268 4762 151320 4768
rect 151452 4820 151504 4826
rect 151452 4762 151504 4768
rect 151280 4593 151308 4762
rect 151266 4584 151322 4593
rect 151266 4519 151322 4528
rect 151268 4072 151320 4078
rect 151320 4032 151400 4060
rect 151268 4014 151320 4020
rect 151268 3392 151320 3398
rect 151268 3334 151320 3340
rect 151280 2922 151308 3334
rect 151372 3058 151400 4032
rect 151464 3126 151492 4762
rect 151556 4146 151584 5646
rect 151648 4554 151676 5766
rect 151832 5386 151860 7686
rect 151924 5710 151952 12038
rect 152096 10668 152148 10674
rect 152096 10610 152148 10616
rect 152004 9988 152056 9994
rect 152108 9976 152136 10610
rect 152292 10470 152320 12940
rect 152384 11626 152412 13126
rect 152476 12918 152504 13262
rect 152464 12912 152516 12918
rect 152464 12854 152516 12860
rect 152372 11620 152424 11626
rect 152372 11562 152424 11568
rect 152476 11218 152504 12854
rect 152568 11898 152596 14214
rect 152660 12714 152688 14622
rect 153384 14340 153436 14346
rect 153384 14282 153436 14288
rect 153200 14136 153252 14142
rect 153200 14078 153252 14084
rect 153212 13546 153240 14078
rect 153292 13728 153344 13734
rect 153292 13670 153344 13676
rect 153120 13518 153240 13546
rect 152832 13320 152884 13326
rect 152832 13262 152884 13268
rect 152740 13252 152792 13258
rect 152740 13194 152792 13200
rect 152648 12708 152700 12714
rect 152648 12650 152700 12656
rect 152752 12646 152780 13194
rect 152740 12640 152792 12646
rect 152740 12582 152792 12588
rect 152648 12232 152700 12238
rect 152648 12174 152700 12180
rect 152556 11892 152608 11898
rect 152556 11834 152608 11840
rect 152660 11529 152688 12174
rect 152646 11520 152702 11529
rect 152646 11455 152702 11464
rect 152464 11212 152516 11218
rect 152464 11154 152516 11160
rect 152370 11112 152426 11121
rect 152370 11047 152426 11056
rect 152280 10464 152332 10470
rect 152280 10406 152332 10412
rect 152056 9948 152136 9976
rect 152004 9930 152056 9936
rect 152188 9920 152240 9926
rect 152186 9888 152188 9897
rect 152280 9920 152332 9926
rect 152240 9888 152242 9897
rect 152280 9862 152332 9868
rect 152186 9823 152242 9832
rect 152002 9616 152058 9625
rect 152002 9551 152058 9560
rect 152096 9580 152148 9586
rect 152016 9042 152044 9551
rect 152148 9540 152228 9568
rect 152096 9522 152148 9528
rect 152004 9036 152056 9042
rect 152004 8978 152056 8984
rect 152096 8968 152148 8974
rect 152096 8910 152148 8916
rect 152004 8424 152056 8430
rect 152002 8392 152004 8401
rect 152056 8392 152058 8401
rect 152002 8327 152058 8336
rect 152002 7576 152058 7585
rect 152002 7511 152058 7520
rect 151912 5704 151964 5710
rect 151912 5646 151964 5652
rect 152016 5409 152044 7511
rect 152108 6798 152136 8910
rect 152200 7750 152228 9540
rect 152292 9382 152320 9862
rect 152280 9376 152332 9382
rect 152280 9318 152332 9324
rect 152384 8809 152412 11047
rect 152476 10674 152504 11154
rect 152556 10804 152608 10810
rect 152556 10746 152608 10752
rect 152464 10668 152516 10674
rect 152464 10610 152516 10616
rect 152568 10418 152596 10746
rect 152646 10704 152702 10713
rect 152646 10639 152702 10648
rect 152660 10538 152688 10639
rect 152648 10532 152700 10538
rect 152648 10474 152700 10480
rect 152568 10390 152688 10418
rect 152554 9616 152610 9625
rect 152554 9551 152556 9560
rect 152608 9551 152610 9560
rect 152556 9522 152608 9528
rect 152660 9518 152688 10390
rect 152648 9512 152700 9518
rect 152648 9454 152700 9460
rect 152464 8968 152516 8974
rect 152464 8910 152516 8916
rect 152556 8968 152608 8974
rect 152556 8910 152608 8916
rect 152370 8800 152426 8809
rect 152370 8735 152426 8744
rect 152280 8424 152332 8430
rect 152280 8366 152332 8372
rect 152292 8090 152320 8366
rect 152280 8084 152332 8090
rect 152280 8026 152332 8032
rect 152372 8084 152424 8090
rect 152372 8026 152424 8032
rect 152384 7886 152412 8026
rect 152280 7880 152332 7886
rect 152280 7822 152332 7828
rect 152372 7880 152424 7886
rect 152372 7822 152424 7828
rect 152188 7744 152240 7750
rect 152188 7686 152240 7692
rect 152188 7336 152240 7342
rect 152188 7278 152240 7284
rect 152200 6866 152228 7278
rect 152188 6860 152240 6866
rect 152188 6802 152240 6808
rect 152096 6792 152148 6798
rect 152096 6734 152148 6740
rect 152200 6730 152228 6802
rect 152188 6724 152240 6730
rect 152188 6666 152240 6672
rect 151740 5358 151860 5386
rect 152002 5400 152058 5409
rect 151636 4548 151688 4554
rect 151636 4490 151688 4496
rect 151544 4140 151596 4146
rect 151544 4082 151596 4088
rect 151542 3496 151598 3505
rect 151542 3431 151544 3440
rect 151596 3431 151598 3440
rect 151544 3402 151596 3408
rect 151452 3120 151504 3126
rect 151452 3062 151504 3068
rect 151360 3052 151412 3058
rect 151360 2994 151412 3000
rect 151268 2916 151320 2922
rect 151268 2858 151320 2864
rect 151740 2310 151768 5358
rect 152002 5335 152058 5344
rect 151820 5296 151872 5302
rect 151872 5256 151952 5284
rect 151820 5238 151872 5244
rect 151820 4616 151872 4622
rect 151820 4558 151872 4564
rect 151832 4214 151860 4558
rect 151820 4208 151872 4214
rect 151820 4150 151872 4156
rect 151832 3602 151860 4150
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 151924 2990 151952 5256
rect 152016 4146 152044 5335
rect 152200 5166 152228 6666
rect 152188 5160 152240 5166
rect 152292 5137 152320 7822
rect 152384 6633 152412 7822
rect 152370 6624 152426 6633
rect 152370 6559 152426 6568
rect 152476 6497 152504 8910
rect 152568 6633 152596 8910
rect 152554 6624 152610 6633
rect 152554 6559 152610 6568
rect 152462 6488 152518 6497
rect 152462 6423 152518 6432
rect 152372 6316 152424 6322
rect 152372 6258 152424 6264
rect 152384 5846 152412 6258
rect 152568 5930 152596 6559
rect 152648 6112 152700 6118
rect 152648 6054 152700 6060
rect 152476 5902 152596 5930
rect 152372 5840 152424 5846
rect 152372 5782 152424 5788
rect 152476 5545 152504 5902
rect 152462 5536 152518 5545
rect 152462 5471 152518 5480
rect 152372 5228 152424 5234
rect 152372 5170 152424 5176
rect 152188 5102 152240 5108
rect 152278 5128 152334 5137
rect 152278 5063 152334 5072
rect 152188 4752 152240 4758
rect 152094 4720 152150 4729
rect 152188 4694 152240 4700
rect 152094 4655 152150 4664
rect 152108 4622 152136 4655
rect 152096 4616 152148 4622
rect 152096 4558 152148 4564
rect 152004 4140 152056 4146
rect 152004 4082 152056 4088
rect 152004 3120 152056 3126
rect 152004 3062 152056 3068
rect 151820 2984 151872 2990
rect 151818 2952 151820 2961
rect 151912 2984 151964 2990
rect 151872 2952 151874 2961
rect 151912 2926 151964 2932
rect 151818 2887 151874 2896
rect 151728 2304 151780 2310
rect 151728 2246 151780 2252
rect 152016 1358 152044 3062
rect 152200 2650 152228 4694
rect 152280 4480 152332 4486
rect 152280 4422 152332 4428
rect 152292 3126 152320 4422
rect 152280 3120 152332 3126
rect 152280 3062 152332 3068
rect 152188 2644 152240 2650
rect 152188 2586 152240 2592
rect 152384 2553 152412 5170
rect 152476 4758 152504 5471
rect 152660 5166 152688 6054
rect 152648 5160 152700 5166
rect 152648 5102 152700 5108
rect 152556 5092 152608 5098
rect 152556 5034 152608 5040
rect 152464 4752 152516 4758
rect 152464 4694 152516 4700
rect 152464 4072 152516 4078
rect 152568 4060 152596 5034
rect 152516 4032 152596 4060
rect 152464 4014 152516 4020
rect 152568 3602 152596 4032
rect 152556 3596 152608 3602
rect 152556 3538 152608 3544
rect 152464 3528 152516 3534
rect 152462 3496 152464 3505
rect 152660 3505 152688 5102
rect 152752 4146 152780 12582
rect 152844 11121 152872 13262
rect 152922 13016 152978 13025
rect 153120 13002 153148 13518
rect 153198 13424 153254 13433
rect 153198 13359 153254 13368
rect 153212 13190 153240 13359
rect 153304 13258 153332 13670
rect 153396 13326 153424 14282
rect 153568 13796 153620 13802
rect 153568 13738 153620 13744
rect 153580 13530 153608 13738
rect 154316 13530 154344 14962
rect 153568 13524 153620 13530
rect 153568 13466 153620 13472
rect 154304 13524 154356 13530
rect 154304 13466 154356 13472
rect 153384 13320 153436 13326
rect 153384 13262 153436 13268
rect 153476 13320 153528 13326
rect 153476 13262 153528 13268
rect 154118 13288 154174 13297
rect 153292 13252 153344 13258
rect 153292 13194 153344 13200
rect 153200 13184 153252 13190
rect 153200 13126 153252 13132
rect 153120 12974 153240 13002
rect 153488 12986 153516 13262
rect 154118 13223 154174 13232
rect 153752 13184 153804 13190
rect 153752 13126 153804 13132
rect 152922 12951 152924 12960
rect 152976 12951 152978 12960
rect 152924 12922 152976 12928
rect 152922 12608 152978 12617
rect 152922 12543 152978 12552
rect 152830 11112 152886 11121
rect 152830 11047 152886 11056
rect 152832 9104 152884 9110
rect 152832 9046 152884 9052
rect 152844 8838 152872 9046
rect 152832 8832 152884 8838
rect 152832 8774 152884 8780
rect 152832 8492 152884 8498
rect 152832 8434 152884 8440
rect 152844 6934 152872 8434
rect 152936 7954 152964 12543
rect 153106 12472 153162 12481
rect 153106 12407 153108 12416
rect 153160 12407 153162 12416
rect 153108 12378 153160 12384
rect 153016 12232 153068 12238
rect 153016 12174 153068 12180
rect 153028 9518 153056 12174
rect 153212 11354 153240 12974
rect 153476 12980 153528 12986
rect 153476 12922 153528 12928
rect 153764 12850 153792 13126
rect 153384 12844 153436 12850
rect 153384 12786 153436 12792
rect 153752 12844 153804 12850
rect 153752 12786 153804 12792
rect 153396 12753 153424 12786
rect 154132 12782 154160 13223
rect 154408 13190 154436 15030
rect 157432 14748 157484 14754
rect 157432 14690 157484 14696
rect 156696 14612 156748 14618
rect 156696 14554 156748 14560
rect 154948 14544 155000 14550
rect 154948 14486 155000 14492
rect 154856 14408 154908 14414
rect 154856 14350 154908 14356
rect 154868 13326 154896 14350
rect 154856 13320 154908 13326
rect 154856 13262 154908 13268
rect 154212 13184 154264 13190
rect 154212 13126 154264 13132
rect 154396 13184 154448 13190
rect 154396 13126 154448 13132
rect 154120 12776 154172 12782
rect 153382 12744 153438 12753
rect 154120 12718 154172 12724
rect 153382 12679 153438 12688
rect 153752 12164 153804 12170
rect 153752 12106 153804 12112
rect 153474 12064 153530 12073
rect 153474 11999 153530 12008
rect 153292 11892 153344 11898
rect 153292 11834 153344 11840
rect 153304 11762 153332 11834
rect 153292 11756 153344 11762
rect 153292 11698 153344 11704
rect 153488 11354 153516 11999
rect 153200 11348 153252 11354
rect 153200 11290 153252 11296
rect 153476 11348 153528 11354
rect 153476 11290 153528 11296
rect 153660 10192 153712 10198
rect 153660 10134 153712 10140
rect 153672 9586 153700 10134
rect 153292 9580 153344 9586
rect 153292 9522 153344 9528
rect 153660 9580 153712 9586
rect 153660 9522 153712 9528
rect 153016 9512 153068 9518
rect 153304 9489 153332 9522
rect 153476 9512 153528 9518
rect 153016 9454 153068 9460
rect 153290 9480 153346 9489
rect 153476 9454 153528 9460
rect 153658 9480 153714 9489
rect 153290 9415 153346 9424
rect 153108 9376 153160 9382
rect 153108 9318 153160 9324
rect 153016 8356 153068 8362
rect 153016 8298 153068 8304
rect 152924 7948 152976 7954
rect 152924 7890 152976 7896
rect 152832 6928 152884 6934
rect 152832 6870 152884 6876
rect 152832 6792 152884 6798
rect 152832 6734 152884 6740
rect 152844 6662 152872 6734
rect 152832 6656 152884 6662
rect 152832 6598 152884 6604
rect 152844 4826 152872 6598
rect 152924 6452 152976 6458
rect 152924 6394 152976 6400
rect 152936 6254 152964 6394
rect 152924 6248 152976 6254
rect 152924 6190 152976 6196
rect 153028 5030 153056 8298
rect 153120 8129 153148 9318
rect 153488 8974 153516 9454
rect 153658 9415 153714 9424
rect 153568 9172 153620 9178
rect 153568 9114 153620 9120
rect 153476 8968 153528 8974
rect 153476 8910 153528 8916
rect 153580 8673 153608 9114
rect 153672 9110 153700 9415
rect 153660 9104 153712 9110
rect 153660 9046 153712 9052
rect 153660 8900 153712 8906
rect 153660 8842 153712 8848
rect 153566 8664 153622 8673
rect 153566 8599 153622 8608
rect 153672 8412 153700 8842
rect 153764 8566 153792 12106
rect 154224 11830 154252 13126
rect 154302 12744 154358 12753
rect 154302 12679 154358 12688
rect 154316 12646 154344 12679
rect 154304 12640 154356 12646
rect 154304 12582 154356 12588
rect 154764 12368 154816 12374
rect 154764 12310 154816 12316
rect 154672 12232 154724 12238
rect 154500 12180 154672 12186
rect 154500 12174 154724 12180
rect 154500 12158 154712 12174
rect 154212 11824 154264 11830
rect 154500 11778 154528 12158
rect 154776 12084 154804 12310
rect 154212 11766 154264 11772
rect 153936 11756 153988 11762
rect 153936 11698 153988 11704
rect 154316 11750 154528 11778
rect 154592 12056 154804 12084
rect 154592 11762 154620 12056
rect 153948 10810 153976 11698
rect 154316 11694 154344 11750
rect 154304 11688 154356 11694
rect 154304 11630 154356 11636
rect 154396 11688 154448 11694
rect 154396 11630 154448 11636
rect 154408 11540 154436 11630
rect 154316 11512 154436 11540
rect 154028 11076 154080 11082
rect 154028 11018 154080 11024
rect 153936 10804 153988 10810
rect 153936 10746 153988 10752
rect 154040 10606 154068 11018
rect 154028 10600 154080 10606
rect 154028 10542 154080 10548
rect 154212 10600 154264 10606
rect 154212 10542 154264 10548
rect 153844 10192 153896 10198
rect 153842 10160 153844 10169
rect 153896 10160 153898 10169
rect 153842 10095 153898 10104
rect 153936 10124 153988 10130
rect 153936 10066 153988 10072
rect 153948 9654 153976 10066
rect 154040 9926 154068 10542
rect 154028 9920 154080 9926
rect 154028 9862 154080 9868
rect 153936 9648 153988 9654
rect 153936 9590 153988 9596
rect 154040 9450 154068 9862
rect 154028 9444 154080 9450
rect 154028 9386 154080 9392
rect 154120 9444 154172 9450
rect 154120 9386 154172 9392
rect 153844 9376 153896 9382
rect 153844 9318 153896 9324
rect 153752 8560 153804 8566
rect 153752 8502 153804 8508
rect 153672 8384 153792 8412
rect 153476 8288 153528 8294
rect 153476 8230 153528 8236
rect 153660 8288 153712 8294
rect 153660 8230 153712 8236
rect 153106 8120 153162 8129
rect 153106 8055 153162 8064
rect 153384 7744 153436 7750
rect 153384 7686 153436 7692
rect 153292 7336 153344 7342
rect 153292 7278 153344 7284
rect 153198 6896 153254 6905
rect 153198 6831 153254 6840
rect 153212 5778 153240 6831
rect 153108 5772 153160 5778
rect 153108 5714 153160 5720
rect 153200 5772 153252 5778
rect 153200 5714 153252 5720
rect 153016 5024 153068 5030
rect 153016 4966 153068 4972
rect 152832 4820 152884 4826
rect 152832 4762 152884 4768
rect 152924 4820 152976 4826
rect 152924 4762 152976 4768
rect 152936 4593 152964 4762
rect 152922 4584 152978 4593
rect 152922 4519 152978 4528
rect 152740 4140 152792 4146
rect 152740 4082 152792 4088
rect 152516 3496 152518 3505
rect 152462 3431 152518 3440
rect 152646 3496 152702 3505
rect 152646 3431 152702 3440
rect 152752 2650 152780 4082
rect 152830 3768 152886 3777
rect 152830 3703 152832 3712
rect 152884 3703 152886 3712
rect 153014 3768 153070 3777
rect 153014 3703 153070 3712
rect 152832 3674 152884 3680
rect 153028 2990 153056 3703
rect 153120 3534 153148 5714
rect 153304 4026 153332 7278
rect 153396 6322 153424 7686
rect 153488 7274 153516 8230
rect 153672 7410 153700 8230
rect 153764 7886 153792 8384
rect 153752 7880 153804 7886
rect 153752 7822 153804 7828
rect 153660 7404 153712 7410
rect 153660 7346 153712 7352
rect 153568 7336 153620 7342
rect 153568 7278 153620 7284
rect 153476 7268 153528 7274
rect 153476 7210 153528 7216
rect 153474 6760 153530 6769
rect 153474 6695 153530 6704
rect 153488 6662 153516 6695
rect 153476 6656 153528 6662
rect 153476 6598 153528 6604
rect 153580 6474 153608 7278
rect 153764 7018 153792 7822
rect 153488 6446 153608 6474
rect 153672 6990 153792 7018
rect 153384 6316 153436 6322
rect 153384 6258 153436 6264
rect 153488 6254 153516 6446
rect 153566 6352 153622 6361
rect 153566 6287 153622 6296
rect 153476 6248 153528 6254
rect 153476 6190 153528 6196
rect 153384 5160 153436 5166
rect 153384 5102 153436 5108
rect 153212 3998 153332 4026
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 153016 2984 153068 2990
rect 153016 2926 153068 2932
rect 153212 2922 153240 3998
rect 153292 3936 153344 3942
rect 153292 3878 153344 3884
rect 153304 3233 153332 3878
rect 153396 3398 153424 5102
rect 153488 4604 153516 6190
rect 153580 5710 153608 6287
rect 153672 6118 153700 6990
rect 153752 6928 153804 6934
rect 153752 6870 153804 6876
rect 153764 6322 153792 6870
rect 153752 6316 153804 6322
rect 153752 6258 153804 6264
rect 153660 6112 153712 6118
rect 153660 6054 153712 6060
rect 153672 5710 153700 6054
rect 153568 5704 153620 5710
rect 153568 5646 153620 5652
rect 153660 5704 153712 5710
rect 153660 5646 153712 5652
rect 153568 4616 153620 4622
rect 153488 4576 153568 4604
rect 153568 4558 153620 4564
rect 153660 4616 153712 4622
rect 153660 4558 153712 4564
rect 153580 4049 153608 4558
rect 153566 4040 153622 4049
rect 153566 3975 153622 3984
rect 153384 3392 153436 3398
rect 153384 3334 153436 3340
rect 153474 3360 153530 3369
rect 153474 3295 153530 3304
rect 153290 3224 153346 3233
rect 153290 3159 153346 3168
rect 153488 2922 153516 3295
rect 153200 2916 153252 2922
rect 153200 2858 153252 2864
rect 153476 2916 153528 2922
rect 153476 2858 153528 2864
rect 152740 2644 152792 2650
rect 152740 2586 152792 2592
rect 152370 2544 152426 2553
rect 152370 2479 152426 2488
rect 153672 2417 153700 4558
rect 153752 3392 153804 3398
rect 153752 3334 153804 3340
rect 153658 2408 153714 2417
rect 153658 2343 153714 2352
rect 152004 1352 152056 1358
rect 152004 1294 152056 1300
rect 153764 1193 153792 3334
rect 153856 3058 153884 9318
rect 153936 8968 153988 8974
rect 153936 8910 153988 8916
rect 153948 7342 153976 8910
rect 154040 7886 154068 9386
rect 154028 7880 154080 7886
rect 154028 7822 154080 7828
rect 154028 7744 154080 7750
rect 154028 7686 154080 7692
rect 153936 7336 153988 7342
rect 153936 7278 153988 7284
rect 154040 6474 154068 7686
rect 154132 7041 154160 9386
rect 154224 8974 154252 10542
rect 154316 10538 154344 11512
rect 154396 11076 154448 11082
rect 154500 11064 154528 11750
rect 154580 11756 154632 11762
rect 154580 11698 154632 11704
rect 154672 11756 154724 11762
rect 154672 11698 154724 11704
rect 154684 11393 154712 11698
rect 154670 11384 154726 11393
rect 154670 11319 154726 11328
rect 154448 11036 154528 11064
rect 154856 11076 154908 11082
rect 154396 11018 154448 11024
rect 154856 11018 154908 11024
rect 154580 10804 154632 10810
rect 154580 10746 154632 10752
rect 154396 10668 154448 10674
rect 154396 10610 154448 10616
rect 154304 10532 154356 10538
rect 154304 10474 154356 10480
rect 154316 9518 154344 10474
rect 154304 9512 154356 9518
rect 154304 9454 154356 9460
rect 154212 8968 154264 8974
rect 154212 8910 154264 8916
rect 154316 8820 154344 9454
rect 154224 8792 154344 8820
rect 154224 8566 154252 8792
rect 154212 8560 154264 8566
rect 154212 8502 154264 8508
rect 154304 8492 154356 8498
rect 154304 8434 154356 8440
rect 154212 8424 154264 8430
rect 154316 8401 154344 8434
rect 154212 8366 154264 8372
rect 154302 8392 154358 8401
rect 154118 7032 154174 7041
rect 154118 6967 154174 6976
rect 154040 6446 154160 6474
rect 154028 6316 154080 6322
rect 154028 6258 154080 6264
rect 153934 6216 153990 6225
rect 153934 6151 153936 6160
rect 153988 6151 153990 6160
rect 153936 6122 153988 6128
rect 153936 5840 153988 5846
rect 153936 5782 153988 5788
rect 153948 3398 153976 5782
rect 154040 5234 154068 6258
rect 154132 5846 154160 6446
rect 154120 5840 154172 5846
rect 154120 5782 154172 5788
rect 154120 5704 154172 5710
rect 154120 5646 154172 5652
rect 154028 5228 154080 5234
rect 154028 5170 154080 5176
rect 154132 5166 154160 5646
rect 154120 5160 154172 5166
rect 154120 5102 154172 5108
rect 154120 5024 154172 5030
rect 154120 4966 154172 4972
rect 153936 3392 153988 3398
rect 153936 3334 153988 3340
rect 153844 3052 153896 3058
rect 153844 2994 153896 3000
rect 154028 2984 154080 2990
rect 154026 2952 154028 2961
rect 154080 2952 154082 2961
rect 154026 2887 154082 2896
rect 154132 2514 154160 4966
rect 154224 2854 154252 8366
rect 154302 8327 154358 8336
rect 154304 8288 154356 8294
rect 154304 8230 154356 8236
rect 154316 8022 154344 8230
rect 154304 8016 154356 8022
rect 154304 7958 154356 7964
rect 154302 7440 154358 7449
rect 154302 7375 154304 7384
rect 154356 7375 154358 7384
rect 154304 7346 154356 7352
rect 154408 7290 154436 10610
rect 154592 8673 154620 10746
rect 154672 10668 154724 10674
rect 154672 10610 154724 10616
rect 154684 10305 154712 10610
rect 154670 10296 154726 10305
rect 154670 10231 154726 10240
rect 154672 10056 154724 10062
rect 154670 10024 154672 10033
rect 154724 10024 154726 10033
rect 154670 9959 154726 9968
rect 154672 9580 154724 9586
rect 154672 9522 154724 9528
rect 154684 9178 154712 9522
rect 154764 9512 154816 9518
rect 154764 9454 154816 9460
rect 154672 9172 154724 9178
rect 154672 9114 154724 9120
rect 154578 8664 154634 8673
rect 154578 8599 154634 8608
rect 154488 8356 154540 8362
rect 154488 8298 154540 8304
rect 154316 7262 154436 7290
rect 154316 6118 154344 7262
rect 154396 7200 154448 7206
rect 154396 7142 154448 7148
rect 154304 6112 154356 6118
rect 154304 6054 154356 6060
rect 154302 5536 154358 5545
rect 154302 5471 154358 5480
rect 154316 5302 154344 5471
rect 154304 5296 154356 5302
rect 154304 5238 154356 5244
rect 154302 5128 154358 5137
rect 154302 5063 154358 5072
rect 154316 4758 154344 5063
rect 154304 4752 154356 4758
rect 154304 4694 154356 4700
rect 154304 3528 154356 3534
rect 154304 3470 154356 3476
rect 154316 3369 154344 3470
rect 154302 3360 154358 3369
rect 154302 3295 154358 3304
rect 154408 3194 154436 7142
rect 154500 6322 154528 8298
rect 154592 7546 154620 8599
rect 154580 7540 154632 7546
rect 154580 7482 154632 7488
rect 154580 6724 154632 6730
rect 154580 6666 154632 6672
rect 154488 6316 154540 6322
rect 154488 6258 154540 6264
rect 154592 6202 154620 6666
rect 154500 6174 154620 6202
rect 154500 5846 154528 6174
rect 154684 5930 154712 9114
rect 154776 9110 154804 9454
rect 154764 9104 154816 9110
rect 154764 9046 154816 9052
rect 154764 8424 154816 8430
rect 154764 8366 154816 8372
rect 154776 8090 154804 8366
rect 154764 8084 154816 8090
rect 154764 8026 154816 8032
rect 154764 7336 154816 7342
rect 154764 7278 154816 7284
rect 154776 7206 154804 7278
rect 154764 7200 154816 7206
rect 154764 7142 154816 7148
rect 154776 6633 154804 7142
rect 154762 6624 154818 6633
rect 154762 6559 154818 6568
rect 154868 6361 154896 11018
rect 154854 6352 154910 6361
rect 154854 6287 154910 6296
rect 154592 5902 154712 5930
rect 154488 5840 154540 5846
rect 154488 5782 154540 5788
rect 154592 4706 154620 5902
rect 154960 5846 154988 14486
rect 156052 14204 156104 14210
rect 156052 14146 156104 14152
rect 155960 14068 156012 14074
rect 155960 14010 156012 14016
rect 155866 13696 155922 13705
rect 155866 13631 155922 13640
rect 155774 13560 155830 13569
rect 155880 13530 155908 13631
rect 155774 13495 155830 13504
rect 155868 13524 155920 13530
rect 155788 13462 155816 13495
rect 155868 13466 155920 13472
rect 155684 13456 155736 13462
rect 155684 13398 155736 13404
rect 155776 13456 155828 13462
rect 155776 13398 155828 13404
rect 155408 12912 155460 12918
rect 155408 12854 155460 12860
rect 155592 12912 155644 12918
rect 155592 12854 155644 12860
rect 155224 12232 155276 12238
rect 155224 12174 155276 12180
rect 155236 11218 155264 12174
rect 155316 11824 155368 11830
rect 155314 11792 155316 11801
rect 155368 11792 155370 11801
rect 155314 11727 155370 11736
rect 155420 11558 155448 12854
rect 155500 12232 155552 12238
rect 155500 12174 155552 12180
rect 155512 11626 155540 12174
rect 155500 11620 155552 11626
rect 155500 11562 155552 11568
rect 155316 11552 155368 11558
rect 155316 11494 155368 11500
rect 155408 11552 155460 11558
rect 155408 11494 155460 11500
rect 155224 11212 155276 11218
rect 155224 11154 155276 11160
rect 155222 10840 155278 10849
rect 155328 10810 155356 11494
rect 155500 11212 155552 11218
rect 155500 11154 155552 11160
rect 155408 11008 155460 11014
rect 155408 10950 155460 10956
rect 155222 10775 155278 10784
rect 155316 10804 155368 10810
rect 155236 10470 155264 10775
rect 155316 10746 155368 10752
rect 155224 10464 155276 10470
rect 155224 10406 155276 10412
rect 155328 9654 155356 10746
rect 155420 10742 155448 10950
rect 155408 10736 155460 10742
rect 155408 10678 155460 10684
rect 155408 10464 155460 10470
rect 155408 10406 155460 10412
rect 155420 10130 155448 10406
rect 155408 10124 155460 10130
rect 155408 10066 155460 10072
rect 155408 9920 155460 9926
rect 155408 9862 155460 9868
rect 155316 9648 155368 9654
rect 155316 9590 155368 9596
rect 155040 9580 155092 9586
rect 155040 9522 155092 9528
rect 155052 9042 155080 9522
rect 155040 9036 155092 9042
rect 155040 8978 155092 8984
rect 155224 8968 155276 8974
rect 155224 8910 155276 8916
rect 155040 8832 155092 8838
rect 155236 8809 155264 8910
rect 155040 8774 155092 8780
rect 155222 8800 155278 8809
rect 154948 5840 155000 5846
rect 154670 5808 154726 5817
rect 154948 5782 155000 5788
rect 154670 5743 154726 5752
rect 154684 5710 154712 5743
rect 154672 5704 154724 5710
rect 154672 5646 154724 5652
rect 155052 5250 155080 8774
rect 155222 8735 155278 8744
rect 155328 8634 155356 9590
rect 155316 8628 155368 8634
rect 155316 8570 155368 8576
rect 155224 6860 155276 6866
rect 155328 6848 155356 8570
rect 155420 8401 155448 9862
rect 155512 9518 155540 11154
rect 155500 9512 155552 9518
rect 155500 9454 155552 9460
rect 155406 8392 155462 8401
rect 155406 8327 155462 8336
rect 155408 8288 155460 8294
rect 155408 8230 155460 8236
rect 155420 6866 155448 8230
rect 155500 7812 155552 7818
rect 155500 7754 155552 7760
rect 155276 6820 155356 6848
rect 155408 6860 155460 6866
rect 155224 6802 155276 6808
rect 155408 6802 155460 6808
rect 155224 6248 155276 6254
rect 155222 6216 155224 6225
rect 155276 6216 155278 6225
rect 155222 6151 155278 6160
rect 155316 6180 155368 6186
rect 154672 5228 154724 5234
rect 154672 5170 154724 5176
rect 154960 5222 155080 5250
rect 154684 5030 154712 5170
rect 154672 5024 154724 5030
rect 154672 4966 154724 4972
rect 154592 4678 154712 4706
rect 154580 4616 154632 4622
rect 154580 4558 154632 4564
rect 154486 3496 154542 3505
rect 154486 3431 154542 3440
rect 154396 3188 154448 3194
rect 154396 3130 154448 3136
rect 154500 3058 154528 3431
rect 154592 3194 154620 4558
rect 154684 4214 154712 4678
rect 154960 4672 154988 5222
rect 155236 5114 155264 6151
rect 155316 6122 155368 6128
rect 155328 5953 155356 6122
rect 155314 5944 155370 5953
rect 155314 5879 155370 5888
rect 155420 5642 155448 6802
rect 155512 6798 155540 7754
rect 155604 7546 155632 12854
rect 155696 12434 155724 13398
rect 155972 13326 156000 14010
rect 155960 13320 156012 13326
rect 155960 13262 156012 13268
rect 156064 12850 156092 14146
rect 156144 13796 156196 13802
rect 156144 13738 156196 13744
rect 156156 12986 156184 13738
rect 156708 13326 156736 14554
rect 156788 13388 156840 13394
rect 156788 13330 156840 13336
rect 156696 13320 156748 13326
rect 156696 13262 156748 13268
rect 156800 12986 156828 13330
rect 157444 13326 157472 14690
rect 157616 14000 157668 14006
rect 157616 13942 157668 13948
rect 157432 13320 157484 13326
rect 157432 13262 157484 13268
rect 156144 12980 156196 12986
rect 156144 12922 156196 12928
rect 156788 12980 156840 12986
rect 156788 12922 156840 12928
rect 156694 12880 156750 12889
rect 156052 12844 156104 12850
rect 156694 12815 156696 12824
rect 156052 12786 156104 12792
rect 156748 12815 156750 12824
rect 156696 12786 156748 12792
rect 155696 12406 155816 12434
rect 155684 11824 155736 11830
rect 155684 11766 155736 11772
rect 155696 11694 155724 11766
rect 155684 11688 155736 11694
rect 155684 11630 155736 11636
rect 155684 11552 155736 11558
rect 155684 11494 155736 11500
rect 155696 11354 155724 11494
rect 155684 11348 155736 11354
rect 155684 11290 155736 11296
rect 155684 10804 155736 10810
rect 155684 10746 155736 10752
rect 155592 7540 155644 7546
rect 155592 7482 155644 7488
rect 155696 7478 155724 10746
rect 155788 10062 155816 12406
rect 156326 12336 156382 12345
rect 155868 12300 155920 12306
rect 156326 12271 156382 12280
rect 155868 12242 155920 12248
rect 155880 11558 155908 12242
rect 156142 11792 156198 11801
rect 156142 11727 156144 11736
rect 156196 11727 156198 11736
rect 156144 11698 156196 11704
rect 156144 11620 156196 11626
rect 156144 11562 156196 11568
rect 155868 11552 155920 11558
rect 155868 11494 155920 11500
rect 155880 10470 155908 11494
rect 156052 11348 156104 11354
rect 156052 11290 156104 11296
rect 155960 11144 156012 11150
rect 155960 11086 156012 11092
rect 155868 10464 155920 10470
rect 155868 10406 155920 10412
rect 155776 10056 155828 10062
rect 155776 9998 155828 10004
rect 155880 9518 155908 10406
rect 155972 10062 156000 11086
rect 155960 10056 156012 10062
rect 155960 9998 156012 10004
rect 156064 9674 156092 11290
rect 156156 11082 156184 11562
rect 156236 11144 156288 11150
rect 156236 11086 156288 11092
rect 156144 11076 156196 11082
rect 156144 11018 156196 11024
rect 156144 10668 156196 10674
rect 156144 10610 156196 10616
rect 156156 10577 156184 10610
rect 156142 10568 156198 10577
rect 156142 10503 156198 10512
rect 156248 10198 156276 11086
rect 156236 10192 156288 10198
rect 156236 10134 156288 10140
rect 156064 9646 156276 9674
rect 156144 9580 156196 9586
rect 156144 9522 156196 9528
rect 155868 9512 155920 9518
rect 155868 9454 155920 9460
rect 156050 9344 156106 9353
rect 156050 9279 156106 9288
rect 155866 9208 155922 9217
rect 155866 9143 155922 9152
rect 155776 8424 155828 8430
rect 155776 8366 155828 8372
rect 155788 7954 155816 8366
rect 155880 8090 155908 9143
rect 155960 9036 156012 9042
rect 155960 8978 156012 8984
rect 155972 8634 156000 8978
rect 156064 8974 156092 9279
rect 156156 9081 156184 9522
rect 156248 9466 156276 9646
rect 156340 9586 156368 12271
rect 157064 12096 157116 12102
rect 157064 12038 157116 12044
rect 156512 11552 156564 11558
rect 156512 11494 156564 11500
rect 156420 11076 156472 11082
rect 156420 11018 156472 11024
rect 156328 9580 156380 9586
rect 156328 9522 156380 9528
rect 156248 9438 156368 9466
rect 156236 9376 156288 9382
rect 156236 9318 156288 9324
rect 156142 9072 156198 9081
rect 156142 9007 156198 9016
rect 156052 8968 156104 8974
rect 156052 8910 156104 8916
rect 156144 8968 156196 8974
rect 156144 8910 156196 8916
rect 155960 8628 156012 8634
rect 155960 8570 156012 8576
rect 156156 8362 156184 8910
rect 155960 8356 156012 8362
rect 155960 8298 156012 8304
rect 156144 8356 156196 8362
rect 156144 8298 156196 8304
rect 155868 8084 155920 8090
rect 155868 8026 155920 8032
rect 155776 7948 155828 7954
rect 155776 7890 155828 7896
rect 155788 7478 155816 7890
rect 155868 7744 155920 7750
rect 155866 7712 155868 7721
rect 155920 7712 155922 7721
rect 155866 7647 155922 7656
rect 155868 7540 155920 7546
rect 155868 7482 155920 7488
rect 155684 7472 155736 7478
rect 155684 7414 155736 7420
rect 155776 7472 155828 7478
rect 155776 7414 155828 7420
rect 155592 7404 155644 7410
rect 155592 7346 155644 7352
rect 155500 6792 155552 6798
rect 155500 6734 155552 6740
rect 155500 5704 155552 5710
rect 155498 5672 155500 5681
rect 155552 5672 155554 5681
rect 155408 5636 155460 5642
rect 155498 5607 155554 5616
rect 155408 5578 155460 5584
rect 154776 4644 154988 4672
rect 155144 5086 155264 5114
rect 155316 5092 155368 5098
rect 154672 4208 154724 4214
rect 154672 4150 154724 4156
rect 154672 4072 154724 4078
rect 154672 4014 154724 4020
rect 154684 3777 154712 4014
rect 154670 3768 154726 3777
rect 154670 3703 154726 3712
rect 154670 3496 154726 3505
rect 154670 3431 154672 3440
rect 154724 3431 154726 3440
rect 154672 3402 154724 3408
rect 154580 3188 154632 3194
rect 154580 3130 154632 3136
rect 154488 3052 154540 3058
rect 154488 2994 154540 3000
rect 154212 2848 154264 2854
rect 154212 2790 154264 2796
rect 154776 2774 154804 4644
rect 155144 4622 155172 5086
rect 155316 5034 155368 5040
rect 155132 4616 155184 4622
rect 155132 4558 155184 4564
rect 155224 4616 155276 4622
rect 155224 4558 155276 4564
rect 154948 4548 155000 4554
rect 154948 4490 155000 4496
rect 154960 4128 154988 4490
rect 155236 4321 155264 4558
rect 155328 4486 155356 5034
rect 155420 5030 155448 5578
rect 155498 5264 155554 5273
rect 155498 5199 155554 5208
rect 155512 5098 155540 5199
rect 155500 5092 155552 5098
rect 155500 5034 155552 5040
rect 155408 5024 155460 5030
rect 155408 4966 155460 4972
rect 155316 4480 155368 4486
rect 155316 4422 155368 4428
rect 155222 4312 155278 4321
rect 155222 4247 155278 4256
rect 155224 4140 155276 4146
rect 154960 4100 155224 4128
rect 155224 4082 155276 4088
rect 155130 4040 155186 4049
rect 155130 3975 155132 3984
rect 155184 3975 155186 3984
rect 155132 3946 155184 3952
rect 154948 3936 155000 3942
rect 154948 3878 155000 3884
rect 154960 2990 154988 3878
rect 155038 3768 155094 3777
rect 155038 3703 155094 3712
rect 155052 3466 155080 3703
rect 155132 3528 155184 3534
rect 155130 3496 155132 3505
rect 155184 3496 155186 3505
rect 155040 3460 155092 3466
rect 155130 3431 155186 3440
rect 155224 3460 155276 3466
rect 155040 3402 155092 3408
rect 155224 3402 155276 3408
rect 155236 3074 155264 3402
rect 155144 3058 155264 3074
rect 155132 3052 155264 3058
rect 155184 3046 155264 3052
rect 155408 3052 155460 3058
rect 155132 2994 155184 3000
rect 155408 2994 155460 3000
rect 154948 2984 155000 2990
rect 154948 2926 155000 2932
rect 154776 2746 154988 2774
rect 154302 2680 154358 2689
rect 154302 2615 154358 2624
rect 154120 2508 154172 2514
rect 154120 2450 154172 2456
rect 154316 2446 154344 2615
rect 154304 2440 154356 2446
rect 154304 2382 154356 2388
rect 154960 1766 154988 2746
rect 155132 2440 155184 2446
rect 155132 2382 155184 2388
rect 154948 1760 155000 1766
rect 154948 1702 155000 1708
rect 155144 1698 155172 2382
rect 155132 1692 155184 1698
rect 155132 1634 155184 1640
rect 155420 1222 155448 2994
rect 155604 2922 155632 7346
rect 155880 7290 155908 7482
rect 155972 7313 156000 8298
rect 156052 7880 156104 7886
rect 156052 7822 156104 7828
rect 156064 7410 156092 7822
rect 156144 7744 156196 7750
rect 156144 7686 156196 7692
rect 156052 7404 156104 7410
rect 156052 7346 156104 7352
rect 155684 7268 155736 7274
rect 155684 7210 155736 7216
rect 155788 7262 155908 7290
rect 155958 7304 156014 7313
rect 155696 3670 155724 7210
rect 155788 7206 155816 7262
rect 155958 7239 156014 7248
rect 155776 7200 155828 7206
rect 155776 7142 155828 7148
rect 155788 5710 155816 7142
rect 156052 6792 156104 6798
rect 156052 6734 156104 6740
rect 155960 6656 156012 6662
rect 155960 6598 156012 6604
rect 155868 6112 155920 6118
rect 155868 6054 155920 6060
rect 155776 5704 155828 5710
rect 155776 5646 155828 5652
rect 155788 5234 155816 5646
rect 155880 5642 155908 6054
rect 155972 5681 156000 6598
rect 155958 5672 156014 5681
rect 155868 5636 155920 5642
rect 155958 5607 156014 5616
rect 155868 5578 155920 5584
rect 155868 5364 155920 5370
rect 155868 5306 155920 5312
rect 155776 5228 155828 5234
rect 155776 5170 155828 5176
rect 155774 4040 155830 4049
rect 155774 3975 155830 3984
rect 155684 3664 155736 3670
rect 155684 3606 155736 3612
rect 155788 3534 155816 3975
rect 155776 3528 155828 3534
rect 155776 3470 155828 3476
rect 155592 2916 155644 2922
rect 155592 2858 155644 2864
rect 155776 2848 155828 2854
rect 155776 2790 155828 2796
rect 155788 2582 155816 2790
rect 155776 2576 155828 2582
rect 155776 2518 155828 2524
rect 155880 2446 155908 5306
rect 156064 4865 156092 6734
rect 156050 4856 156106 4865
rect 156050 4791 156106 4800
rect 156156 4622 156184 7686
rect 156248 7426 156276 9318
rect 156340 8974 156368 9438
rect 156328 8968 156380 8974
rect 156328 8910 156380 8916
rect 156340 7546 156368 8910
rect 156328 7540 156380 7546
rect 156328 7482 156380 7488
rect 156248 7398 156368 7426
rect 156236 7336 156288 7342
rect 156236 7278 156288 7284
rect 156144 4616 156196 4622
rect 156144 4558 156196 4564
rect 156052 4004 156104 4010
rect 156052 3946 156104 3952
rect 155960 2916 156012 2922
rect 155960 2858 156012 2864
rect 155972 2825 156000 2858
rect 155958 2816 156014 2825
rect 155958 2751 156014 2760
rect 155960 2576 156012 2582
rect 155960 2518 156012 2524
rect 155868 2440 155920 2446
rect 155868 2382 155920 2388
rect 155868 2304 155920 2310
rect 155868 2246 155920 2252
rect 155880 2009 155908 2246
rect 155866 2000 155922 2009
rect 155866 1935 155922 1944
rect 155972 1630 156000 2518
rect 156064 1834 156092 3946
rect 156248 2990 156276 7278
rect 156340 6202 156368 7398
rect 156432 6322 156460 11018
rect 156420 6316 156472 6322
rect 156420 6258 156472 6264
rect 156340 6174 156460 6202
rect 156328 6112 156380 6118
rect 156328 6054 156380 6060
rect 156340 2990 156368 6054
rect 156432 4146 156460 6174
rect 156524 4146 156552 11494
rect 157076 11257 157104 12038
rect 157628 11898 157656 13942
rect 158076 13932 158128 13938
rect 158076 13874 158128 13880
rect 158088 12986 158116 13874
rect 158729 13084 159037 13093
rect 158729 13082 158735 13084
rect 158791 13082 158815 13084
rect 158871 13082 158895 13084
rect 158951 13082 158975 13084
rect 159031 13082 159037 13084
rect 158791 13030 158793 13082
rect 158973 13030 158975 13082
rect 158729 13028 158735 13030
rect 158791 13028 158815 13030
rect 158871 13028 158895 13030
rect 158951 13028 158975 13030
rect 159031 13028 159037 13030
rect 158729 13019 159037 13028
rect 158076 12980 158128 12986
rect 158076 12922 158128 12928
rect 158352 12776 158404 12782
rect 158352 12718 158404 12724
rect 158168 12708 158220 12714
rect 158168 12650 158220 12656
rect 157616 11892 157668 11898
rect 157616 11834 157668 11840
rect 157062 11248 157118 11257
rect 157062 11183 157118 11192
rect 157432 11008 157484 11014
rect 156970 10976 157026 10985
rect 157432 10950 157484 10956
rect 156970 10911 157026 10920
rect 156984 10674 157012 10911
rect 156972 10668 157024 10674
rect 156972 10610 157024 10616
rect 157156 10464 157208 10470
rect 157156 10406 157208 10412
rect 156604 10056 156656 10062
rect 156604 9998 156656 10004
rect 156616 8344 156644 9998
rect 156878 9480 156934 9489
rect 156878 9415 156934 9424
rect 156972 9444 157024 9450
rect 156892 9110 156920 9415
rect 156972 9386 157024 9392
rect 156880 9104 156932 9110
rect 156880 9046 156932 9052
rect 156788 8968 156840 8974
rect 156708 8928 156788 8956
rect 156708 8673 156736 8928
rect 156788 8910 156840 8916
rect 156880 8832 156932 8838
rect 156880 8774 156932 8780
rect 156694 8664 156750 8673
rect 156694 8599 156750 8608
rect 156788 8628 156840 8634
rect 156788 8570 156840 8576
rect 156800 8498 156828 8570
rect 156788 8492 156840 8498
rect 156788 8434 156840 8440
rect 156616 8316 156736 8344
rect 156602 7984 156658 7993
rect 156602 7919 156658 7928
rect 156616 7886 156644 7919
rect 156604 7880 156656 7886
rect 156604 7822 156656 7828
rect 156708 7342 156736 8316
rect 156696 7336 156748 7342
rect 156696 7278 156748 7284
rect 156800 6866 156828 8434
rect 156788 6860 156840 6866
rect 156788 6802 156840 6808
rect 156800 6254 156828 6802
rect 156788 6248 156840 6254
rect 156788 6190 156840 6196
rect 156788 6112 156840 6118
rect 156694 6080 156750 6089
rect 156788 6054 156840 6060
rect 156694 6015 156750 6024
rect 156708 5846 156736 6015
rect 156800 5914 156828 6054
rect 156788 5908 156840 5914
rect 156788 5850 156840 5856
rect 156696 5840 156748 5846
rect 156696 5782 156748 5788
rect 156786 5400 156842 5409
rect 156786 5335 156788 5344
rect 156840 5335 156842 5344
rect 156788 5306 156840 5312
rect 156604 5228 156656 5234
rect 156604 5170 156656 5176
rect 156420 4140 156472 4146
rect 156420 4082 156472 4088
rect 156512 4140 156564 4146
rect 156512 4082 156564 4088
rect 156432 3942 156460 4082
rect 156420 3936 156472 3942
rect 156420 3878 156472 3884
rect 156236 2984 156288 2990
rect 156236 2926 156288 2932
rect 156328 2984 156380 2990
rect 156328 2926 156380 2932
rect 156432 2938 156460 3878
rect 156616 3194 156644 5170
rect 156892 4622 156920 8774
rect 156984 8634 157012 9386
rect 157064 9376 157116 9382
rect 157064 9318 157116 9324
rect 156972 8628 157024 8634
rect 156972 8570 157024 8576
rect 156970 8528 157026 8537
rect 156970 8463 156972 8472
rect 157024 8463 157026 8472
rect 156972 8434 157024 8440
rect 156970 7576 157026 7585
rect 156970 7511 157026 7520
rect 156984 7410 157012 7511
rect 156972 7404 157024 7410
rect 156972 7346 157024 7352
rect 156972 7200 157024 7206
rect 156972 7142 157024 7148
rect 156880 4616 156932 4622
rect 156880 4558 156932 4564
rect 156788 3936 156840 3942
rect 156786 3904 156788 3913
rect 156880 3936 156932 3942
rect 156840 3904 156842 3913
rect 156880 3878 156932 3884
rect 156786 3839 156842 3848
rect 156892 3738 156920 3878
rect 156880 3732 156932 3738
rect 156880 3674 156932 3680
rect 156984 3534 157012 7142
rect 157076 6798 157104 9318
rect 157064 6792 157116 6798
rect 157064 6734 157116 6740
rect 157064 6112 157116 6118
rect 157064 6054 157116 6060
rect 157076 5545 157104 6054
rect 157168 5710 157196 10406
rect 157340 8356 157392 8362
rect 157340 8298 157392 8304
rect 157246 7168 157302 7177
rect 157246 7103 157302 7112
rect 157260 5846 157288 7103
rect 157248 5840 157300 5846
rect 157248 5782 157300 5788
rect 157156 5704 157208 5710
rect 157156 5646 157208 5652
rect 157062 5536 157118 5545
rect 157062 5471 157118 5480
rect 157156 5364 157208 5370
rect 157156 5306 157208 5312
rect 157064 5024 157116 5030
rect 157064 4966 157116 4972
rect 156972 3528 157024 3534
rect 156972 3470 157024 3476
rect 156604 3188 156656 3194
rect 156604 3130 156656 3136
rect 157076 3058 157104 4966
rect 157064 3052 157116 3058
rect 157064 2994 157116 3000
rect 157168 2938 157196 5306
rect 157352 5234 157380 8298
rect 157444 8242 157472 10950
rect 157708 10124 157760 10130
rect 157708 10066 157760 10072
rect 157524 10056 157576 10062
rect 157522 10024 157524 10033
rect 157576 10024 157578 10033
rect 157522 9959 157578 9968
rect 157614 9752 157670 9761
rect 157614 9687 157670 9696
rect 157524 9376 157576 9382
rect 157524 9318 157576 9324
rect 157536 8362 157564 9318
rect 157524 8356 157576 8362
rect 157524 8298 157576 8304
rect 157444 8214 157564 8242
rect 157536 7750 157564 8214
rect 157524 7744 157576 7750
rect 157524 7686 157576 7692
rect 157628 7546 157656 9687
rect 157720 8974 157748 10066
rect 157892 9920 157944 9926
rect 157892 9862 157944 9868
rect 157800 9580 157852 9586
rect 157800 9522 157852 9528
rect 157812 9178 157840 9522
rect 157800 9172 157852 9178
rect 157800 9114 157852 9120
rect 157708 8968 157760 8974
rect 157708 8910 157760 8916
rect 157616 7540 157668 7546
rect 157616 7482 157668 7488
rect 157800 7404 157852 7410
rect 157800 7346 157852 7352
rect 157524 7268 157576 7274
rect 157524 7210 157576 7216
rect 157536 5710 157564 7210
rect 157708 6724 157760 6730
rect 157708 6666 157760 6672
rect 157616 6656 157668 6662
rect 157616 6598 157668 6604
rect 157524 5704 157576 5710
rect 157524 5646 157576 5652
rect 157340 5228 157392 5234
rect 157340 5170 157392 5176
rect 157248 5024 157300 5030
rect 157628 5001 157656 6598
rect 157248 4966 157300 4972
rect 157614 4992 157670 5001
rect 157260 4758 157288 4966
rect 157614 4927 157670 4936
rect 157248 4752 157300 4758
rect 157248 4694 157300 4700
rect 157248 4480 157300 4486
rect 157248 4422 157300 4428
rect 157260 4282 157288 4422
rect 157248 4276 157300 4282
rect 157248 4218 157300 4224
rect 157720 4146 157748 6666
rect 157812 6390 157840 7346
rect 157904 6798 157932 9862
rect 158076 9716 158128 9722
rect 158076 9658 158128 9664
rect 157984 9444 158036 9450
rect 157984 9386 158036 9392
rect 157892 6792 157944 6798
rect 157892 6734 157944 6740
rect 157800 6384 157852 6390
rect 157800 6326 157852 6332
rect 157996 4622 158024 9386
rect 158088 8498 158116 9658
rect 158076 8492 158128 8498
rect 158076 8434 158128 8440
rect 158076 8356 158128 8362
rect 158076 8298 158128 8304
rect 157984 4616 158036 4622
rect 157984 4558 158036 4564
rect 157708 4140 157760 4146
rect 157708 4082 157760 4088
rect 157616 3528 157668 3534
rect 157616 3470 157668 3476
rect 157432 3392 157484 3398
rect 157628 3369 157656 3470
rect 157432 3334 157484 3340
rect 157614 3360 157670 3369
rect 156432 2910 156552 2938
rect 156524 2854 156552 2910
rect 156984 2910 157196 2938
rect 156420 2848 156472 2854
rect 156420 2790 156472 2796
rect 156512 2848 156564 2854
rect 156512 2790 156564 2796
rect 156052 1828 156104 1834
rect 156052 1770 156104 1776
rect 155960 1624 156012 1630
rect 155960 1566 156012 1572
rect 155408 1216 155460 1222
rect 153750 1184 153806 1193
rect 155408 1158 155460 1164
rect 153750 1119 153806 1128
rect 151176 1080 151228 1086
rect 145746 1048 145802 1057
rect 113548 1012 113600 1018
rect 113548 954 113600 960
rect 138112 1012 138164 1018
rect 156432 1057 156460 2790
rect 156604 2304 156656 2310
rect 156604 2246 156656 2252
rect 156616 2106 156644 2246
rect 156604 2100 156656 2106
rect 156604 2042 156656 2048
rect 156984 1562 157012 2910
rect 157156 2848 157208 2854
rect 157156 2790 157208 2796
rect 157168 2514 157196 2790
rect 157444 2582 157472 3334
rect 157614 3295 157670 3304
rect 158088 3097 158116 8298
rect 158180 6322 158208 12650
rect 158364 12434 158392 12718
rect 158364 12406 159404 12434
rect 159180 12232 159232 12238
rect 159180 12174 159232 12180
rect 158729 11996 159037 12005
rect 158729 11994 158735 11996
rect 158791 11994 158815 11996
rect 158871 11994 158895 11996
rect 158951 11994 158975 11996
rect 159031 11994 159037 11996
rect 158791 11942 158793 11994
rect 158973 11942 158975 11994
rect 158729 11940 158735 11942
rect 158791 11940 158815 11942
rect 158871 11940 158895 11942
rect 158951 11940 158975 11942
rect 159031 11940 159037 11942
rect 158729 11931 159037 11940
rect 158260 11552 158312 11558
rect 158260 11494 158312 11500
rect 158272 10810 158300 11494
rect 158352 11280 158404 11286
rect 158352 11222 158404 11228
rect 158260 10804 158312 10810
rect 158260 10746 158312 10752
rect 158272 9722 158300 10746
rect 158260 9716 158312 9722
rect 158260 9658 158312 9664
rect 158260 8356 158312 8362
rect 158260 8298 158312 8304
rect 158272 7993 158300 8298
rect 158258 7984 158314 7993
rect 158258 7919 158314 7928
rect 158260 7744 158312 7750
rect 158260 7686 158312 7692
rect 158168 6316 158220 6322
rect 158168 6258 158220 6264
rect 158272 6202 158300 7686
rect 158180 6174 158300 6202
rect 158180 3194 158208 6174
rect 158260 5772 158312 5778
rect 158260 5714 158312 5720
rect 158272 4146 158300 5714
rect 158260 4140 158312 4146
rect 158260 4082 158312 4088
rect 158168 3188 158220 3194
rect 158168 3130 158220 3136
rect 158074 3088 158130 3097
rect 158074 3023 158130 3032
rect 158364 2774 158392 11222
rect 158628 11144 158680 11150
rect 158628 11086 158680 11092
rect 158444 10532 158496 10538
rect 158444 10474 158496 10480
rect 158456 6390 158484 10474
rect 158536 8900 158588 8906
rect 158536 8842 158588 8848
rect 158444 6384 158496 6390
rect 158444 6326 158496 6332
rect 158548 5234 158576 8842
rect 158640 5574 158668 11086
rect 158729 10908 159037 10917
rect 158729 10906 158735 10908
rect 158791 10906 158815 10908
rect 158871 10906 158895 10908
rect 158951 10906 158975 10908
rect 159031 10906 159037 10908
rect 158791 10854 158793 10906
rect 158973 10854 158975 10906
rect 158729 10852 158735 10854
rect 158791 10852 158815 10854
rect 158871 10852 158895 10854
rect 158951 10852 158975 10854
rect 159031 10852 159037 10854
rect 158729 10843 159037 10852
rect 159088 10668 159140 10674
rect 159088 10610 159140 10616
rect 158729 9820 159037 9829
rect 158729 9818 158735 9820
rect 158791 9818 158815 9820
rect 158871 9818 158895 9820
rect 158951 9818 158975 9820
rect 159031 9818 159037 9820
rect 158791 9766 158793 9818
rect 158973 9766 158975 9818
rect 158729 9764 158735 9766
rect 158791 9764 158815 9766
rect 158871 9764 158895 9766
rect 158951 9764 158975 9766
rect 159031 9764 159037 9766
rect 158729 9755 159037 9764
rect 158729 8732 159037 8741
rect 158729 8730 158735 8732
rect 158791 8730 158815 8732
rect 158871 8730 158895 8732
rect 158951 8730 158975 8732
rect 159031 8730 159037 8732
rect 158791 8678 158793 8730
rect 158973 8678 158975 8730
rect 158729 8676 158735 8678
rect 158791 8676 158815 8678
rect 158871 8676 158895 8678
rect 158951 8676 158975 8678
rect 159031 8676 159037 8678
rect 158729 8667 159037 8676
rect 158729 7644 159037 7653
rect 158729 7642 158735 7644
rect 158791 7642 158815 7644
rect 158871 7642 158895 7644
rect 158951 7642 158975 7644
rect 159031 7642 159037 7644
rect 158791 7590 158793 7642
rect 158973 7590 158975 7642
rect 158729 7588 158735 7590
rect 158791 7588 158815 7590
rect 158871 7588 158895 7590
rect 158951 7588 158975 7590
rect 159031 7588 159037 7590
rect 158729 7579 159037 7588
rect 158729 6556 159037 6565
rect 158729 6554 158735 6556
rect 158791 6554 158815 6556
rect 158871 6554 158895 6556
rect 158951 6554 158975 6556
rect 159031 6554 159037 6556
rect 158791 6502 158793 6554
rect 158973 6502 158975 6554
rect 158729 6500 158735 6502
rect 158791 6500 158815 6502
rect 158871 6500 158895 6502
rect 158951 6500 158975 6502
rect 159031 6500 159037 6502
rect 158729 6491 159037 6500
rect 158628 5568 158680 5574
rect 158628 5510 158680 5516
rect 158729 5468 159037 5477
rect 158729 5466 158735 5468
rect 158791 5466 158815 5468
rect 158871 5466 158895 5468
rect 158951 5466 158975 5468
rect 159031 5466 159037 5468
rect 158791 5414 158793 5466
rect 158973 5414 158975 5466
rect 158729 5412 158735 5414
rect 158791 5412 158815 5414
rect 158871 5412 158895 5414
rect 158951 5412 158975 5414
rect 159031 5412 159037 5414
rect 158729 5403 159037 5412
rect 158536 5228 158588 5234
rect 158536 5170 158588 5176
rect 158729 4380 159037 4389
rect 158729 4378 158735 4380
rect 158791 4378 158815 4380
rect 158871 4378 158895 4380
rect 158951 4378 158975 4380
rect 159031 4378 159037 4380
rect 158791 4326 158793 4378
rect 158973 4326 158975 4378
rect 158729 4324 158735 4326
rect 158791 4324 158815 4326
rect 158871 4324 158895 4326
rect 158951 4324 158975 4326
rect 159031 4324 159037 4326
rect 158729 4315 159037 4324
rect 158729 3292 159037 3301
rect 158729 3290 158735 3292
rect 158791 3290 158815 3292
rect 158871 3290 158895 3292
rect 158951 3290 158975 3292
rect 159031 3290 159037 3292
rect 158791 3238 158793 3290
rect 158973 3238 158975 3290
rect 158729 3236 158735 3238
rect 158791 3236 158815 3238
rect 158871 3236 158895 3238
rect 158951 3236 158975 3238
rect 159031 3236 159037 3238
rect 158729 3227 159037 3236
rect 158180 2746 158392 2774
rect 157432 2576 157484 2582
rect 157432 2518 157484 2524
rect 157156 2508 157208 2514
rect 157156 2450 157208 2456
rect 157800 2304 157852 2310
rect 158180 2281 158208 2746
rect 159100 2650 159128 10610
rect 159192 5302 159220 12174
rect 159270 10296 159326 10305
rect 159270 10231 159326 10240
rect 159180 5296 159232 5302
rect 159180 5238 159232 5244
rect 159284 4826 159312 10231
rect 159272 4820 159324 4826
rect 159272 4762 159324 4768
rect 159376 4690 159404 12406
rect 159456 11348 159508 11354
rect 159456 11290 159508 11296
rect 159364 4684 159416 4690
rect 159364 4626 159416 4632
rect 159468 2774 159496 11290
rect 159192 2746 159496 2774
rect 159088 2644 159140 2650
rect 159088 2586 159140 2592
rect 157800 2246 157852 2252
rect 158166 2272 158222 2281
rect 157812 2145 157840 2246
rect 158166 2207 158222 2216
rect 158729 2204 159037 2213
rect 158729 2202 158735 2204
rect 158791 2202 158815 2204
rect 158871 2202 158895 2204
rect 158951 2202 158975 2204
rect 159031 2202 159037 2204
rect 158791 2150 158793 2202
rect 158973 2150 158975 2202
rect 158729 2148 158735 2150
rect 158791 2148 158815 2150
rect 158871 2148 158895 2150
rect 158951 2148 158975 2150
rect 159031 2148 159037 2150
rect 157798 2136 157854 2145
rect 158729 2139 159037 2148
rect 157798 2071 157854 2080
rect 159192 1970 159220 2746
rect 159180 1964 159232 1970
rect 159180 1906 159232 1912
rect 156972 1556 157024 1562
rect 156972 1498 157024 1504
rect 151176 1022 151228 1028
rect 156418 1048 156474 1057
rect 145746 983 145802 992
rect 156418 983 156474 992
rect 138112 954 138164 960
<< via2 >>
rect 4066 13812 4068 13832
rect 4068 13812 4120 13832
rect 4120 13812 4122 13832
rect 4066 13776 4122 13812
rect 10230 13268 10232 13288
rect 10232 13268 10284 13288
rect 10284 13268 10286 13288
rect 10230 13232 10286 13268
rect 9862 12180 9864 12200
rect 9864 12180 9916 12200
rect 9916 12180 9918 12200
rect 1582 9832 1638 9888
rect 9862 12144 9918 12180
rect 1582 5888 1638 5944
rect 10322 6160 10378 6216
rect 10690 11600 10746 11656
rect 10506 11212 10562 11248
rect 10506 11192 10508 11212
rect 10508 11192 10560 11212
rect 10560 11192 10562 11212
rect 11886 11756 11942 11792
rect 11886 11736 11888 11756
rect 11888 11736 11940 11756
rect 11940 11736 11942 11756
rect 12070 12280 12126 12336
rect 12438 12280 12494 12336
rect 12438 10512 12494 10568
rect 12898 11636 12900 11656
rect 12900 11636 12952 11656
rect 12952 11636 12954 11656
rect 12898 11600 12954 11636
rect 13358 10512 13414 10568
rect 14830 12180 14832 12200
rect 14832 12180 14884 12200
rect 14884 12180 14886 12200
rect 14830 12144 14886 12180
rect 14094 11192 14150 11248
rect 14278 9036 14334 9072
rect 14278 9016 14280 9036
rect 14280 9016 14332 9036
rect 14332 9016 14334 9036
rect 16394 13232 16450 13288
rect 15934 11736 15990 11792
rect 17958 12144 18014 12200
rect 17222 10648 17278 10704
rect 16302 5364 16358 5400
rect 16302 5344 16304 5364
rect 16304 5344 16356 5364
rect 16356 5344 16358 5364
rect 16946 9036 17002 9072
rect 16946 9016 16948 9036
rect 16948 9016 17000 9036
rect 17000 9016 17002 9036
rect 16762 8372 16764 8392
rect 16764 8372 16816 8392
rect 16816 8372 16818 8392
rect 16762 8336 16818 8372
rect 17314 5344 17370 5400
rect 19338 11056 19394 11112
rect 19430 8336 19486 8392
rect 20678 13626 20734 13628
rect 20758 13626 20814 13628
rect 20838 13626 20894 13628
rect 20918 13626 20974 13628
rect 20678 13574 20724 13626
rect 20724 13574 20734 13626
rect 20758 13574 20788 13626
rect 20788 13574 20800 13626
rect 20800 13574 20814 13626
rect 20838 13574 20852 13626
rect 20852 13574 20864 13626
rect 20864 13574 20894 13626
rect 20918 13574 20928 13626
rect 20928 13574 20974 13626
rect 20678 13572 20734 13574
rect 20758 13572 20814 13574
rect 20838 13572 20894 13574
rect 20918 13572 20974 13574
rect 21362 13096 21418 13152
rect 20678 12538 20734 12540
rect 20758 12538 20814 12540
rect 20838 12538 20894 12540
rect 20918 12538 20974 12540
rect 20678 12486 20724 12538
rect 20724 12486 20734 12538
rect 20758 12486 20788 12538
rect 20788 12486 20800 12538
rect 20800 12486 20814 12538
rect 20838 12486 20852 12538
rect 20852 12486 20864 12538
rect 20864 12486 20894 12538
rect 20918 12486 20928 12538
rect 20928 12486 20974 12538
rect 20678 12484 20734 12486
rect 20758 12484 20814 12486
rect 20838 12484 20894 12486
rect 20918 12484 20974 12486
rect 21546 12688 21602 12744
rect 20626 11600 20682 11656
rect 19798 9444 19854 9480
rect 19798 9424 19800 9444
rect 19800 9424 19852 9444
rect 19852 9424 19854 9444
rect 20678 11450 20734 11452
rect 20758 11450 20814 11452
rect 20838 11450 20894 11452
rect 20918 11450 20974 11452
rect 20678 11398 20724 11450
rect 20724 11398 20734 11450
rect 20758 11398 20788 11450
rect 20788 11398 20800 11450
rect 20800 11398 20814 11450
rect 20838 11398 20852 11450
rect 20852 11398 20864 11450
rect 20864 11398 20894 11450
rect 20918 11398 20928 11450
rect 20928 11398 20974 11450
rect 20678 11396 20734 11398
rect 20758 11396 20814 11398
rect 20838 11396 20894 11398
rect 20918 11396 20974 11398
rect 20678 10362 20734 10364
rect 20758 10362 20814 10364
rect 20838 10362 20894 10364
rect 20918 10362 20974 10364
rect 20678 10310 20724 10362
rect 20724 10310 20734 10362
rect 20758 10310 20788 10362
rect 20788 10310 20800 10362
rect 20800 10310 20814 10362
rect 20838 10310 20852 10362
rect 20852 10310 20864 10362
rect 20864 10310 20894 10362
rect 20918 10310 20928 10362
rect 20928 10310 20974 10362
rect 20678 10308 20734 10310
rect 20758 10308 20814 10310
rect 20838 10308 20894 10310
rect 20918 10308 20974 10310
rect 20678 9274 20734 9276
rect 20758 9274 20814 9276
rect 20838 9274 20894 9276
rect 20918 9274 20974 9276
rect 20678 9222 20724 9274
rect 20724 9222 20734 9274
rect 20758 9222 20788 9274
rect 20788 9222 20800 9274
rect 20800 9222 20814 9274
rect 20838 9222 20852 9274
rect 20852 9222 20864 9274
rect 20864 9222 20894 9274
rect 20918 9222 20928 9274
rect 20928 9222 20974 9274
rect 20678 9220 20734 9222
rect 20758 9220 20814 9222
rect 20838 9220 20894 9222
rect 20918 9220 20974 9222
rect 20678 8186 20734 8188
rect 20758 8186 20814 8188
rect 20838 8186 20894 8188
rect 20918 8186 20974 8188
rect 20678 8134 20724 8186
rect 20724 8134 20734 8186
rect 20758 8134 20788 8186
rect 20788 8134 20800 8186
rect 20800 8134 20814 8186
rect 20838 8134 20852 8186
rect 20852 8134 20864 8186
rect 20864 8134 20894 8186
rect 20918 8134 20928 8186
rect 20928 8134 20974 8186
rect 20678 8132 20734 8134
rect 20758 8132 20814 8134
rect 20838 8132 20894 8134
rect 20918 8132 20974 8134
rect 20678 7098 20734 7100
rect 20758 7098 20814 7100
rect 20838 7098 20894 7100
rect 20918 7098 20974 7100
rect 20678 7046 20724 7098
rect 20724 7046 20734 7098
rect 20758 7046 20788 7098
rect 20788 7046 20800 7098
rect 20800 7046 20814 7098
rect 20838 7046 20852 7098
rect 20852 7046 20864 7098
rect 20864 7046 20894 7098
rect 20918 7046 20928 7098
rect 20928 7046 20974 7098
rect 20678 7044 20734 7046
rect 20758 7044 20814 7046
rect 20838 7044 20894 7046
rect 20918 7044 20974 7046
rect 20678 6010 20734 6012
rect 20758 6010 20814 6012
rect 20838 6010 20894 6012
rect 20918 6010 20974 6012
rect 20678 5958 20724 6010
rect 20724 5958 20734 6010
rect 20758 5958 20788 6010
rect 20788 5958 20800 6010
rect 20800 5958 20814 6010
rect 20838 5958 20852 6010
rect 20852 5958 20864 6010
rect 20864 5958 20894 6010
rect 20918 5958 20928 6010
rect 20928 5958 20974 6010
rect 20678 5956 20734 5958
rect 20758 5956 20814 5958
rect 20838 5956 20894 5958
rect 20918 5956 20974 5958
rect 20678 4922 20734 4924
rect 20758 4922 20814 4924
rect 20838 4922 20894 4924
rect 20918 4922 20974 4924
rect 20678 4870 20724 4922
rect 20724 4870 20734 4922
rect 20758 4870 20788 4922
rect 20788 4870 20800 4922
rect 20800 4870 20814 4922
rect 20838 4870 20852 4922
rect 20852 4870 20864 4922
rect 20864 4870 20894 4922
rect 20918 4870 20928 4922
rect 20928 4870 20974 4922
rect 20678 4868 20734 4870
rect 20758 4868 20814 4870
rect 20838 4868 20894 4870
rect 20918 4868 20974 4870
rect 20678 3834 20734 3836
rect 20758 3834 20814 3836
rect 20838 3834 20894 3836
rect 20918 3834 20974 3836
rect 20678 3782 20724 3834
rect 20724 3782 20734 3834
rect 20758 3782 20788 3834
rect 20788 3782 20800 3834
rect 20800 3782 20814 3834
rect 20838 3782 20852 3834
rect 20852 3782 20864 3834
rect 20864 3782 20894 3834
rect 20918 3782 20928 3834
rect 20928 3782 20974 3834
rect 20678 3780 20734 3782
rect 20758 3780 20814 3782
rect 20838 3780 20894 3782
rect 20918 3780 20974 3782
rect 20534 3068 20536 3088
rect 20536 3068 20588 3088
rect 20588 3068 20590 3088
rect 20534 3032 20590 3068
rect 20678 2746 20734 2748
rect 20758 2746 20814 2748
rect 20838 2746 20894 2748
rect 20918 2746 20974 2748
rect 20678 2694 20724 2746
rect 20724 2694 20734 2746
rect 20758 2694 20788 2746
rect 20788 2694 20800 2746
rect 20800 2694 20814 2746
rect 20838 2694 20852 2746
rect 20852 2694 20864 2746
rect 20864 2694 20894 2746
rect 20918 2694 20928 2746
rect 20928 2694 20974 2746
rect 20678 2692 20734 2694
rect 20758 2692 20814 2694
rect 20838 2692 20894 2694
rect 20918 2692 20974 2694
rect 22742 12844 22798 12880
rect 22742 12824 22744 12844
rect 22744 12824 22796 12844
rect 22796 12824 22798 12844
rect 22466 11600 22522 11656
rect 21914 8472 21970 8528
rect 22098 5616 22154 5672
rect 24030 12708 24086 12744
rect 24030 12688 24032 12708
rect 24032 12688 24084 12708
rect 24084 12688 24086 12708
rect 26238 12688 26294 12744
rect 26882 10920 26938 10976
rect 24766 3032 24822 3088
rect 27802 10648 27858 10704
rect 27066 8356 27122 8392
rect 27066 8336 27068 8356
rect 27068 8336 27120 8356
rect 27120 8336 27122 8356
rect 27710 8492 27766 8528
rect 27710 8472 27712 8492
rect 27712 8472 27764 8492
rect 27764 8472 27766 8492
rect 27986 13096 28042 13152
rect 28906 11056 28962 11112
rect 28630 9424 28686 9480
rect 28170 8372 28172 8392
rect 28172 8372 28224 8392
rect 28224 8372 28226 8392
rect 28170 8336 28226 8372
rect 29734 12708 29790 12744
rect 29734 12688 29736 12708
rect 29736 12688 29788 12708
rect 29788 12688 29790 12708
rect 30102 13232 30158 13288
rect 30654 12824 30710 12880
rect 30378 10920 30434 10976
rect 29366 6180 29422 6216
rect 29366 6160 29368 6180
rect 29368 6160 29420 6180
rect 29420 6160 29422 6180
rect 30378 5652 30380 5672
rect 30380 5652 30432 5672
rect 30432 5652 30434 5672
rect 30378 5616 30434 5652
rect 31758 13232 31814 13288
rect 32034 9696 32090 9752
rect 34794 11620 34850 11656
rect 34794 11600 34796 11620
rect 34796 11600 34848 11620
rect 34848 11600 34850 11620
rect 34426 10548 34428 10568
rect 34428 10548 34480 10568
rect 34480 10548 34482 10568
rect 34426 10512 34482 10548
rect 37186 9696 37242 9752
rect 39762 8880 39818 8936
rect 40222 12280 40278 12336
rect 40400 13082 40456 13084
rect 40480 13082 40536 13084
rect 40560 13082 40616 13084
rect 40640 13082 40696 13084
rect 40400 13030 40446 13082
rect 40446 13030 40456 13082
rect 40480 13030 40510 13082
rect 40510 13030 40522 13082
rect 40522 13030 40536 13082
rect 40560 13030 40574 13082
rect 40574 13030 40586 13082
rect 40586 13030 40616 13082
rect 40640 13030 40650 13082
rect 40650 13030 40696 13082
rect 40400 13028 40456 13030
rect 40480 13028 40536 13030
rect 40560 13028 40616 13030
rect 40640 13028 40696 13030
rect 40400 11994 40456 11996
rect 40480 11994 40536 11996
rect 40560 11994 40616 11996
rect 40640 11994 40696 11996
rect 40400 11942 40446 11994
rect 40446 11942 40456 11994
rect 40480 11942 40510 11994
rect 40510 11942 40522 11994
rect 40522 11942 40536 11994
rect 40560 11942 40574 11994
rect 40574 11942 40586 11994
rect 40586 11942 40616 11994
rect 40640 11942 40650 11994
rect 40650 11942 40696 11994
rect 40400 11940 40456 11942
rect 40480 11940 40536 11942
rect 40560 11940 40616 11942
rect 40640 11940 40696 11942
rect 40866 12280 40922 12336
rect 40400 10906 40456 10908
rect 40480 10906 40536 10908
rect 40560 10906 40616 10908
rect 40640 10906 40696 10908
rect 40400 10854 40446 10906
rect 40446 10854 40456 10906
rect 40480 10854 40510 10906
rect 40510 10854 40522 10906
rect 40522 10854 40536 10906
rect 40560 10854 40574 10906
rect 40574 10854 40586 10906
rect 40586 10854 40616 10906
rect 40640 10854 40650 10906
rect 40650 10854 40696 10906
rect 40400 10852 40456 10854
rect 40480 10852 40536 10854
rect 40560 10852 40616 10854
rect 40640 10852 40696 10854
rect 40400 9818 40456 9820
rect 40480 9818 40536 9820
rect 40560 9818 40616 9820
rect 40640 9818 40696 9820
rect 40400 9766 40446 9818
rect 40446 9766 40456 9818
rect 40480 9766 40510 9818
rect 40510 9766 40522 9818
rect 40522 9766 40536 9818
rect 40560 9766 40574 9818
rect 40574 9766 40586 9818
rect 40586 9766 40616 9818
rect 40640 9766 40650 9818
rect 40650 9766 40696 9818
rect 40400 9764 40456 9766
rect 40480 9764 40536 9766
rect 40560 9764 40616 9766
rect 40640 9764 40696 9766
rect 40400 8730 40456 8732
rect 40480 8730 40536 8732
rect 40560 8730 40616 8732
rect 40640 8730 40696 8732
rect 40400 8678 40446 8730
rect 40446 8678 40456 8730
rect 40480 8678 40510 8730
rect 40510 8678 40522 8730
rect 40522 8678 40536 8730
rect 40560 8678 40574 8730
rect 40574 8678 40586 8730
rect 40586 8678 40616 8730
rect 40640 8678 40650 8730
rect 40650 8678 40696 8730
rect 40400 8676 40456 8678
rect 40480 8676 40536 8678
rect 40560 8676 40616 8678
rect 40640 8676 40696 8678
rect 40400 7642 40456 7644
rect 40480 7642 40536 7644
rect 40560 7642 40616 7644
rect 40640 7642 40696 7644
rect 40400 7590 40446 7642
rect 40446 7590 40456 7642
rect 40480 7590 40510 7642
rect 40510 7590 40522 7642
rect 40522 7590 40536 7642
rect 40560 7590 40574 7642
rect 40574 7590 40586 7642
rect 40586 7590 40616 7642
rect 40640 7590 40650 7642
rect 40650 7590 40696 7642
rect 40400 7588 40456 7590
rect 40480 7588 40536 7590
rect 40560 7588 40616 7590
rect 40640 7588 40696 7590
rect 40400 6554 40456 6556
rect 40480 6554 40536 6556
rect 40560 6554 40616 6556
rect 40640 6554 40696 6556
rect 40400 6502 40446 6554
rect 40446 6502 40456 6554
rect 40480 6502 40510 6554
rect 40510 6502 40522 6554
rect 40522 6502 40536 6554
rect 40560 6502 40574 6554
rect 40574 6502 40586 6554
rect 40586 6502 40616 6554
rect 40640 6502 40650 6554
rect 40650 6502 40696 6554
rect 40400 6500 40456 6502
rect 40480 6500 40536 6502
rect 40560 6500 40616 6502
rect 40640 6500 40696 6502
rect 41050 8472 41106 8528
rect 41234 9016 41290 9072
rect 40400 5466 40456 5468
rect 40480 5466 40536 5468
rect 40560 5466 40616 5468
rect 40640 5466 40696 5468
rect 40400 5414 40446 5466
rect 40446 5414 40456 5466
rect 40480 5414 40510 5466
rect 40510 5414 40522 5466
rect 40522 5414 40536 5466
rect 40560 5414 40574 5466
rect 40574 5414 40586 5466
rect 40586 5414 40616 5466
rect 40640 5414 40650 5466
rect 40650 5414 40696 5466
rect 40400 5412 40456 5414
rect 40480 5412 40536 5414
rect 40560 5412 40616 5414
rect 40640 5412 40696 5414
rect 40400 4378 40456 4380
rect 40480 4378 40536 4380
rect 40560 4378 40616 4380
rect 40640 4378 40696 4380
rect 40400 4326 40446 4378
rect 40446 4326 40456 4378
rect 40480 4326 40510 4378
rect 40510 4326 40522 4378
rect 40522 4326 40536 4378
rect 40560 4326 40574 4378
rect 40574 4326 40586 4378
rect 40586 4326 40616 4378
rect 40640 4326 40650 4378
rect 40650 4326 40696 4378
rect 40400 4324 40456 4326
rect 40480 4324 40536 4326
rect 40560 4324 40616 4326
rect 40640 4324 40696 4326
rect 40400 3290 40456 3292
rect 40480 3290 40536 3292
rect 40560 3290 40616 3292
rect 40640 3290 40696 3292
rect 40400 3238 40446 3290
rect 40446 3238 40456 3290
rect 40480 3238 40510 3290
rect 40510 3238 40522 3290
rect 40522 3238 40536 3290
rect 40560 3238 40574 3290
rect 40574 3238 40586 3290
rect 40586 3238 40616 3290
rect 40640 3238 40650 3290
rect 40650 3238 40696 3290
rect 40400 3236 40456 3238
rect 40480 3236 40536 3238
rect 40560 3236 40616 3238
rect 40640 3236 40696 3238
rect 41694 12688 41750 12744
rect 42154 12316 42156 12336
rect 42156 12316 42208 12336
rect 42208 12316 42210 12336
rect 42154 12280 42210 12316
rect 42062 11328 42118 11384
rect 41602 8880 41658 8936
rect 42062 9288 42118 9344
rect 42614 11464 42670 11520
rect 43074 11464 43130 11520
rect 43994 13368 44050 13424
rect 45558 12436 45614 12472
rect 45558 12416 45560 12436
rect 45560 12416 45612 12436
rect 45612 12416 45614 12436
rect 45466 12180 45468 12200
rect 45468 12180 45520 12200
rect 45520 12180 45522 12200
rect 45466 12144 45522 12180
rect 45374 11328 45430 11384
rect 44730 8492 44786 8528
rect 44730 8472 44732 8492
rect 44732 8472 44784 8492
rect 44784 8472 44786 8492
rect 46294 12688 46350 12744
rect 46938 12416 46994 12472
rect 46754 12280 46810 12336
rect 46294 9324 46296 9344
rect 46296 9324 46348 9344
rect 46348 9324 46350 9344
rect 46294 9288 46350 9324
rect 47674 9288 47730 9344
rect 48778 11872 48834 11928
rect 47950 9016 48006 9072
rect 48778 10376 48834 10432
rect 48870 8492 48926 8528
rect 48870 8472 48872 8492
rect 48872 8472 48924 8492
rect 48924 8472 48926 8492
rect 49790 13404 49792 13424
rect 49792 13404 49844 13424
rect 49844 13404 49846 13424
rect 49790 13368 49846 13404
rect 49146 10920 49202 10976
rect 49146 10240 49202 10296
rect 50158 10784 50214 10840
rect 50710 12824 50766 12880
rect 50894 12960 50950 13016
rect 50894 12280 50950 12336
rect 51170 12960 51226 13016
rect 50710 11464 50766 11520
rect 51170 10920 51226 10976
rect 49606 3340 49608 3360
rect 49608 3340 49660 3360
rect 49660 3340 49662 3360
rect 49606 3304 49662 3340
rect 51630 11192 51686 11248
rect 51538 10104 51594 10160
rect 52182 10104 52238 10160
rect 52550 11500 52552 11520
rect 52552 11500 52604 11520
rect 52604 11500 52606 11520
rect 52550 11464 52606 11500
rect 52826 11892 52882 11928
rect 52826 11872 52828 11892
rect 52828 11872 52880 11892
rect 52880 11872 52882 11892
rect 52550 10648 52606 10704
rect 53102 10648 53158 10704
rect 53930 11600 53986 11656
rect 53838 10784 53894 10840
rect 54390 10124 54446 10160
rect 54390 10104 54392 10124
rect 54392 10104 54444 10124
rect 54444 10104 54446 10124
rect 54206 9968 54262 10024
rect 55126 12144 55182 12200
rect 54114 9832 54170 9888
rect 55402 13096 55458 13152
rect 56046 12844 56102 12880
rect 56046 12824 56048 12844
rect 56048 12824 56100 12844
rect 56100 12824 56102 12844
rect 55954 12280 56010 12336
rect 55954 10140 55956 10160
rect 55956 10140 56008 10160
rect 56008 10140 56010 10160
rect 55954 10104 56010 10140
rect 56322 13232 56378 13288
rect 56230 9580 56286 9616
rect 56230 9560 56232 9580
rect 56232 9560 56284 9580
rect 56284 9560 56286 9580
rect 56690 13268 56692 13288
rect 56692 13268 56744 13288
rect 56744 13268 56746 13288
rect 56690 13232 56746 13268
rect 56506 10376 56562 10432
rect 53562 3340 53564 3360
rect 53564 3340 53616 3360
rect 53616 3340 53618 3360
rect 53562 3304 53618 3340
rect 57150 12300 57206 12336
rect 57150 12280 57152 12300
rect 57152 12280 57204 12300
rect 57204 12280 57206 12300
rect 57518 10240 57574 10296
rect 57058 9968 57114 10024
rect 57150 9596 57152 9616
rect 57152 9596 57204 9616
rect 57204 9596 57206 9616
rect 57150 9560 57206 9596
rect 57794 9832 57850 9888
rect 58346 10784 58402 10840
rect 58622 12960 58678 13016
rect 58622 11192 58678 11248
rect 58806 12280 58862 12336
rect 59450 13368 59506 13424
rect 58990 10104 59046 10160
rect 60123 13626 60179 13628
rect 60203 13626 60259 13628
rect 60283 13626 60339 13628
rect 60363 13626 60419 13628
rect 60123 13574 60169 13626
rect 60169 13574 60179 13626
rect 60203 13574 60233 13626
rect 60233 13574 60245 13626
rect 60245 13574 60259 13626
rect 60283 13574 60297 13626
rect 60297 13574 60309 13626
rect 60309 13574 60339 13626
rect 60363 13574 60373 13626
rect 60373 13574 60419 13626
rect 60123 13572 60179 13574
rect 60203 13572 60259 13574
rect 60283 13572 60339 13574
rect 60363 13572 60419 13574
rect 60370 13252 60426 13288
rect 60370 13232 60372 13252
rect 60372 13232 60424 13252
rect 60424 13232 60426 13252
rect 60123 12538 60179 12540
rect 60203 12538 60259 12540
rect 60283 12538 60339 12540
rect 60363 12538 60419 12540
rect 60123 12486 60169 12538
rect 60169 12486 60179 12538
rect 60203 12486 60233 12538
rect 60233 12486 60245 12538
rect 60245 12486 60259 12538
rect 60283 12486 60297 12538
rect 60297 12486 60309 12538
rect 60309 12486 60339 12538
rect 60363 12486 60373 12538
rect 60373 12486 60419 12538
rect 60123 12484 60179 12486
rect 60203 12484 60259 12486
rect 60283 12484 60339 12486
rect 60363 12484 60419 12486
rect 60646 13132 60648 13152
rect 60648 13132 60700 13152
rect 60700 13132 60702 13152
rect 60646 13096 60702 13132
rect 60830 12960 60886 13016
rect 60123 11450 60179 11452
rect 60203 11450 60259 11452
rect 60283 11450 60339 11452
rect 60363 11450 60419 11452
rect 60123 11398 60169 11450
rect 60169 11398 60179 11450
rect 60203 11398 60233 11450
rect 60233 11398 60245 11450
rect 60245 11398 60259 11450
rect 60283 11398 60297 11450
rect 60297 11398 60309 11450
rect 60309 11398 60339 11450
rect 60363 11398 60373 11450
rect 60373 11398 60419 11450
rect 60123 11396 60179 11398
rect 60203 11396 60259 11398
rect 60283 11396 60339 11398
rect 60363 11396 60419 11398
rect 60123 10362 60179 10364
rect 60203 10362 60259 10364
rect 60283 10362 60339 10364
rect 60363 10362 60419 10364
rect 60123 10310 60169 10362
rect 60169 10310 60179 10362
rect 60203 10310 60233 10362
rect 60233 10310 60245 10362
rect 60245 10310 60259 10362
rect 60283 10310 60297 10362
rect 60297 10310 60309 10362
rect 60309 10310 60339 10362
rect 60363 10310 60373 10362
rect 60373 10310 60419 10362
rect 60123 10308 60179 10310
rect 60203 10308 60259 10310
rect 60283 10308 60339 10310
rect 60363 10308 60419 10310
rect 60002 10104 60058 10160
rect 60462 9696 60518 9752
rect 60123 9274 60179 9276
rect 60203 9274 60259 9276
rect 60283 9274 60339 9276
rect 60363 9274 60419 9276
rect 60123 9222 60169 9274
rect 60169 9222 60179 9274
rect 60203 9222 60233 9274
rect 60233 9222 60245 9274
rect 60245 9222 60259 9274
rect 60283 9222 60297 9274
rect 60297 9222 60309 9274
rect 60309 9222 60339 9274
rect 60363 9222 60373 9274
rect 60373 9222 60419 9274
rect 60123 9220 60179 9222
rect 60203 9220 60259 9222
rect 60283 9220 60339 9222
rect 60363 9220 60419 9222
rect 60123 8186 60179 8188
rect 60203 8186 60259 8188
rect 60283 8186 60339 8188
rect 60363 8186 60419 8188
rect 60123 8134 60169 8186
rect 60169 8134 60179 8186
rect 60203 8134 60233 8186
rect 60233 8134 60245 8186
rect 60245 8134 60259 8186
rect 60283 8134 60297 8186
rect 60297 8134 60309 8186
rect 60309 8134 60339 8186
rect 60363 8134 60373 8186
rect 60373 8134 60419 8186
rect 60123 8132 60179 8134
rect 60203 8132 60259 8134
rect 60283 8132 60339 8134
rect 60363 8132 60419 8134
rect 60830 10104 60886 10160
rect 61566 11756 61622 11792
rect 61566 11736 61568 11756
rect 61568 11736 61620 11756
rect 61620 11736 61622 11756
rect 60123 7098 60179 7100
rect 60203 7098 60259 7100
rect 60283 7098 60339 7100
rect 60363 7098 60419 7100
rect 60123 7046 60169 7098
rect 60169 7046 60179 7098
rect 60203 7046 60233 7098
rect 60233 7046 60245 7098
rect 60245 7046 60259 7098
rect 60283 7046 60297 7098
rect 60297 7046 60309 7098
rect 60309 7046 60339 7098
rect 60363 7046 60373 7098
rect 60373 7046 60419 7098
rect 60123 7044 60179 7046
rect 60203 7044 60259 7046
rect 60283 7044 60339 7046
rect 60363 7044 60419 7046
rect 60123 6010 60179 6012
rect 60203 6010 60259 6012
rect 60283 6010 60339 6012
rect 60363 6010 60419 6012
rect 60123 5958 60169 6010
rect 60169 5958 60179 6010
rect 60203 5958 60233 6010
rect 60233 5958 60245 6010
rect 60245 5958 60259 6010
rect 60283 5958 60297 6010
rect 60297 5958 60309 6010
rect 60309 5958 60339 6010
rect 60363 5958 60373 6010
rect 60373 5958 60419 6010
rect 60123 5956 60179 5958
rect 60203 5956 60259 5958
rect 60283 5956 60339 5958
rect 60363 5956 60419 5958
rect 60123 4922 60179 4924
rect 60203 4922 60259 4924
rect 60283 4922 60339 4924
rect 60363 4922 60419 4924
rect 60123 4870 60169 4922
rect 60169 4870 60179 4922
rect 60203 4870 60233 4922
rect 60233 4870 60245 4922
rect 60245 4870 60259 4922
rect 60283 4870 60297 4922
rect 60297 4870 60309 4922
rect 60309 4870 60339 4922
rect 60363 4870 60373 4922
rect 60373 4870 60419 4922
rect 60123 4868 60179 4870
rect 60203 4868 60259 4870
rect 60283 4868 60339 4870
rect 60363 4868 60419 4870
rect 60123 3834 60179 3836
rect 60203 3834 60259 3836
rect 60283 3834 60339 3836
rect 60363 3834 60419 3836
rect 60123 3782 60169 3834
rect 60169 3782 60179 3834
rect 60203 3782 60233 3834
rect 60233 3782 60245 3834
rect 60245 3782 60259 3834
rect 60283 3782 60297 3834
rect 60297 3782 60309 3834
rect 60309 3782 60339 3834
rect 60363 3782 60373 3834
rect 60373 3782 60419 3834
rect 60123 3780 60179 3782
rect 60203 3780 60259 3782
rect 60283 3780 60339 3782
rect 60363 3780 60419 3782
rect 62578 9696 62634 9752
rect 62670 8900 62726 8936
rect 62670 8880 62672 8900
rect 62672 8880 62724 8900
rect 62724 8880 62726 8900
rect 63682 13232 63738 13288
rect 63866 10784 63922 10840
rect 63866 10668 63922 10704
rect 63866 10648 63868 10668
rect 63868 10648 63920 10668
rect 63920 10648 63922 10668
rect 60123 2746 60179 2748
rect 60203 2746 60259 2748
rect 60283 2746 60339 2748
rect 60363 2746 60419 2748
rect 60123 2694 60169 2746
rect 60169 2694 60179 2746
rect 60203 2694 60233 2746
rect 60233 2694 60245 2746
rect 60245 2694 60259 2746
rect 60283 2694 60297 2746
rect 60297 2694 60309 2746
rect 60309 2694 60339 2746
rect 60363 2694 60373 2746
rect 60373 2694 60419 2746
rect 60123 2692 60179 2694
rect 60203 2692 60259 2694
rect 60283 2692 60339 2694
rect 60363 2692 60419 2694
rect 66166 12688 66222 12744
rect 67730 10920 67786 10976
rect 67638 9968 67694 10024
rect 67638 9696 67694 9752
rect 69662 13096 69718 13152
rect 70490 10104 70546 10160
rect 70214 8336 70270 8392
rect 71226 10104 71282 10160
rect 72974 11092 72976 11112
rect 72976 11092 73028 11112
rect 73028 11092 73030 11112
rect 72974 11056 73030 11092
rect 72882 7404 72938 7440
rect 72882 7384 72884 7404
rect 72884 7384 72936 7404
rect 72936 7384 72938 7404
rect 74814 12552 74870 12608
rect 74630 10920 74686 10976
rect 74722 9988 74778 10024
rect 74722 9968 74724 9988
rect 74724 9968 74776 9988
rect 74776 9968 74778 9988
rect 77482 13504 77538 13560
rect 76838 13096 76894 13152
rect 77390 12980 77446 13016
rect 77390 12960 77392 12980
rect 77392 12960 77444 12980
rect 77444 12960 77446 12980
rect 77298 12416 77354 12472
rect 77298 12164 77354 12200
rect 77298 12144 77300 12164
rect 77300 12144 77352 12164
rect 77352 12144 77354 12164
rect 78586 12280 78642 12336
rect 79966 13232 80022 13288
rect 80242 13096 80298 13152
rect 79845 13082 79901 13084
rect 79925 13082 79981 13084
rect 80005 13082 80061 13084
rect 80085 13082 80141 13084
rect 79845 13030 79891 13082
rect 79891 13030 79901 13082
rect 79925 13030 79955 13082
rect 79955 13030 79967 13082
rect 79967 13030 79981 13082
rect 80005 13030 80019 13082
rect 80019 13030 80031 13082
rect 80031 13030 80061 13082
rect 80085 13030 80095 13082
rect 80095 13030 80141 13082
rect 79845 13028 79901 13030
rect 79925 13028 79981 13030
rect 80005 13028 80061 13030
rect 80085 13028 80141 13030
rect 79506 12980 79562 13016
rect 79506 12960 79508 12980
rect 79508 12960 79560 12980
rect 79560 12960 79562 12980
rect 80242 12416 80298 12472
rect 77850 9560 77906 9616
rect 78770 11600 78826 11656
rect 74814 3440 74870 3496
rect 76378 4548 76434 4584
rect 76378 4528 76380 4548
rect 76380 4528 76432 4548
rect 76432 4528 76434 4548
rect 79845 11994 79901 11996
rect 79925 11994 79981 11996
rect 80005 11994 80061 11996
rect 80085 11994 80141 11996
rect 79845 11942 79891 11994
rect 79891 11942 79901 11994
rect 79925 11942 79955 11994
rect 79955 11942 79967 11994
rect 79967 11942 79981 11994
rect 80005 11942 80019 11994
rect 80019 11942 80031 11994
rect 80031 11942 80061 11994
rect 80085 11942 80095 11994
rect 80095 11942 80141 11994
rect 79845 11940 79901 11942
rect 79925 11940 79981 11942
rect 80005 11940 80061 11942
rect 80085 11940 80141 11942
rect 79845 10906 79901 10908
rect 79925 10906 79981 10908
rect 80005 10906 80061 10908
rect 80085 10906 80141 10908
rect 79845 10854 79891 10906
rect 79891 10854 79901 10906
rect 79925 10854 79955 10906
rect 79955 10854 79967 10906
rect 79967 10854 79981 10906
rect 80005 10854 80019 10906
rect 80019 10854 80031 10906
rect 80031 10854 80061 10906
rect 80085 10854 80095 10906
rect 80095 10854 80141 10906
rect 79845 10852 79901 10854
rect 79925 10852 79981 10854
rect 80005 10852 80061 10854
rect 80085 10852 80141 10854
rect 79874 10684 79876 10704
rect 79876 10684 79928 10704
rect 79928 10684 79930 10704
rect 79874 10648 79930 10684
rect 79845 9818 79901 9820
rect 79925 9818 79981 9820
rect 80005 9818 80061 9820
rect 80085 9818 80141 9820
rect 79845 9766 79891 9818
rect 79891 9766 79901 9818
rect 79925 9766 79955 9818
rect 79955 9766 79967 9818
rect 79967 9766 79981 9818
rect 80005 9766 80019 9818
rect 80019 9766 80031 9818
rect 80031 9766 80061 9818
rect 80085 9766 80095 9818
rect 80095 9766 80141 9818
rect 79845 9764 79901 9766
rect 79925 9764 79981 9766
rect 80005 9764 80061 9766
rect 80085 9764 80141 9766
rect 79845 8730 79901 8732
rect 79925 8730 79981 8732
rect 80005 8730 80061 8732
rect 80085 8730 80141 8732
rect 79845 8678 79891 8730
rect 79891 8678 79901 8730
rect 79925 8678 79955 8730
rect 79955 8678 79967 8730
rect 79967 8678 79981 8730
rect 80005 8678 80019 8730
rect 80019 8678 80031 8730
rect 80031 8678 80061 8730
rect 80085 8678 80095 8730
rect 80095 8678 80141 8730
rect 79845 8676 79901 8678
rect 79925 8676 79981 8678
rect 80005 8676 80061 8678
rect 80085 8676 80141 8678
rect 79845 7642 79901 7644
rect 79925 7642 79981 7644
rect 80005 7642 80061 7644
rect 80085 7642 80141 7644
rect 79845 7590 79891 7642
rect 79891 7590 79901 7642
rect 79925 7590 79955 7642
rect 79955 7590 79967 7642
rect 79967 7590 79981 7642
rect 80005 7590 80019 7642
rect 80019 7590 80031 7642
rect 80031 7590 80061 7642
rect 80085 7590 80095 7642
rect 80095 7590 80141 7642
rect 79845 7588 79901 7590
rect 79925 7588 79981 7590
rect 80005 7588 80061 7590
rect 80085 7588 80141 7590
rect 79845 6554 79901 6556
rect 79925 6554 79981 6556
rect 80005 6554 80061 6556
rect 80085 6554 80141 6556
rect 79845 6502 79891 6554
rect 79891 6502 79901 6554
rect 79925 6502 79955 6554
rect 79955 6502 79967 6554
rect 79967 6502 79981 6554
rect 80005 6502 80019 6554
rect 80019 6502 80031 6554
rect 80031 6502 80061 6554
rect 80085 6502 80095 6554
rect 80095 6502 80141 6554
rect 79845 6500 79901 6502
rect 79925 6500 79981 6502
rect 80005 6500 80061 6502
rect 80085 6500 80141 6502
rect 79845 5466 79901 5468
rect 79925 5466 79981 5468
rect 80005 5466 80061 5468
rect 80085 5466 80141 5468
rect 79845 5414 79891 5466
rect 79891 5414 79901 5466
rect 79925 5414 79955 5466
rect 79955 5414 79967 5466
rect 79967 5414 79981 5466
rect 80005 5414 80019 5466
rect 80019 5414 80031 5466
rect 80031 5414 80061 5466
rect 80085 5414 80095 5466
rect 80095 5414 80141 5466
rect 79845 5412 79901 5414
rect 79925 5412 79981 5414
rect 80005 5412 80061 5414
rect 80085 5412 80141 5414
rect 79845 4378 79901 4380
rect 79925 4378 79981 4380
rect 80005 4378 80061 4380
rect 80085 4378 80141 4380
rect 79845 4326 79891 4378
rect 79891 4326 79901 4378
rect 79925 4326 79955 4378
rect 79955 4326 79967 4378
rect 79967 4326 79981 4378
rect 80005 4326 80019 4378
rect 80019 4326 80031 4378
rect 80031 4326 80061 4378
rect 80085 4326 80095 4378
rect 80095 4326 80141 4378
rect 79845 4324 79901 4326
rect 79925 4324 79981 4326
rect 80005 4324 80061 4326
rect 80085 4324 80141 4326
rect 81530 13232 81586 13288
rect 81346 12416 81402 12472
rect 82174 13504 82230 13560
rect 81898 12280 81954 12336
rect 82082 12280 82138 12336
rect 81254 10956 81256 10976
rect 81256 10956 81308 10976
rect 81308 10956 81310 10976
rect 81254 10920 81310 10956
rect 81254 9832 81310 9888
rect 79845 3290 79901 3292
rect 79925 3290 79981 3292
rect 80005 3290 80061 3292
rect 80085 3290 80141 3292
rect 79845 3238 79891 3290
rect 79891 3238 79901 3290
rect 79925 3238 79955 3290
rect 79955 3238 79967 3290
rect 79967 3238 79981 3290
rect 80005 3238 80019 3290
rect 80019 3238 80031 3290
rect 80031 3238 80061 3290
rect 80085 3238 80095 3290
rect 80095 3238 80141 3290
rect 79845 3236 79901 3238
rect 79925 3236 79981 3238
rect 80005 3236 80061 3238
rect 80085 3236 80141 3238
rect 83186 12416 83242 12472
rect 83370 8472 83426 8528
rect 85486 12280 85542 12336
rect 86682 11600 86738 11656
rect 86222 11328 86278 11384
rect 84842 9832 84898 9888
rect 86866 10920 86922 10976
rect 87234 10532 87290 10568
rect 87234 10512 87236 10532
rect 87236 10512 87288 10532
rect 87288 10512 87290 10532
rect 88154 11464 88210 11520
rect 87786 9288 87842 9344
rect 88890 13132 88892 13152
rect 88892 13132 88944 13152
rect 88944 13132 88946 13152
rect 88890 13096 88946 13132
rect 88982 12552 89038 12608
rect 88246 9696 88302 9752
rect 88338 8780 88340 8800
rect 88340 8780 88392 8800
rect 88392 8780 88394 8800
rect 88338 8744 88394 8780
rect 89258 13252 89314 13288
rect 89258 13232 89260 13252
rect 89260 13232 89312 13252
rect 89312 13232 89314 13252
rect 90362 11464 90418 11520
rect 89350 7520 89406 7576
rect 90086 9696 90142 9752
rect 89718 9016 89774 9072
rect 90454 9324 90456 9344
rect 90456 9324 90508 9344
rect 90508 9324 90510 9344
rect 90454 9288 90510 9324
rect 89810 7520 89866 7576
rect 90914 9016 90970 9072
rect 91098 8608 91154 8664
rect 90730 7812 90786 7848
rect 90730 7792 90732 7812
rect 90732 7792 90784 7812
rect 90784 7792 90786 7812
rect 90822 7692 90824 7712
rect 90824 7692 90876 7712
rect 90876 7692 90878 7712
rect 90822 7656 90878 7692
rect 90822 7520 90878 7576
rect 91374 7248 91430 7304
rect 91466 6316 91522 6352
rect 91466 6296 91468 6316
rect 91468 6296 91520 6316
rect 91520 6296 91522 6316
rect 93398 12688 93454 12744
rect 92846 11192 92902 11248
rect 92754 9424 92810 9480
rect 92478 8744 92534 8800
rect 93214 10240 93270 10296
rect 93214 8744 93270 8800
rect 94410 13096 94466 13152
rect 93674 11328 93730 11384
rect 93490 7540 93546 7576
rect 93490 7520 93492 7540
rect 93492 7520 93544 7540
rect 93544 7520 93546 7540
rect 95882 13368 95938 13424
rect 93858 9016 93914 9072
rect 93766 7792 93822 7848
rect 93950 7520 94006 7576
rect 93858 7248 93914 7304
rect 96986 13268 96988 13288
rect 96988 13268 97040 13288
rect 97040 13268 97042 13288
rect 96986 13232 97042 13268
rect 95330 9832 95386 9888
rect 95514 10240 95570 10296
rect 95330 8880 95386 8936
rect 95146 7692 95148 7712
rect 95148 7692 95200 7712
rect 95200 7692 95202 7712
rect 95146 7656 95202 7692
rect 93490 3032 93546 3088
rect 97722 13096 97778 13152
rect 96802 12280 96858 12336
rect 96802 11736 96858 11792
rect 98458 11736 98514 11792
rect 99568 13626 99624 13628
rect 99648 13626 99704 13628
rect 99728 13626 99784 13628
rect 99808 13626 99864 13628
rect 99568 13574 99614 13626
rect 99614 13574 99624 13626
rect 99648 13574 99678 13626
rect 99678 13574 99690 13626
rect 99690 13574 99704 13626
rect 99728 13574 99742 13626
rect 99742 13574 99754 13626
rect 99754 13574 99784 13626
rect 99808 13574 99818 13626
rect 99818 13574 99864 13626
rect 99568 13572 99624 13574
rect 99648 13572 99704 13574
rect 99728 13572 99784 13574
rect 99808 13572 99864 13574
rect 96710 2896 96766 2952
rect 99378 11636 99380 11656
rect 99380 11636 99432 11656
rect 99432 11636 99434 11656
rect 99378 11600 99434 11636
rect 99930 13232 99986 13288
rect 99568 12538 99624 12540
rect 99648 12538 99704 12540
rect 99728 12538 99784 12540
rect 99808 12538 99864 12540
rect 99568 12486 99614 12538
rect 99614 12486 99624 12538
rect 99648 12486 99678 12538
rect 99678 12486 99690 12538
rect 99690 12486 99704 12538
rect 99728 12486 99742 12538
rect 99742 12486 99754 12538
rect 99754 12486 99784 12538
rect 99808 12486 99818 12538
rect 99818 12486 99864 12538
rect 99568 12484 99624 12486
rect 99648 12484 99704 12486
rect 99728 12484 99784 12486
rect 99808 12484 99864 12486
rect 100298 13096 100354 13152
rect 99568 11450 99624 11452
rect 99648 11450 99704 11452
rect 99728 11450 99784 11452
rect 99808 11450 99864 11452
rect 99568 11398 99614 11450
rect 99614 11398 99624 11450
rect 99648 11398 99678 11450
rect 99678 11398 99690 11450
rect 99690 11398 99704 11450
rect 99728 11398 99742 11450
rect 99742 11398 99754 11450
rect 99754 11398 99784 11450
rect 99808 11398 99818 11450
rect 99818 11398 99864 11450
rect 99568 11396 99624 11398
rect 99648 11396 99704 11398
rect 99728 11396 99784 11398
rect 99808 11396 99864 11398
rect 99568 10362 99624 10364
rect 99648 10362 99704 10364
rect 99728 10362 99784 10364
rect 99808 10362 99864 10364
rect 99568 10310 99614 10362
rect 99614 10310 99624 10362
rect 99648 10310 99678 10362
rect 99678 10310 99690 10362
rect 99690 10310 99704 10362
rect 99728 10310 99742 10362
rect 99742 10310 99754 10362
rect 99754 10310 99784 10362
rect 99808 10310 99818 10362
rect 99818 10310 99864 10362
rect 99568 10308 99624 10310
rect 99648 10308 99704 10310
rect 99728 10308 99784 10310
rect 99808 10308 99864 10310
rect 99568 9274 99624 9276
rect 99648 9274 99704 9276
rect 99728 9274 99784 9276
rect 99808 9274 99864 9276
rect 99568 9222 99614 9274
rect 99614 9222 99624 9274
rect 99648 9222 99678 9274
rect 99678 9222 99690 9274
rect 99690 9222 99704 9274
rect 99728 9222 99742 9274
rect 99742 9222 99754 9274
rect 99754 9222 99784 9274
rect 99808 9222 99818 9274
rect 99818 9222 99864 9274
rect 99568 9220 99624 9222
rect 99648 9220 99704 9222
rect 99728 9220 99784 9222
rect 99808 9220 99864 9222
rect 99568 8186 99624 8188
rect 99648 8186 99704 8188
rect 99728 8186 99784 8188
rect 99808 8186 99864 8188
rect 99568 8134 99614 8186
rect 99614 8134 99624 8186
rect 99648 8134 99678 8186
rect 99678 8134 99690 8186
rect 99690 8134 99704 8186
rect 99728 8134 99742 8186
rect 99742 8134 99754 8186
rect 99754 8134 99784 8186
rect 99808 8134 99818 8186
rect 99818 8134 99864 8186
rect 99568 8132 99624 8134
rect 99648 8132 99704 8134
rect 99728 8132 99784 8134
rect 99808 8132 99864 8134
rect 99568 7098 99624 7100
rect 99648 7098 99704 7100
rect 99728 7098 99784 7100
rect 99808 7098 99864 7100
rect 99568 7046 99614 7098
rect 99614 7046 99624 7098
rect 99648 7046 99678 7098
rect 99678 7046 99690 7098
rect 99690 7046 99704 7098
rect 99728 7046 99742 7098
rect 99742 7046 99754 7098
rect 99754 7046 99784 7098
rect 99808 7046 99818 7098
rect 99818 7046 99864 7098
rect 99568 7044 99624 7046
rect 99648 7044 99704 7046
rect 99728 7044 99784 7046
rect 99808 7044 99864 7046
rect 99568 6010 99624 6012
rect 99648 6010 99704 6012
rect 99728 6010 99784 6012
rect 99808 6010 99864 6012
rect 99568 5958 99614 6010
rect 99614 5958 99624 6010
rect 99648 5958 99678 6010
rect 99678 5958 99690 6010
rect 99690 5958 99704 6010
rect 99728 5958 99742 6010
rect 99742 5958 99754 6010
rect 99754 5958 99784 6010
rect 99808 5958 99818 6010
rect 99818 5958 99864 6010
rect 99568 5956 99624 5958
rect 99648 5956 99704 5958
rect 99728 5956 99784 5958
rect 99808 5956 99864 5958
rect 99930 5208 99986 5264
rect 100666 11056 100722 11112
rect 100666 8880 100722 8936
rect 100390 7656 100446 7712
rect 100758 6840 100814 6896
rect 100298 6160 100354 6216
rect 100022 5072 100078 5128
rect 99568 4922 99624 4924
rect 99648 4922 99704 4924
rect 99728 4922 99784 4924
rect 99808 4922 99864 4924
rect 99568 4870 99614 4922
rect 99614 4870 99624 4922
rect 99648 4870 99678 4922
rect 99678 4870 99690 4922
rect 99690 4870 99704 4922
rect 99728 4870 99742 4922
rect 99742 4870 99754 4922
rect 99754 4870 99784 4922
rect 99808 4870 99818 4922
rect 99818 4870 99864 4922
rect 99568 4868 99624 4870
rect 99648 4868 99704 4870
rect 99728 4868 99784 4870
rect 99808 4868 99864 4870
rect 99568 3834 99624 3836
rect 99648 3834 99704 3836
rect 99728 3834 99784 3836
rect 99808 3834 99864 3836
rect 99568 3782 99614 3834
rect 99614 3782 99624 3834
rect 99648 3782 99678 3834
rect 99678 3782 99690 3834
rect 99690 3782 99704 3834
rect 99728 3782 99742 3834
rect 99742 3782 99754 3834
rect 99754 3782 99784 3834
rect 99808 3782 99818 3834
rect 99818 3782 99864 3834
rect 99568 3780 99624 3782
rect 99648 3780 99704 3782
rect 99728 3780 99784 3782
rect 99808 3780 99864 3782
rect 101862 10240 101918 10296
rect 101862 6024 101918 6080
rect 99568 2746 99624 2748
rect 99648 2746 99704 2748
rect 99728 2746 99784 2748
rect 99808 2746 99864 2748
rect 99568 2694 99614 2746
rect 99614 2694 99624 2746
rect 99648 2694 99678 2746
rect 99678 2694 99690 2746
rect 99690 2694 99704 2746
rect 99728 2694 99742 2746
rect 99742 2694 99754 2746
rect 99754 2694 99784 2746
rect 99808 2694 99818 2746
rect 99818 2694 99864 2746
rect 99568 2692 99624 2694
rect 99648 2692 99704 2694
rect 99728 2692 99784 2694
rect 99808 2692 99864 2694
rect 95606 2352 95662 2408
rect 40400 2202 40456 2204
rect 40480 2202 40536 2204
rect 40560 2202 40616 2204
rect 40640 2202 40696 2204
rect 40400 2150 40446 2202
rect 40446 2150 40456 2202
rect 40480 2150 40510 2202
rect 40510 2150 40522 2202
rect 40522 2150 40536 2202
rect 40560 2150 40574 2202
rect 40574 2150 40586 2202
rect 40586 2150 40616 2202
rect 40640 2150 40650 2202
rect 40650 2150 40696 2202
rect 40400 2148 40456 2150
rect 40480 2148 40536 2150
rect 40560 2148 40616 2150
rect 40640 2148 40696 2150
rect 79845 2202 79901 2204
rect 79925 2202 79981 2204
rect 80005 2202 80061 2204
rect 80085 2202 80141 2204
rect 79845 2150 79891 2202
rect 79891 2150 79901 2202
rect 79925 2150 79955 2202
rect 79955 2150 79967 2202
rect 79967 2150 79981 2202
rect 80005 2150 80019 2202
rect 80019 2150 80031 2202
rect 80031 2150 80061 2202
rect 80085 2150 80095 2202
rect 80095 2150 80141 2202
rect 79845 2148 79901 2150
rect 79925 2148 79981 2150
rect 80005 2148 80061 2150
rect 80085 2148 80141 2150
rect 1674 1944 1730 2000
rect 103886 12724 103888 12744
rect 103888 12724 103940 12744
rect 103940 12724 103942 12744
rect 103886 12688 103942 12724
rect 102506 6840 102562 6896
rect 104346 12008 104402 12064
rect 104162 10376 104218 10432
rect 104162 9832 104218 9888
rect 104714 10104 104770 10160
rect 104990 10240 105046 10296
rect 105174 10240 105230 10296
rect 104714 7928 104770 7984
rect 105818 12044 105820 12064
rect 105820 12044 105872 12064
rect 105872 12044 105874 12064
rect 105818 12008 105874 12044
rect 106462 6704 106518 6760
rect 107842 10784 107898 10840
rect 107750 10648 107806 10704
rect 107750 10104 107806 10160
rect 107842 9696 107898 9752
rect 107658 8608 107714 8664
rect 107842 8608 107898 8664
rect 107106 6432 107162 6488
rect 106922 5888 106978 5944
rect 106002 3884 106004 3904
rect 106004 3884 106056 3904
rect 106056 3884 106058 3904
rect 106002 3848 106058 3884
rect 107934 8064 107990 8120
rect 107382 5636 107438 5672
rect 107382 5616 107384 5636
rect 107384 5616 107436 5636
rect 107436 5616 107438 5636
rect 109038 10804 109094 10840
rect 109038 10784 109040 10804
rect 109040 10784 109092 10804
rect 109092 10784 109094 10804
rect 108854 7792 108910 7848
rect 109222 4392 109278 4448
rect 110418 13132 110420 13152
rect 110420 13132 110472 13152
rect 110472 13132 110474 13152
rect 110418 13096 110474 13132
rect 110418 12416 110474 12472
rect 110050 8200 110106 8256
rect 110326 7268 110382 7304
rect 110326 7248 110328 7268
rect 110328 7248 110380 7268
rect 110380 7248 110382 7268
rect 110602 6976 110658 7032
rect 110602 6568 110658 6624
rect 108302 1944 108358 2000
rect 111614 10104 111670 10160
rect 112626 9560 112682 9616
rect 112534 8064 112590 8120
rect 111982 5888 112038 5944
rect 113086 13096 113142 13152
rect 113086 9868 113088 9888
rect 113088 9868 113140 9888
rect 113140 9868 113142 9888
rect 113086 9832 113142 9868
rect 113454 10648 113510 10704
rect 113546 10104 113602 10160
rect 113362 8064 113418 8120
rect 112442 7284 112444 7304
rect 112444 7284 112496 7304
rect 112496 7284 112498 7304
rect 112442 7248 112498 7284
rect 112626 7248 112682 7304
rect 113270 7792 113326 7848
rect 112718 4120 112774 4176
rect 113730 5652 113732 5672
rect 113732 5652 113784 5672
rect 113784 5652 113786 5672
rect 113730 5616 113786 5652
rect 114006 6704 114062 6760
rect 114466 8744 114522 8800
rect 114466 6976 114522 7032
rect 115662 12824 115718 12880
rect 114926 9560 114982 9616
rect 114742 7656 114798 7712
rect 114742 6704 114798 6760
rect 114282 1672 114338 1728
rect 116122 12588 116124 12608
rect 116124 12588 116176 12608
rect 116176 12588 116178 12608
rect 116122 12552 116178 12588
rect 116950 13640 117006 13696
rect 116490 12008 116546 12064
rect 115294 9152 115350 9208
rect 115294 8336 115350 8392
rect 115570 9288 115626 9344
rect 115570 8608 115626 8664
rect 115478 6568 115534 6624
rect 115386 6432 115442 6488
rect 115386 6296 115442 6352
rect 115386 5616 115442 5672
rect 115386 4392 115442 4448
rect 115294 3984 115350 4040
rect 116030 10784 116086 10840
rect 115846 9696 115902 9752
rect 115938 8472 115994 8528
rect 116950 11056 117006 11112
rect 117318 11736 117374 11792
rect 116950 9696 117006 9752
rect 116858 8744 116914 8800
rect 116214 7812 116270 7848
rect 116214 7792 116216 7812
rect 116216 7792 116268 7812
rect 116268 7792 116270 7812
rect 116766 8336 116822 8392
rect 117226 8744 117282 8800
rect 117410 6976 117466 7032
rect 116950 5752 117006 5808
rect 117410 5908 117466 5944
rect 117410 5888 117412 5908
rect 117412 5888 117464 5908
rect 117464 5888 117466 5908
rect 117226 4820 117282 4856
rect 117226 4800 117228 4820
rect 117228 4800 117280 4820
rect 117280 4800 117282 4820
rect 117778 4664 117834 4720
rect 118514 10648 118570 10704
rect 119290 13082 119346 13084
rect 119370 13082 119426 13084
rect 119450 13082 119506 13084
rect 119530 13082 119586 13084
rect 119290 13030 119336 13082
rect 119336 13030 119346 13082
rect 119370 13030 119400 13082
rect 119400 13030 119412 13082
rect 119412 13030 119426 13082
rect 119450 13030 119464 13082
rect 119464 13030 119476 13082
rect 119476 13030 119506 13082
rect 119530 13030 119540 13082
rect 119540 13030 119586 13082
rect 119290 13028 119346 13030
rect 119370 13028 119426 13030
rect 119450 13028 119506 13030
rect 119530 13028 119586 13030
rect 119066 12008 119122 12064
rect 118882 11872 118938 11928
rect 120906 12960 120962 13016
rect 121366 14048 121422 14104
rect 121458 13232 121514 13288
rect 119290 11994 119346 11996
rect 119370 11994 119426 11996
rect 119450 11994 119506 11996
rect 119530 11994 119586 11996
rect 119290 11942 119336 11994
rect 119336 11942 119346 11994
rect 119370 11942 119400 11994
rect 119400 11942 119412 11994
rect 119412 11942 119426 11994
rect 119450 11942 119464 11994
rect 119464 11942 119476 11994
rect 119476 11942 119506 11994
rect 119530 11942 119540 11994
rect 119540 11942 119586 11994
rect 119290 11940 119346 11942
rect 119370 11940 119426 11942
rect 119450 11940 119506 11942
rect 119530 11940 119586 11942
rect 118238 9968 118294 10024
rect 118422 8336 118478 8392
rect 118974 10784 119030 10840
rect 119290 10906 119346 10908
rect 119370 10906 119426 10908
rect 119450 10906 119506 10908
rect 119530 10906 119586 10908
rect 119290 10854 119336 10906
rect 119336 10854 119346 10906
rect 119370 10854 119400 10906
rect 119400 10854 119412 10906
rect 119412 10854 119426 10906
rect 119450 10854 119464 10906
rect 119464 10854 119476 10906
rect 119476 10854 119506 10906
rect 119530 10854 119540 10906
rect 119540 10854 119586 10906
rect 119290 10852 119346 10854
rect 119370 10852 119426 10854
rect 119450 10852 119506 10854
rect 119530 10852 119586 10854
rect 118974 8492 119030 8528
rect 118974 8472 118976 8492
rect 118976 8472 119028 8492
rect 119028 8472 119030 8492
rect 119290 9818 119346 9820
rect 119370 9818 119426 9820
rect 119450 9818 119506 9820
rect 119530 9818 119586 9820
rect 119290 9766 119336 9818
rect 119336 9766 119346 9818
rect 119370 9766 119400 9818
rect 119400 9766 119412 9818
rect 119412 9766 119426 9818
rect 119450 9766 119464 9818
rect 119464 9766 119476 9818
rect 119476 9766 119506 9818
rect 119530 9766 119540 9818
rect 119540 9766 119586 9818
rect 119290 9764 119346 9766
rect 119370 9764 119426 9766
rect 119450 9764 119506 9766
rect 119530 9764 119586 9766
rect 119158 9696 119214 9752
rect 119158 8780 119160 8800
rect 119160 8780 119212 8800
rect 119212 8780 119214 8800
rect 119158 8744 119214 8780
rect 119290 8730 119346 8732
rect 119370 8730 119426 8732
rect 119450 8730 119506 8732
rect 119530 8730 119586 8732
rect 119290 8678 119336 8730
rect 119336 8678 119346 8730
rect 119370 8678 119400 8730
rect 119400 8678 119412 8730
rect 119412 8678 119426 8730
rect 119450 8678 119464 8730
rect 119464 8678 119476 8730
rect 119476 8678 119506 8730
rect 119530 8678 119540 8730
rect 119540 8678 119586 8730
rect 119290 8676 119346 8678
rect 119370 8676 119426 8678
rect 119450 8676 119506 8678
rect 119530 8676 119586 8678
rect 118698 4800 118754 4856
rect 118238 3712 118294 3768
rect 119290 7642 119346 7644
rect 119370 7642 119426 7644
rect 119450 7642 119506 7644
rect 119530 7642 119586 7644
rect 119290 7590 119336 7642
rect 119336 7590 119346 7642
rect 119370 7590 119400 7642
rect 119400 7590 119412 7642
rect 119412 7590 119426 7642
rect 119450 7590 119464 7642
rect 119464 7590 119476 7642
rect 119476 7590 119506 7642
rect 119530 7590 119540 7642
rect 119540 7590 119586 7642
rect 119290 7588 119346 7590
rect 119370 7588 119426 7590
rect 119450 7588 119506 7590
rect 119530 7588 119586 7590
rect 119290 6554 119346 6556
rect 119370 6554 119426 6556
rect 119450 6554 119506 6556
rect 119530 6554 119586 6556
rect 119290 6502 119336 6554
rect 119336 6502 119346 6554
rect 119370 6502 119400 6554
rect 119400 6502 119412 6554
rect 119412 6502 119426 6554
rect 119450 6502 119464 6554
rect 119464 6502 119476 6554
rect 119476 6502 119506 6554
rect 119530 6502 119540 6554
rect 119540 6502 119586 6554
rect 119290 6500 119346 6502
rect 119370 6500 119426 6502
rect 119450 6500 119506 6502
rect 119530 6500 119586 6502
rect 119290 5466 119346 5468
rect 119370 5466 119426 5468
rect 119450 5466 119506 5468
rect 119530 5466 119586 5468
rect 119290 5414 119336 5466
rect 119336 5414 119346 5466
rect 119370 5414 119400 5466
rect 119400 5414 119412 5466
rect 119412 5414 119426 5466
rect 119450 5414 119464 5466
rect 119464 5414 119476 5466
rect 119476 5414 119506 5466
rect 119530 5414 119540 5466
rect 119540 5414 119586 5466
rect 119290 5412 119346 5414
rect 119370 5412 119426 5414
rect 119450 5412 119506 5414
rect 119530 5412 119586 5414
rect 119290 4378 119346 4380
rect 119370 4378 119426 4380
rect 119450 4378 119506 4380
rect 119530 4378 119586 4380
rect 119290 4326 119336 4378
rect 119336 4326 119346 4378
rect 119370 4326 119400 4378
rect 119400 4326 119412 4378
rect 119412 4326 119426 4378
rect 119450 4326 119464 4378
rect 119464 4326 119476 4378
rect 119476 4326 119506 4378
rect 119530 4326 119540 4378
rect 119540 4326 119586 4378
rect 119290 4324 119346 4326
rect 119370 4324 119426 4326
rect 119450 4324 119506 4326
rect 119530 4324 119586 4326
rect 119250 3712 119306 3768
rect 118790 3576 118846 3632
rect 117594 2796 117596 2816
rect 117596 2796 117648 2816
rect 117648 2796 117650 2816
rect 117594 2760 117650 2796
rect 118514 2624 118570 2680
rect 119290 3290 119346 3292
rect 119370 3290 119426 3292
rect 119450 3290 119506 3292
rect 119530 3290 119586 3292
rect 119290 3238 119336 3290
rect 119336 3238 119346 3290
rect 119370 3238 119400 3290
rect 119400 3238 119412 3290
rect 119412 3238 119426 3290
rect 119450 3238 119464 3290
rect 119464 3238 119476 3290
rect 119476 3238 119506 3290
rect 119530 3238 119540 3290
rect 119540 3238 119586 3290
rect 119290 3236 119346 3238
rect 119370 3236 119426 3238
rect 119450 3236 119506 3238
rect 119530 3236 119586 3238
rect 117410 2352 117466 2408
rect 119290 2202 119346 2204
rect 119370 2202 119426 2204
rect 119450 2202 119506 2204
rect 119530 2202 119586 2204
rect 119290 2150 119336 2202
rect 119336 2150 119346 2202
rect 119370 2150 119400 2202
rect 119400 2150 119412 2202
rect 119412 2150 119426 2202
rect 119450 2150 119464 2202
rect 119464 2150 119476 2202
rect 119476 2150 119506 2202
rect 119530 2150 119540 2202
rect 119540 2150 119586 2202
rect 119290 2148 119346 2150
rect 119370 2148 119426 2150
rect 119450 2148 119506 2150
rect 119530 2148 119586 2150
rect 120262 12416 120318 12472
rect 120814 12824 120870 12880
rect 122378 13096 122434 13152
rect 120170 11872 120226 11928
rect 120814 12044 120816 12064
rect 120816 12044 120868 12064
rect 120868 12044 120870 12064
rect 120814 12008 120870 12044
rect 121642 11736 121698 11792
rect 121366 11328 121422 11384
rect 121182 11192 121238 11248
rect 120354 10412 120356 10432
rect 120356 10412 120408 10432
rect 120408 10412 120410 10432
rect 120354 10376 120410 10412
rect 120722 9968 120778 10024
rect 120170 8472 120226 8528
rect 120078 6432 120134 6488
rect 120170 2760 120226 2816
rect 120722 8608 120778 8664
rect 120354 4428 120356 4448
rect 120356 4428 120408 4448
rect 120408 4428 120410 4448
rect 120354 4392 120410 4428
rect 121366 8064 121422 8120
rect 122838 12144 122894 12200
rect 121734 10376 121790 10432
rect 123298 12416 123354 12472
rect 123206 10648 123262 10704
rect 121826 9016 121882 9072
rect 122378 8780 122380 8800
rect 122380 8780 122432 8800
rect 122432 8780 122434 8800
rect 122378 8744 122434 8780
rect 121826 7112 121882 7168
rect 122930 9968 122986 10024
rect 124770 13232 124826 13288
rect 124402 13132 124404 13152
rect 124404 13132 124456 13152
rect 124456 13132 124458 13152
rect 124402 13096 124458 13132
rect 124862 12824 124918 12880
rect 123850 12180 123852 12200
rect 123852 12180 123904 12200
rect 123904 12180 123906 12200
rect 123850 12144 123906 12180
rect 123666 11192 123722 11248
rect 124310 11736 124366 11792
rect 123942 11464 123998 11520
rect 122930 8472 122986 8528
rect 122838 6976 122894 7032
rect 122746 6024 122802 6080
rect 122746 4684 122802 4720
rect 122746 4664 122748 4684
rect 122748 4664 122800 4684
rect 122800 4664 122802 4684
rect 123114 5480 123170 5536
rect 119986 2488 120042 2544
rect 123022 2624 123078 2680
rect 123574 8608 123630 8664
rect 123758 8744 123814 8800
rect 124218 11328 124274 11384
rect 124310 11192 124366 11248
rect 125690 14456 125746 14512
rect 125322 13268 125324 13288
rect 125324 13268 125376 13288
rect 125376 13268 125378 13288
rect 125322 13232 125378 13268
rect 125322 12144 125378 12200
rect 124770 10920 124826 10976
rect 124402 9696 124458 9752
rect 124402 9424 124458 9480
rect 124402 8472 124458 8528
rect 124954 11736 125010 11792
rect 124954 11328 125010 11384
rect 125506 11872 125562 11928
rect 124862 7656 124918 7712
rect 123390 3032 123446 3088
rect 124126 7112 124182 7168
rect 124402 6180 124458 6216
rect 124402 6160 124404 6180
rect 124404 6160 124456 6180
rect 124456 6160 124458 6180
rect 124586 5752 124642 5808
rect 125690 10804 125746 10840
rect 125690 10784 125692 10804
rect 125692 10784 125744 10804
rect 125744 10784 125746 10804
rect 125598 9968 125654 10024
rect 125506 7112 125562 7168
rect 125690 5752 125746 5808
rect 126334 12960 126390 13016
rect 125966 6432 126022 6488
rect 126150 10784 126206 10840
rect 126150 9968 126206 10024
rect 126150 9696 126206 9752
rect 126334 9968 126390 10024
rect 126426 8472 126482 8528
rect 127346 12960 127402 13016
rect 126610 7284 126612 7304
rect 126612 7284 126664 7304
rect 126664 7284 126666 7304
rect 126610 7248 126666 7284
rect 125874 5480 125930 5536
rect 125230 3984 125286 4040
rect 126518 6296 126574 6352
rect 127162 12280 127218 12336
rect 128450 14320 128506 14376
rect 128634 12824 128690 12880
rect 127346 11872 127402 11928
rect 126610 4256 126666 4312
rect 127070 10532 127126 10568
rect 127070 10512 127072 10532
rect 127072 10512 127124 10532
rect 127124 10512 127126 10532
rect 127070 6568 127126 6624
rect 126978 5344 127034 5400
rect 127162 5228 127218 5264
rect 127162 5208 127164 5228
rect 127164 5208 127216 5228
rect 127216 5208 127218 5228
rect 127714 12144 127770 12200
rect 127898 11192 127954 11248
rect 128082 11092 128084 11112
rect 128084 11092 128136 11112
rect 128136 11092 128138 11112
rect 128082 11056 128138 11092
rect 127990 10512 128046 10568
rect 128266 9016 128322 9072
rect 128634 10920 128690 10976
rect 129554 13232 129610 13288
rect 130382 13232 130438 13288
rect 130198 12280 130254 12336
rect 131302 12960 131358 13016
rect 130014 12008 130070 12064
rect 129094 9288 129150 9344
rect 128818 9016 128874 9072
rect 128082 8608 128138 8664
rect 128174 5888 128230 5944
rect 127990 4256 128046 4312
rect 128358 3712 128414 3768
rect 123206 1264 123262 1320
rect 128542 7248 128598 7304
rect 128634 3984 128690 4040
rect 128910 8064 128966 8120
rect 128910 7656 128966 7712
rect 129186 7656 129242 7712
rect 129094 6296 129150 6352
rect 129646 10240 129702 10296
rect 129646 7520 129702 7576
rect 128910 4664 128966 4720
rect 129922 7928 129978 7984
rect 129738 6024 129794 6080
rect 129922 6024 129978 6080
rect 129738 5480 129794 5536
rect 130290 7248 130346 7304
rect 130198 4528 130254 4584
rect 130658 12144 130714 12200
rect 130658 11056 130714 11112
rect 131210 11872 131266 11928
rect 130842 9152 130898 9208
rect 131118 9052 131120 9072
rect 131120 9052 131172 9072
rect 131172 9052 131174 9072
rect 131118 9016 131174 9052
rect 131762 10240 131818 10296
rect 131026 7792 131082 7848
rect 130842 7248 130898 7304
rect 131762 7112 131818 7168
rect 131302 5888 131358 5944
rect 130842 4256 130898 4312
rect 130750 3440 130806 3496
rect 130198 2916 130254 2952
rect 130198 2896 130200 2916
rect 130200 2896 130252 2916
rect 130252 2896 130254 2916
rect 129554 2508 129610 2544
rect 129554 2488 129556 2508
rect 129556 2488 129608 2508
rect 129608 2488 129610 2508
rect 131118 4120 131174 4176
rect 131118 3440 131174 3496
rect 132130 8900 132186 8936
rect 132130 8880 132132 8900
rect 132132 8880 132184 8900
rect 132184 8880 132186 8900
rect 132038 4120 132094 4176
rect 133142 13232 133198 13288
rect 133142 12688 133198 12744
rect 133050 11500 133052 11520
rect 133052 11500 133104 11520
rect 133104 11500 133106 11520
rect 133050 11464 133106 11500
rect 133970 12144 134026 12200
rect 134338 12688 134394 12744
rect 134522 10376 134578 10432
rect 133878 9696 133934 9752
rect 133418 6840 133474 6896
rect 133142 4120 133198 4176
rect 132774 3712 132830 3768
rect 132958 3576 133014 3632
rect 133878 7520 133934 7576
rect 133602 4120 133658 4176
rect 133878 6160 133934 6216
rect 133970 4256 134026 4312
rect 133694 3848 133750 3904
rect 131302 2488 131358 2544
rect 134430 6160 134486 6216
rect 134522 5652 134524 5672
rect 134524 5652 134576 5672
rect 134576 5652 134578 5672
rect 134522 5616 134578 5652
rect 134890 12824 134946 12880
rect 135166 10920 135222 10976
rect 134154 3168 134210 3224
rect 135166 9424 135222 9480
rect 135718 12724 135720 12744
rect 135720 12724 135772 12744
rect 135772 12724 135774 12744
rect 135718 12688 135774 12724
rect 135534 10512 135590 10568
rect 135350 6296 135406 6352
rect 135074 2624 135130 2680
rect 135626 9696 135682 9752
rect 136914 14048 136970 14104
rect 136730 12552 136786 12608
rect 136638 12416 136694 12472
rect 136914 12280 136970 12336
rect 135994 8064 136050 8120
rect 135994 2896 136050 2952
rect 136638 10512 136694 10568
rect 136362 8608 136418 8664
rect 136362 7812 136418 7848
rect 136362 7792 136364 7812
rect 136364 7792 136416 7812
rect 136416 7792 136418 7812
rect 137190 10240 137246 10296
rect 136638 7384 136694 7440
rect 138018 10784 138074 10840
rect 138018 9424 138074 9480
rect 137466 9288 137522 9344
rect 137926 9152 137982 9208
rect 137374 8900 137430 8936
rect 137374 8880 137376 8900
rect 137376 8880 137428 8900
rect 137428 8880 137430 8900
rect 137098 7384 137154 7440
rect 137098 7112 137154 7168
rect 137282 6976 137338 7032
rect 137742 5752 137798 5808
rect 137926 6840 137982 6896
rect 137834 4528 137890 4584
rect 137926 4256 137982 4312
rect 137926 3612 137928 3632
rect 137928 3612 137980 3632
rect 137980 3612 137982 3632
rect 137926 3576 137982 3612
rect 137742 3032 137798 3088
rect 134062 2216 134118 2272
rect 136638 2624 136694 2680
rect 138018 2372 138074 2408
rect 138018 2352 138020 2372
rect 138020 2352 138072 2372
rect 138072 2352 138074 2372
rect 138202 9172 138258 9208
rect 138202 9152 138204 9172
rect 138204 9152 138256 9172
rect 138256 9152 138258 9172
rect 138662 13640 138718 13696
rect 139013 13626 139069 13628
rect 139093 13626 139149 13628
rect 139173 13626 139229 13628
rect 139253 13626 139309 13628
rect 139013 13574 139059 13626
rect 139059 13574 139069 13626
rect 139093 13574 139123 13626
rect 139123 13574 139135 13626
rect 139135 13574 139149 13626
rect 139173 13574 139187 13626
rect 139187 13574 139199 13626
rect 139199 13574 139229 13626
rect 139253 13574 139263 13626
rect 139263 13574 139309 13626
rect 139013 13572 139069 13574
rect 139093 13572 139149 13574
rect 139173 13572 139229 13574
rect 139253 13572 139309 13574
rect 139013 12538 139069 12540
rect 139093 12538 139149 12540
rect 139173 12538 139229 12540
rect 139253 12538 139309 12540
rect 139013 12486 139059 12538
rect 139059 12486 139069 12538
rect 139093 12486 139123 12538
rect 139123 12486 139135 12538
rect 139135 12486 139149 12538
rect 139173 12486 139187 12538
rect 139187 12486 139199 12538
rect 139199 12486 139229 12538
rect 139253 12486 139263 12538
rect 139263 12486 139309 12538
rect 139013 12484 139069 12486
rect 139093 12484 139149 12486
rect 139173 12484 139229 12486
rect 139253 12484 139309 12486
rect 139013 11450 139069 11452
rect 139093 11450 139149 11452
rect 139173 11450 139229 11452
rect 139253 11450 139309 11452
rect 139013 11398 139059 11450
rect 139059 11398 139069 11450
rect 139093 11398 139123 11450
rect 139123 11398 139135 11450
rect 139135 11398 139149 11450
rect 139173 11398 139187 11450
rect 139187 11398 139199 11450
rect 139199 11398 139229 11450
rect 139253 11398 139263 11450
rect 139263 11398 139309 11450
rect 139013 11396 139069 11398
rect 139093 11396 139149 11398
rect 139173 11396 139229 11398
rect 139253 11396 139309 11398
rect 138754 10804 138810 10840
rect 138754 10784 138756 10804
rect 138756 10784 138808 10804
rect 138808 10784 138810 10804
rect 139013 10362 139069 10364
rect 139093 10362 139149 10364
rect 139173 10362 139229 10364
rect 139253 10362 139309 10364
rect 139013 10310 139059 10362
rect 139059 10310 139069 10362
rect 139093 10310 139123 10362
rect 139123 10310 139135 10362
rect 139135 10310 139149 10362
rect 139173 10310 139187 10362
rect 139187 10310 139199 10362
rect 139199 10310 139229 10362
rect 139253 10310 139263 10362
rect 139263 10310 139309 10362
rect 139013 10308 139069 10310
rect 139093 10308 139149 10310
rect 139173 10308 139229 10310
rect 139253 10308 139309 10310
rect 138570 9560 138626 9616
rect 139306 9560 139362 9616
rect 138846 9288 138902 9344
rect 139013 9274 139069 9276
rect 139093 9274 139149 9276
rect 139173 9274 139229 9276
rect 139253 9274 139309 9276
rect 139013 9222 139059 9274
rect 139059 9222 139069 9274
rect 139093 9222 139123 9274
rect 139123 9222 139135 9274
rect 139135 9222 139149 9274
rect 139173 9222 139187 9274
rect 139187 9222 139199 9274
rect 139199 9222 139229 9274
rect 139253 9222 139263 9274
rect 139263 9222 139309 9274
rect 139013 9220 139069 9222
rect 139093 9220 139149 9222
rect 139173 9220 139229 9222
rect 139253 9220 139309 9222
rect 138386 6568 138442 6624
rect 138294 4140 138350 4176
rect 138294 4120 138296 4140
rect 138296 4120 138348 4140
rect 138348 4120 138350 4140
rect 139013 8186 139069 8188
rect 139093 8186 139149 8188
rect 139173 8186 139229 8188
rect 139253 8186 139309 8188
rect 139013 8134 139059 8186
rect 139059 8134 139069 8186
rect 139093 8134 139123 8186
rect 139123 8134 139135 8186
rect 139135 8134 139149 8186
rect 139173 8134 139187 8186
rect 139187 8134 139199 8186
rect 139199 8134 139229 8186
rect 139253 8134 139263 8186
rect 139263 8134 139309 8186
rect 139013 8132 139069 8134
rect 139093 8132 139149 8134
rect 139173 8132 139229 8134
rect 139253 8132 139309 8134
rect 139013 7098 139069 7100
rect 139093 7098 139149 7100
rect 139173 7098 139229 7100
rect 139253 7098 139309 7100
rect 139013 7046 139059 7098
rect 139059 7046 139069 7098
rect 139093 7046 139123 7098
rect 139123 7046 139135 7098
rect 139135 7046 139149 7098
rect 139173 7046 139187 7098
rect 139187 7046 139199 7098
rect 139199 7046 139229 7098
rect 139253 7046 139263 7098
rect 139263 7046 139309 7098
rect 139013 7044 139069 7046
rect 139093 7044 139149 7046
rect 139173 7044 139229 7046
rect 139253 7044 139309 7046
rect 139013 6010 139069 6012
rect 139093 6010 139149 6012
rect 139173 6010 139229 6012
rect 139253 6010 139309 6012
rect 139013 5958 139059 6010
rect 139059 5958 139069 6010
rect 139093 5958 139123 6010
rect 139123 5958 139135 6010
rect 139135 5958 139149 6010
rect 139173 5958 139187 6010
rect 139187 5958 139199 6010
rect 139199 5958 139229 6010
rect 139253 5958 139263 6010
rect 139263 5958 139309 6010
rect 139013 5956 139069 5958
rect 139093 5956 139149 5958
rect 139173 5956 139229 5958
rect 139253 5956 139309 5958
rect 139013 4922 139069 4924
rect 139093 4922 139149 4924
rect 139173 4922 139229 4924
rect 139253 4922 139309 4924
rect 139013 4870 139059 4922
rect 139059 4870 139069 4922
rect 139093 4870 139123 4922
rect 139123 4870 139135 4922
rect 139135 4870 139149 4922
rect 139173 4870 139187 4922
rect 139187 4870 139199 4922
rect 139199 4870 139229 4922
rect 139253 4870 139263 4922
rect 139263 4870 139309 4922
rect 139013 4868 139069 4870
rect 139093 4868 139149 4870
rect 139173 4868 139229 4870
rect 139253 4868 139309 4870
rect 139490 11328 139546 11384
rect 139490 8880 139546 8936
rect 139950 12416 140006 12472
rect 140594 12280 140650 12336
rect 139766 10376 139822 10432
rect 139858 10240 139914 10296
rect 139766 9696 139822 9752
rect 139858 9324 139860 9344
rect 139860 9324 139912 9344
rect 139912 9324 139914 9344
rect 139858 9288 139914 9324
rect 139674 7112 139730 7168
rect 139582 6024 139638 6080
rect 139490 5208 139546 5264
rect 139013 3834 139069 3836
rect 139093 3834 139149 3836
rect 139173 3834 139229 3836
rect 139253 3834 139309 3836
rect 139013 3782 139059 3834
rect 139059 3782 139069 3834
rect 139093 3782 139123 3834
rect 139123 3782 139135 3834
rect 139135 3782 139149 3834
rect 139173 3782 139187 3834
rect 139187 3782 139199 3834
rect 139199 3782 139229 3834
rect 139253 3782 139263 3834
rect 139263 3782 139309 3834
rect 139013 3780 139069 3782
rect 139093 3780 139149 3782
rect 139173 3780 139229 3782
rect 139253 3780 139309 3782
rect 139582 4972 139584 4992
rect 139584 4972 139636 4992
rect 139636 4972 139638 4992
rect 139582 4936 139638 4972
rect 140410 11056 140466 11112
rect 140042 9580 140098 9616
rect 140042 9560 140044 9580
rect 140044 9560 140096 9580
rect 140096 9560 140098 9580
rect 140042 4528 140098 4584
rect 139950 4120 140006 4176
rect 140134 4120 140190 4176
rect 141330 11328 141386 11384
rect 141238 10920 141294 10976
rect 141146 7656 141202 7712
rect 140778 7112 140834 7168
rect 140778 6604 140780 6624
rect 140780 6604 140832 6624
rect 140832 6604 140834 6624
rect 140778 6568 140834 6604
rect 140594 5092 140650 5128
rect 140594 5072 140596 5092
rect 140596 5072 140648 5092
rect 140648 5072 140650 5092
rect 140686 4392 140742 4448
rect 140686 3712 140742 3768
rect 139013 2746 139069 2748
rect 139093 2746 139149 2748
rect 139173 2746 139229 2748
rect 139253 2746 139309 2748
rect 139013 2694 139059 2746
rect 139059 2694 139069 2746
rect 139093 2694 139123 2746
rect 139123 2694 139135 2746
rect 139135 2694 139149 2746
rect 139173 2694 139187 2746
rect 139187 2694 139199 2746
rect 139199 2694 139229 2746
rect 139253 2694 139263 2746
rect 139263 2694 139309 2746
rect 139013 2692 139069 2694
rect 139093 2692 139149 2694
rect 139173 2692 139229 2694
rect 139253 2692 139309 2694
rect 140594 2352 140650 2408
rect 141514 11192 141570 11248
rect 141790 8608 141846 8664
rect 141330 7384 141386 7440
rect 141422 6840 141478 6896
rect 141146 6296 141202 6352
rect 141054 4528 141110 4584
rect 141054 2624 141110 2680
rect 141790 4004 141846 4040
rect 141790 3984 141792 4004
rect 141792 3984 141844 4004
rect 141844 3984 141846 4004
rect 143078 12008 143134 12064
rect 142618 11872 142674 11928
rect 142066 7928 142122 7984
rect 142066 7656 142122 7712
rect 141974 7384 142030 7440
rect 142066 7112 142122 7168
rect 142342 9288 142398 9344
rect 142342 6976 142398 7032
rect 142802 9832 142858 9888
rect 142802 9152 142858 9208
rect 143170 11600 143226 11656
rect 143262 11500 143264 11520
rect 143264 11500 143316 11520
rect 143316 11500 143318 11520
rect 143262 11464 143318 11500
rect 142250 6568 142306 6624
rect 142158 5888 142214 5944
rect 141974 5480 142030 5536
rect 143078 4256 143134 4312
rect 143998 14184 144054 14240
rect 143906 14048 143962 14104
rect 144274 12960 144330 13016
rect 144182 12280 144238 12336
rect 145654 13232 145710 13288
rect 145102 12552 145158 12608
rect 143446 11056 143502 11112
rect 143722 9324 143724 9344
rect 143724 9324 143776 9344
rect 143776 9324 143778 9344
rect 143722 9288 143778 9324
rect 143722 8744 143778 8800
rect 143998 9696 144054 9752
rect 144090 8744 144146 8800
rect 143814 7928 143870 7984
rect 143814 6332 143816 6352
rect 143816 6332 143868 6352
rect 143868 6332 143870 6352
rect 143814 6296 143870 6332
rect 143630 4256 143686 4312
rect 143630 3576 143686 3632
rect 141054 2216 141110 2272
rect 143722 2524 143724 2544
rect 143724 2524 143776 2544
rect 143776 2524 143778 2544
rect 143722 2488 143778 2524
rect 143722 1808 143778 1864
rect 144642 11192 144698 11248
rect 145010 11872 145066 11928
rect 145286 11328 145342 11384
rect 144734 10784 144790 10840
rect 144642 9696 144698 9752
rect 144182 6840 144238 6896
rect 144918 9696 144974 9752
rect 144826 8608 144882 8664
rect 144550 6296 144606 6352
rect 144918 7656 144974 7712
rect 144826 6976 144882 7032
rect 145010 6976 145066 7032
rect 144734 4120 144790 4176
rect 144918 4120 144974 4176
rect 145286 8880 145342 8936
rect 145838 13096 145894 13152
rect 145838 11600 145894 11656
rect 146206 13912 146262 13968
rect 147034 13640 147090 13696
rect 147586 13504 147642 13560
rect 146298 12688 146354 12744
rect 145562 9560 145618 9616
rect 145286 6976 145342 7032
rect 145194 5888 145250 5944
rect 145286 5480 145342 5536
rect 145562 8880 145618 8936
rect 145838 8064 145894 8120
rect 145654 7520 145710 7576
rect 145654 5888 145710 5944
rect 145562 4428 145564 4448
rect 145564 4428 145616 4448
rect 145616 4428 145618 4448
rect 145562 4392 145618 4428
rect 145562 4256 145618 4312
rect 145654 4120 145710 4176
rect 145470 3068 145472 3088
rect 145472 3068 145524 3088
rect 145524 3068 145526 3088
rect 145470 3032 145526 3068
rect 145010 1944 145066 2000
rect 145838 7520 145894 7576
rect 146206 9016 146262 9072
rect 145838 7112 145894 7168
rect 146022 4820 146078 4856
rect 146022 4800 146024 4820
rect 146024 4800 146076 4820
rect 146076 4800 146078 4820
rect 145930 4256 145986 4312
rect 145930 2216 145986 2272
rect 146482 6568 146538 6624
rect 146758 6568 146814 6624
rect 146298 4936 146354 4992
rect 146482 4936 146538 4992
rect 146206 3848 146262 3904
rect 146298 3732 146354 3768
rect 146298 3712 146300 3732
rect 146300 3712 146352 3732
rect 146352 3712 146354 3732
rect 147310 12280 147366 12336
rect 148046 13368 148102 13424
rect 148506 11872 148562 11928
rect 147678 11328 147734 11384
rect 148046 11328 148102 11384
rect 147770 11056 147826 11112
rect 147218 8064 147274 8120
rect 147402 8916 147404 8936
rect 147404 8916 147456 8936
rect 147456 8916 147458 8936
rect 147402 8880 147458 8916
rect 147770 8880 147826 8936
rect 147126 7112 147182 7168
rect 146942 6432 146998 6488
rect 147034 5888 147090 5944
rect 146942 5652 146944 5672
rect 146944 5652 146996 5672
rect 146996 5652 146998 5672
rect 146942 5616 146998 5652
rect 146942 5072 146998 5128
rect 146942 4428 146944 4448
rect 146944 4428 146996 4448
rect 146996 4428 146998 4448
rect 146942 4392 146998 4428
rect 147034 4120 147090 4176
rect 147678 6840 147734 6896
rect 148138 9016 148194 9072
rect 148322 10784 148378 10840
rect 148782 12960 148838 13016
rect 149242 11600 149298 11656
rect 148782 10804 148838 10840
rect 148782 10784 148784 10804
rect 148784 10784 148836 10804
rect 148836 10784 148838 10804
rect 148598 9832 148654 9888
rect 148690 9424 148746 9480
rect 148874 9424 148930 9480
rect 148782 9172 148838 9208
rect 148782 9152 148784 9172
rect 148784 9152 148836 9172
rect 148836 9152 148838 9172
rect 148690 8880 148746 8936
rect 148046 8200 148102 8256
rect 148046 7112 148102 7168
rect 147862 6160 147918 6216
rect 147310 5616 147366 5672
rect 147310 5072 147366 5128
rect 146942 3576 146998 3632
rect 147310 3304 147366 3360
rect 147954 4256 148010 4312
rect 147494 3576 147550 3632
rect 147678 3576 147734 3632
rect 147862 3304 147918 3360
rect 147862 3068 147864 3088
rect 147864 3068 147916 3088
rect 147916 3068 147918 3088
rect 147862 3032 147918 3068
rect 148322 5888 148378 5944
rect 148782 8744 148838 8800
rect 148230 5208 148286 5264
rect 148230 3460 148286 3496
rect 148230 3440 148232 3460
rect 148232 3440 148284 3460
rect 148284 3440 148286 3460
rect 149426 11600 149482 11656
rect 149426 10240 149482 10296
rect 149242 9152 149298 9208
rect 149150 8744 149206 8800
rect 149058 8608 149114 8664
rect 149058 8200 149114 8256
rect 148690 3304 148746 3360
rect 148874 3440 148930 3496
rect 148782 3032 148838 3088
rect 148506 2896 148562 2952
rect 148690 2796 148692 2816
rect 148692 2796 148744 2816
rect 148744 2796 148746 2816
rect 148690 2760 148746 2796
rect 150070 13096 150126 13152
rect 150438 11772 150440 11792
rect 150440 11772 150492 11792
rect 150492 11772 150494 11792
rect 150438 11736 150494 11772
rect 149610 8608 149666 8664
rect 149518 5652 149520 5672
rect 149520 5652 149572 5672
rect 149572 5652 149574 5672
rect 149518 5616 149574 5652
rect 150254 10240 150310 10296
rect 150070 9968 150126 10024
rect 150438 9968 150494 10024
rect 150622 11872 150678 11928
rect 150162 8608 150218 8664
rect 150162 8200 150218 8256
rect 150530 8608 150586 8664
rect 149886 6160 149942 6216
rect 149702 5616 149758 5672
rect 149058 3984 149114 4040
rect 149242 3984 149298 4040
rect 148138 1944 148194 2000
rect 149794 4392 149850 4448
rect 149702 3576 149758 3632
rect 149610 2488 149666 2544
rect 150254 6160 150310 6216
rect 150438 6296 150494 6352
rect 150070 3440 150126 3496
rect 149610 2080 149666 2136
rect 150438 3304 150494 3360
rect 150990 14320 151046 14376
rect 150806 12708 150862 12744
rect 150806 12688 150808 12708
rect 150808 12688 150860 12708
rect 150860 12688 150862 12708
rect 150898 8744 150954 8800
rect 150806 7540 150862 7576
rect 150806 7520 150808 7540
rect 150808 7520 150860 7540
rect 150860 7520 150862 7540
rect 150346 2080 150402 2136
rect 149242 1672 149298 1728
rect 151450 11600 151506 11656
rect 151266 9968 151322 10024
rect 151174 8880 151230 8936
rect 151082 8064 151138 8120
rect 151266 8064 151322 8120
rect 151082 7112 151138 7168
rect 150990 6160 151046 6216
rect 150898 4392 150954 4448
rect 151082 5208 151138 5264
rect 151082 3304 151138 3360
rect 151726 10376 151782 10432
rect 151542 6568 151598 6624
rect 151358 5208 151414 5264
rect 151266 4528 151322 4584
rect 152646 11464 152702 11520
rect 152370 11056 152426 11112
rect 152186 9868 152188 9888
rect 152188 9868 152240 9888
rect 152240 9868 152242 9888
rect 152186 9832 152242 9868
rect 152002 9560 152058 9616
rect 152002 8372 152004 8392
rect 152004 8372 152056 8392
rect 152056 8372 152058 8392
rect 152002 8336 152058 8372
rect 152002 7520 152058 7576
rect 152646 10648 152702 10704
rect 152554 9580 152610 9616
rect 152554 9560 152556 9580
rect 152556 9560 152608 9580
rect 152608 9560 152610 9580
rect 152370 8744 152426 8800
rect 151542 3460 151598 3496
rect 151542 3440 151544 3460
rect 151544 3440 151596 3460
rect 151596 3440 151598 3460
rect 152002 5344 152058 5400
rect 152370 6568 152426 6624
rect 152554 6568 152610 6624
rect 152462 6432 152518 6488
rect 152462 5480 152518 5536
rect 152278 5072 152334 5128
rect 152094 4664 152150 4720
rect 151818 2932 151820 2952
rect 151820 2932 151872 2952
rect 151872 2932 151874 2952
rect 151818 2896 151874 2932
rect 152922 12980 152978 13016
rect 152922 12960 152924 12980
rect 152924 12960 152976 12980
rect 152976 12960 152978 12980
rect 153198 13368 153254 13424
rect 154118 13232 154174 13288
rect 152922 12552 152978 12608
rect 152830 11056 152886 11112
rect 153106 12436 153162 12472
rect 153106 12416 153108 12436
rect 153108 12416 153160 12436
rect 153160 12416 153162 12436
rect 153382 12688 153438 12744
rect 153474 12008 153530 12064
rect 153290 9424 153346 9480
rect 153658 9424 153714 9480
rect 153566 8608 153622 8664
rect 154302 12688 154358 12744
rect 153842 10140 153844 10160
rect 153844 10140 153896 10160
rect 153896 10140 153898 10160
rect 153842 10104 153898 10140
rect 153106 8064 153162 8120
rect 153198 6840 153254 6896
rect 152922 4528 152978 4584
rect 152462 3476 152464 3496
rect 152464 3476 152516 3496
rect 152516 3476 152518 3496
rect 152462 3440 152518 3476
rect 152646 3440 152702 3496
rect 152830 3732 152886 3768
rect 152830 3712 152832 3732
rect 152832 3712 152884 3732
rect 152884 3712 152886 3732
rect 153014 3712 153070 3768
rect 153474 6704 153530 6760
rect 153566 6296 153622 6352
rect 153566 3984 153622 4040
rect 153474 3304 153530 3360
rect 153290 3168 153346 3224
rect 152370 2488 152426 2544
rect 153658 2352 153714 2408
rect 154670 11328 154726 11384
rect 154118 6976 154174 7032
rect 153934 6180 153990 6216
rect 153934 6160 153936 6180
rect 153936 6160 153988 6180
rect 153988 6160 153990 6180
rect 154026 2932 154028 2952
rect 154028 2932 154080 2952
rect 154080 2932 154082 2952
rect 154026 2896 154082 2932
rect 154302 8336 154358 8392
rect 154302 7404 154358 7440
rect 154302 7384 154304 7404
rect 154304 7384 154356 7404
rect 154356 7384 154358 7404
rect 154670 10240 154726 10296
rect 154670 10004 154672 10024
rect 154672 10004 154724 10024
rect 154724 10004 154726 10024
rect 154670 9968 154726 10004
rect 154578 8608 154634 8664
rect 154302 5480 154358 5536
rect 154302 5072 154358 5128
rect 154302 3304 154358 3360
rect 154762 6568 154818 6624
rect 154854 6296 154910 6352
rect 155866 13640 155922 13696
rect 155774 13504 155830 13560
rect 155314 11772 155316 11792
rect 155316 11772 155368 11792
rect 155368 11772 155370 11792
rect 155314 11736 155370 11772
rect 155222 10784 155278 10840
rect 154670 5752 154726 5808
rect 155222 8744 155278 8800
rect 155406 8336 155462 8392
rect 155222 6196 155224 6216
rect 155224 6196 155276 6216
rect 155276 6196 155278 6216
rect 155222 6160 155278 6196
rect 154486 3440 154542 3496
rect 155314 5888 155370 5944
rect 156694 12844 156750 12880
rect 156694 12824 156696 12844
rect 156696 12824 156748 12844
rect 156748 12824 156750 12844
rect 156326 12280 156382 12336
rect 156142 11756 156198 11792
rect 156142 11736 156144 11756
rect 156144 11736 156196 11756
rect 156196 11736 156198 11756
rect 156142 10512 156198 10568
rect 156050 9288 156106 9344
rect 155866 9152 155922 9208
rect 156142 9016 156198 9072
rect 155866 7692 155868 7712
rect 155868 7692 155920 7712
rect 155920 7692 155922 7712
rect 155866 7656 155922 7692
rect 155498 5652 155500 5672
rect 155500 5652 155552 5672
rect 155552 5652 155554 5672
rect 155498 5616 155554 5652
rect 154670 3712 154726 3768
rect 154670 3460 154726 3496
rect 154670 3440 154672 3460
rect 154672 3440 154724 3460
rect 154724 3440 154726 3460
rect 155498 5208 155554 5264
rect 155222 4256 155278 4312
rect 155130 4004 155186 4040
rect 155130 3984 155132 4004
rect 155132 3984 155184 4004
rect 155184 3984 155186 4004
rect 155038 3712 155094 3768
rect 155130 3476 155132 3496
rect 155132 3476 155184 3496
rect 155184 3476 155186 3496
rect 155130 3440 155186 3476
rect 154302 2624 154358 2680
rect 155958 7248 156014 7304
rect 155958 5616 156014 5672
rect 155774 3984 155830 4040
rect 156050 4800 156106 4856
rect 155958 2760 156014 2816
rect 155866 1944 155922 2000
rect 158735 13082 158791 13084
rect 158815 13082 158871 13084
rect 158895 13082 158951 13084
rect 158975 13082 159031 13084
rect 158735 13030 158781 13082
rect 158781 13030 158791 13082
rect 158815 13030 158845 13082
rect 158845 13030 158857 13082
rect 158857 13030 158871 13082
rect 158895 13030 158909 13082
rect 158909 13030 158921 13082
rect 158921 13030 158951 13082
rect 158975 13030 158985 13082
rect 158985 13030 159031 13082
rect 158735 13028 158791 13030
rect 158815 13028 158871 13030
rect 158895 13028 158951 13030
rect 158975 13028 159031 13030
rect 157062 11192 157118 11248
rect 156970 10920 157026 10976
rect 156878 9424 156934 9480
rect 156694 8608 156750 8664
rect 156602 7928 156658 7984
rect 156694 6024 156750 6080
rect 156786 5364 156842 5400
rect 156786 5344 156788 5364
rect 156788 5344 156840 5364
rect 156840 5344 156842 5364
rect 156970 8492 157026 8528
rect 156970 8472 156972 8492
rect 156972 8472 157024 8492
rect 157024 8472 157026 8492
rect 156970 7520 157026 7576
rect 156786 3884 156788 3904
rect 156788 3884 156840 3904
rect 156840 3884 156842 3904
rect 156786 3848 156842 3884
rect 157246 7112 157302 7168
rect 157062 5480 157118 5536
rect 157522 10004 157524 10024
rect 157524 10004 157576 10024
rect 157576 10004 157578 10024
rect 157522 9968 157578 10004
rect 157614 9696 157670 9752
rect 157614 4936 157670 4992
rect 153750 1128 153806 1184
rect 145746 992 145802 1048
rect 157614 3304 157670 3360
rect 158735 11994 158791 11996
rect 158815 11994 158871 11996
rect 158895 11994 158951 11996
rect 158975 11994 159031 11996
rect 158735 11942 158781 11994
rect 158781 11942 158791 11994
rect 158815 11942 158845 11994
rect 158845 11942 158857 11994
rect 158857 11942 158871 11994
rect 158895 11942 158909 11994
rect 158909 11942 158921 11994
rect 158921 11942 158951 11994
rect 158975 11942 158985 11994
rect 158985 11942 159031 11994
rect 158735 11940 158791 11942
rect 158815 11940 158871 11942
rect 158895 11940 158951 11942
rect 158975 11940 159031 11942
rect 158258 7928 158314 7984
rect 158074 3032 158130 3088
rect 158735 10906 158791 10908
rect 158815 10906 158871 10908
rect 158895 10906 158951 10908
rect 158975 10906 159031 10908
rect 158735 10854 158781 10906
rect 158781 10854 158791 10906
rect 158815 10854 158845 10906
rect 158845 10854 158857 10906
rect 158857 10854 158871 10906
rect 158895 10854 158909 10906
rect 158909 10854 158921 10906
rect 158921 10854 158951 10906
rect 158975 10854 158985 10906
rect 158985 10854 159031 10906
rect 158735 10852 158791 10854
rect 158815 10852 158871 10854
rect 158895 10852 158951 10854
rect 158975 10852 159031 10854
rect 158735 9818 158791 9820
rect 158815 9818 158871 9820
rect 158895 9818 158951 9820
rect 158975 9818 159031 9820
rect 158735 9766 158781 9818
rect 158781 9766 158791 9818
rect 158815 9766 158845 9818
rect 158845 9766 158857 9818
rect 158857 9766 158871 9818
rect 158895 9766 158909 9818
rect 158909 9766 158921 9818
rect 158921 9766 158951 9818
rect 158975 9766 158985 9818
rect 158985 9766 159031 9818
rect 158735 9764 158791 9766
rect 158815 9764 158871 9766
rect 158895 9764 158951 9766
rect 158975 9764 159031 9766
rect 158735 8730 158791 8732
rect 158815 8730 158871 8732
rect 158895 8730 158951 8732
rect 158975 8730 159031 8732
rect 158735 8678 158781 8730
rect 158781 8678 158791 8730
rect 158815 8678 158845 8730
rect 158845 8678 158857 8730
rect 158857 8678 158871 8730
rect 158895 8678 158909 8730
rect 158909 8678 158921 8730
rect 158921 8678 158951 8730
rect 158975 8678 158985 8730
rect 158985 8678 159031 8730
rect 158735 8676 158791 8678
rect 158815 8676 158871 8678
rect 158895 8676 158951 8678
rect 158975 8676 159031 8678
rect 158735 7642 158791 7644
rect 158815 7642 158871 7644
rect 158895 7642 158951 7644
rect 158975 7642 159031 7644
rect 158735 7590 158781 7642
rect 158781 7590 158791 7642
rect 158815 7590 158845 7642
rect 158845 7590 158857 7642
rect 158857 7590 158871 7642
rect 158895 7590 158909 7642
rect 158909 7590 158921 7642
rect 158921 7590 158951 7642
rect 158975 7590 158985 7642
rect 158985 7590 159031 7642
rect 158735 7588 158791 7590
rect 158815 7588 158871 7590
rect 158895 7588 158951 7590
rect 158975 7588 159031 7590
rect 158735 6554 158791 6556
rect 158815 6554 158871 6556
rect 158895 6554 158951 6556
rect 158975 6554 159031 6556
rect 158735 6502 158781 6554
rect 158781 6502 158791 6554
rect 158815 6502 158845 6554
rect 158845 6502 158857 6554
rect 158857 6502 158871 6554
rect 158895 6502 158909 6554
rect 158909 6502 158921 6554
rect 158921 6502 158951 6554
rect 158975 6502 158985 6554
rect 158985 6502 159031 6554
rect 158735 6500 158791 6502
rect 158815 6500 158871 6502
rect 158895 6500 158951 6502
rect 158975 6500 159031 6502
rect 158735 5466 158791 5468
rect 158815 5466 158871 5468
rect 158895 5466 158951 5468
rect 158975 5466 159031 5468
rect 158735 5414 158781 5466
rect 158781 5414 158791 5466
rect 158815 5414 158845 5466
rect 158845 5414 158857 5466
rect 158857 5414 158871 5466
rect 158895 5414 158909 5466
rect 158909 5414 158921 5466
rect 158921 5414 158951 5466
rect 158975 5414 158985 5466
rect 158985 5414 159031 5466
rect 158735 5412 158791 5414
rect 158815 5412 158871 5414
rect 158895 5412 158951 5414
rect 158975 5412 159031 5414
rect 158735 4378 158791 4380
rect 158815 4378 158871 4380
rect 158895 4378 158951 4380
rect 158975 4378 159031 4380
rect 158735 4326 158781 4378
rect 158781 4326 158791 4378
rect 158815 4326 158845 4378
rect 158845 4326 158857 4378
rect 158857 4326 158871 4378
rect 158895 4326 158909 4378
rect 158909 4326 158921 4378
rect 158921 4326 158951 4378
rect 158975 4326 158985 4378
rect 158985 4326 159031 4378
rect 158735 4324 158791 4326
rect 158815 4324 158871 4326
rect 158895 4324 158951 4326
rect 158975 4324 159031 4326
rect 158735 3290 158791 3292
rect 158815 3290 158871 3292
rect 158895 3290 158951 3292
rect 158975 3290 159031 3292
rect 158735 3238 158781 3290
rect 158781 3238 158791 3290
rect 158815 3238 158845 3290
rect 158845 3238 158857 3290
rect 158857 3238 158871 3290
rect 158895 3238 158909 3290
rect 158909 3238 158921 3290
rect 158921 3238 158951 3290
rect 158975 3238 158985 3290
rect 158985 3238 159031 3290
rect 158735 3236 158791 3238
rect 158815 3236 158871 3238
rect 158895 3236 158951 3238
rect 158975 3236 159031 3238
rect 159270 10240 159326 10296
rect 158166 2216 158222 2272
rect 158735 2202 158791 2204
rect 158815 2202 158871 2204
rect 158895 2202 158951 2204
rect 158975 2202 159031 2204
rect 158735 2150 158781 2202
rect 158781 2150 158791 2202
rect 158815 2150 158845 2202
rect 158845 2150 158857 2202
rect 158857 2150 158871 2202
rect 158895 2150 158909 2202
rect 158909 2150 158921 2202
rect 158921 2150 158951 2202
rect 158975 2150 158985 2202
rect 158985 2150 159031 2202
rect 158735 2148 158791 2150
rect 158815 2148 158871 2150
rect 158895 2148 158951 2150
rect 158975 2148 159031 2150
rect 157798 2080 157854 2136
rect 156418 992 156474 1048
<< metal3 >>
rect 125685 14514 125751 14517
rect 150750 14514 150756 14516
rect 125685 14512 150756 14514
rect 125685 14456 125690 14512
rect 125746 14456 150756 14512
rect 125685 14454 150756 14456
rect 125685 14451 125751 14454
rect 150750 14452 150756 14454
rect 150820 14452 150826 14516
rect 128445 14378 128511 14381
rect 150985 14378 151051 14381
rect 128445 14376 151051 14378
rect 128445 14320 128450 14376
rect 128506 14320 150990 14376
rect 151046 14320 151051 14376
rect 128445 14318 151051 14320
rect 128445 14315 128511 14318
rect 150985 14315 151051 14318
rect 143993 14242 144059 14245
rect 156822 14242 156828 14244
rect 143993 14240 156828 14242
rect 143993 14184 143998 14240
rect 144054 14184 156828 14240
rect 143993 14182 156828 14184
rect 143993 14179 144059 14182
rect 156822 14180 156828 14182
rect 156892 14180 156898 14244
rect 121361 14106 121427 14109
rect 136909 14106 136975 14109
rect 121361 14104 136975 14106
rect 121361 14048 121366 14104
rect 121422 14048 136914 14104
rect 136970 14048 136975 14104
rect 121361 14046 136975 14048
rect 121361 14043 121427 14046
rect 136909 14043 136975 14046
rect 143901 14106 143967 14109
rect 155718 14106 155724 14108
rect 143901 14104 155724 14106
rect 143901 14048 143906 14104
rect 143962 14048 155724 14104
rect 143901 14046 155724 14048
rect 143901 14043 143967 14046
rect 155718 14044 155724 14046
rect 155788 14044 155794 14108
rect 146201 13970 146267 13973
rect 155166 13970 155172 13972
rect 146201 13968 155172 13970
rect 146201 13912 146206 13968
rect 146262 13912 155172 13968
rect 146201 13910 155172 13912
rect 146201 13907 146267 13910
rect 155166 13908 155172 13910
rect 155236 13908 155242 13972
rect 0 13834 800 13864
rect 4061 13834 4127 13837
rect 0 13832 4127 13834
rect 0 13776 4066 13832
rect 4122 13776 4127 13832
rect 0 13774 4127 13776
rect 0 13744 800 13774
rect 4061 13771 4127 13774
rect 116945 13698 117011 13701
rect 138657 13698 138723 13701
rect 116945 13696 138723 13698
rect 116945 13640 116950 13696
rect 117006 13640 138662 13696
rect 138718 13640 138723 13696
rect 116945 13638 138723 13640
rect 116945 13635 117011 13638
rect 138657 13635 138723 13638
rect 147029 13698 147095 13701
rect 155861 13698 155927 13701
rect 147029 13696 155927 13698
rect 147029 13640 147034 13696
rect 147090 13640 155866 13696
rect 155922 13640 155927 13696
rect 147029 13638 155927 13640
rect 147029 13635 147095 13638
rect 155861 13635 155927 13638
rect 20668 13632 20984 13633
rect 20668 13568 20674 13632
rect 20738 13568 20754 13632
rect 20818 13568 20834 13632
rect 20898 13568 20914 13632
rect 20978 13568 20984 13632
rect 20668 13567 20984 13568
rect 60113 13632 60429 13633
rect 60113 13568 60119 13632
rect 60183 13568 60199 13632
rect 60263 13568 60279 13632
rect 60343 13568 60359 13632
rect 60423 13568 60429 13632
rect 60113 13567 60429 13568
rect 99558 13632 99874 13633
rect 99558 13568 99564 13632
rect 99628 13568 99644 13632
rect 99708 13568 99724 13632
rect 99788 13568 99804 13632
rect 99868 13568 99874 13632
rect 99558 13567 99874 13568
rect 139003 13632 139319 13633
rect 139003 13568 139009 13632
rect 139073 13568 139089 13632
rect 139153 13568 139169 13632
rect 139233 13568 139249 13632
rect 139313 13568 139319 13632
rect 139003 13567 139319 13568
rect 77477 13562 77543 13565
rect 82169 13562 82235 13565
rect 77477 13560 82235 13562
rect 77477 13504 77482 13560
rect 77538 13504 82174 13560
rect 82230 13504 82235 13560
rect 77477 13502 82235 13504
rect 77477 13499 77543 13502
rect 82169 13499 82235 13502
rect 147581 13562 147647 13565
rect 155769 13562 155835 13565
rect 147581 13560 155835 13562
rect 147581 13504 147586 13560
rect 147642 13504 155774 13560
rect 155830 13504 155835 13560
rect 147581 13502 155835 13504
rect 147581 13499 147647 13502
rect 155769 13499 155835 13502
rect 43989 13426 44055 13429
rect 49785 13426 49851 13429
rect 43989 13424 49851 13426
rect 43989 13368 43994 13424
rect 44050 13368 49790 13424
rect 49846 13368 49851 13424
rect 43989 13366 49851 13368
rect 43989 13363 44055 13366
rect 49785 13363 49851 13366
rect 59445 13426 59511 13429
rect 95877 13426 95943 13429
rect 59445 13424 95943 13426
rect 59445 13368 59450 13424
rect 59506 13368 95882 13424
rect 95938 13368 95943 13424
rect 59445 13366 95943 13368
rect 59445 13363 59511 13366
rect 95877 13363 95943 13366
rect 148041 13426 148107 13429
rect 153193 13426 153259 13429
rect 148041 13424 153259 13426
rect 148041 13368 148046 13424
rect 148102 13368 153198 13424
rect 153254 13368 153259 13424
rect 148041 13366 153259 13368
rect 148041 13363 148107 13366
rect 153193 13363 153259 13366
rect 10225 13290 10291 13293
rect 16389 13290 16455 13293
rect 10225 13288 16455 13290
rect 10225 13232 10230 13288
rect 10286 13232 16394 13288
rect 16450 13232 16455 13288
rect 10225 13230 16455 13232
rect 10225 13227 10291 13230
rect 16389 13227 16455 13230
rect 30097 13290 30163 13293
rect 31753 13290 31819 13293
rect 30097 13288 31819 13290
rect 30097 13232 30102 13288
rect 30158 13232 31758 13288
rect 31814 13232 31819 13288
rect 30097 13230 31819 13232
rect 30097 13227 30163 13230
rect 31753 13227 31819 13230
rect 56317 13290 56383 13293
rect 56685 13290 56751 13293
rect 56317 13288 56751 13290
rect 56317 13232 56322 13288
rect 56378 13232 56690 13288
rect 56746 13232 56751 13288
rect 56317 13230 56751 13232
rect 56317 13227 56383 13230
rect 56685 13227 56751 13230
rect 60365 13290 60431 13293
rect 63677 13290 63743 13293
rect 60365 13288 63743 13290
rect 60365 13232 60370 13288
rect 60426 13232 63682 13288
rect 63738 13232 63743 13288
rect 60365 13230 63743 13232
rect 60365 13227 60431 13230
rect 63677 13227 63743 13230
rect 79961 13290 80027 13293
rect 81525 13290 81591 13293
rect 89253 13290 89319 13293
rect 79961 13288 81591 13290
rect 79961 13232 79966 13288
rect 80022 13232 81530 13288
rect 81586 13232 81591 13288
rect 79961 13230 81591 13232
rect 79961 13227 80027 13230
rect 81525 13227 81591 13230
rect 86910 13288 89319 13290
rect 86910 13232 89258 13288
rect 89314 13232 89319 13288
rect 86910 13230 89319 13232
rect 21357 13154 21423 13157
rect 27981 13154 28047 13157
rect 21357 13152 28047 13154
rect 21357 13096 21362 13152
rect 21418 13096 27986 13152
rect 28042 13096 28047 13152
rect 21357 13094 28047 13096
rect 21357 13091 21423 13094
rect 27981 13091 28047 13094
rect 55397 13154 55463 13157
rect 60641 13154 60707 13157
rect 55397 13152 60707 13154
rect 55397 13096 55402 13152
rect 55458 13096 60646 13152
rect 60702 13096 60707 13152
rect 55397 13094 60707 13096
rect 55397 13091 55463 13094
rect 60641 13091 60707 13094
rect 69657 13154 69723 13157
rect 76833 13154 76899 13157
rect 69657 13152 76899 13154
rect 69657 13096 69662 13152
rect 69718 13096 76838 13152
rect 76894 13096 76899 13152
rect 69657 13094 76899 13096
rect 69657 13091 69723 13094
rect 76833 13091 76899 13094
rect 80237 13154 80303 13157
rect 86910 13154 86970 13230
rect 89253 13227 89319 13230
rect 96981 13290 97047 13293
rect 99925 13290 99991 13293
rect 96981 13288 99991 13290
rect 96981 13232 96986 13288
rect 97042 13232 99930 13288
rect 99986 13232 99991 13288
rect 96981 13230 99991 13232
rect 96981 13227 97047 13230
rect 99925 13227 99991 13230
rect 121453 13290 121519 13293
rect 124765 13290 124831 13293
rect 121453 13288 124831 13290
rect 121453 13232 121458 13288
rect 121514 13232 124770 13288
rect 124826 13232 124831 13288
rect 121453 13230 124831 13232
rect 121453 13227 121519 13230
rect 124765 13227 124831 13230
rect 125317 13290 125383 13293
rect 129549 13290 129615 13293
rect 125317 13288 129615 13290
rect 125317 13232 125322 13288
rect 125378 13232 129554 13288
rect 129610 13232 129615 13288
rect 125317 13230 129615 13232
rect 125317 13227 125383 13230
rect 129549 13227 129615 13230
rect 130377 13290 130443 13293
rect 133137 13290 133203 13293
rect 130377 13288 133203 13290
rect 130377 13232 130382 13288
rect 130438 13232 133142 13288
rect 133198 13232 133203 13288
rect 130377 13230 133203 13232
rect 130377 13227 130443 13230
rect 133137 13227 133203 13230
rect 145649 13290 145715 13293
rect 154113 13290 154179 13293
rect 145649 13288 154179 13290
rect 145649 13232 145654 13288
rect 145710 13232 154118 13288
rect 154174 13232 154179 13288
rect 145649 13230 154179 13232
rect 145649 13227 145715 13230
rect 154113 13227 154179 13230
rect 80237 13152 86970 13154
rect 80237 13096 80242 13152
rect 80298 13096 86970 13152
rect 80237 13094 86970 13096
rect 88885 13154 88951 13157
rect 94405 13154 94471 13157
rect 88885 13152 94471 13154
rect 88885 13096 88890 13152
rect 88946 13096 94410 13152
rect 94466 13096 94471 13152
rect 88885 13094 94471 13096
rect 80237 13091 80303 13094
rect 88885 13091 88951 13094
rect 94405 13091 94471 13094
rect 97717 13154 97783 13157
rect 100293 13154 100359 13157
rect 97717 13152 100359 13154
rect 97717 13096 97722 13152
rect 97778 13096 100298 13152
rect 100354 13096 100359 13152
rect 97717 13094 100359 13096
rect 97717 13091 97783 13094
rect 100293 13091 100359 13094
rect 110413 13154 110479 13157
rect 113081 13154 113147 13157
rect 110413 13152 113147 13154
rect 110413 13096 110418 13152
rect 110474 13096 113086 13152
rect 113142 13096 113147 13152
rect 110413 13094 113147 13096
rect 110413 13091 110479 13094
rect 113081 13091 113147 13094
rect 122373 13154 122439 13157
rect 124397 13154 124463 13157
rect 122373 13152 124463 13154
rect 122373 13096 122378 13152
rect 122434 13096 124402 13152
rect 124458 13096 124463 13152
rect 122373 13094 124463 13096
rect 122373 13091 122439 13094
rect 124397 13091 124463 13094
rect 145833 13154 145899 13157
rect 150065 13154 150131 13157
rect 145833 13152 150131 13154
rect 145833 13096 145838 13152
rect 145894 13096 150070 13152
rect 150126 13096 150131 13152
rect 145833 13094 150131 13096
rect 145833 13091 145899 13094
rect 150065 13091 150131 13094
rect 40390 13088 40706 13089
rect 40390 13024 40396 13088
rect 40460 13024 40476 13088
rect 40540 13024 40556 13088
rect 40620 13024 40636 13088
rect 40700 13024 40706 13088
rect 40390 13023 40706 13024
rect 79835 13088 80151 13089
rect 79835 13024 79841 13088
rect 79905 13024 79921 13088
rect 79985 13024 80001 13088
rect 80065 13024 80081 13088
rect 80145 13024 80151 13088
rect 79835 13023 80151 13024
rect 119280 13088 119596 13089
rect 119280 13024 119286 13088
rect 119350 13024 119366 13088
rect 119430 13024 119446 13088
rect 119510 13024 119526 13088
rect 119590 13024 119596 13088
rect 119280 13023 119596 13024
rect 158725 13088 159041 13089
rect 158725 13024 158731 13088
rect 158795 13024 158811 13088
rect 158875 13024 158891 13088
rect 158955 13024 158971 13088
rect 159035 13024 159041 13088
rect 158725 13023 159041 13024
rect 50889 13018 50955 13021
rect 51165 13018 51231 13021
rect 50889 13016 51231 13018
rect 50889 12960 50894 13016
rect 50950 12960 51170 13016
rect 51226 12960 51231 13016
rect 50889 12958 51231 12960
rect 50889 12955 50955 12958
rect 51165 12955 51231 12958
rect 58617 13018 58683 13021
rect 60825 13018 60891 13021
rect 58617 13016 60891 13018
rect 58617 12960 58622 13016
rect 58678 12960 60830 13016
rect 60886 12960 60891 13016
rect 58617 12958 60891 12960
rect 58617 12955 58683 12958
rect 60825 12955 60891 12958
rect 77385 13018 77451 13021
rect 79501 13018 79567 13021
rect 77385 13016 79567 13018
rect 77385 12960 77390 13016
rect 77446 12960 79506 13016
rect 79562 12960 79567 13016
rect 77385 12958 79567 12960
rect 77385 12955 77451 12958
rect 79501 12955 79567 12958
rect 120901 13018 120967 13021
rect 126329 13018 126395 13021
rect 120901 13016 126395 13018
rect 120901 12960 120906 13016
rect 120962 12960 126334 13016
rect 126390 12960 126395 13016
rect 120901 12958 126395 12960
rect 120901 12955 120967 12958
rect 126329 12955 126395 12958
rect 127341 13018 127407 13021
rect 131297 13018 131363 13021
rect 127341 13016 131363 13018
rect 127341 12960 127346 13016
rect 127402 12960 131302 13016
rect 131358 12960 131363 13016
rect 127341 12958 131363 12960
rect 127341 12955 127407 12958
rect 131297 12955 131363 12958
rect 144269 13018 144335 13021
rect 148777 13018 148843 13021
rect 144269 13016 148843 13018
rect 144269 12960 144274 13016
rect 144330 12960 148782 13016
rect 148838 12960 148843 13016
rect 144269 12958 148843 12960
rect 144269 12955 144335 12958
rect 148777 12955 148843 12958
rect 149646 12956 149652 13020
rect 149716 13018 149722 13020
rect 152917 13018 152983 13021
rect 149716 13016 152983 13018
rect 149716 12960 152922 13016
rect 152978 12960 152983 13016
rect 149716 12958 152983 12960
rect 149716 12956 149722 12958
rect 152917 12955 152983 12958
rect 22737 12882 22803 12885
rect 30649 12882 30715 12885
rect 22737 12880 30715 12882
rect 22737 12824 22742 12880
rect 22798 12824 30654 12880
rect 30710 12824 30715 12880
rect 22737 12822 30715 12824
rect 22737 12819 22803 12822
rect 30649 12819 30715 12822
rect 50705 12882 50771 12885
rect 56041 12882 56107 12885
rect 115657 12882 115723 12885
rect 50705 12880 115723 12882
rect 50705 12824 50710 12880
rect 50766 12824 56046 12880
rect 56102 12824 115662 12880
rect 115718 12824 115723 12880
rect 50705 12822 115723 12824
rect 50705 12819 50771 12822
rect 56041 12819 56107 12822
rect 115657 12819 115723 12822
rect 120809 12882 120875 12885
rect 124857 12882 124923 12885
rect 120809 12880 124923 12882
rect 120809 12824 120814 12880
rect 120870 12824 124862 12880
rect 124918 12824 124923 12880
rect 120809 12822 124923 12824
rect 120809 12819 120875 12822
rect 124857 12819 124923 12822
rect 128629 12882 128695 12885
rect 134885 12882 134951 12885
rect 156689 12882 156755 12885
rect 128629 12880 133890 12882
rect 128629 12824 128634 12880
rect 128690 12824 133890 12880
rect 128629 12822 133890 12824
rect 128629 12819 128695 12822
rect 21541 12746 21607 12749
rect 24025 12746 24091 12749
rect 21541 12744 24091 12746
rect 21541 12688 21546 12744
rect 21602 12688 24030 12744
rect 24086 12688 24091 12744
rect 21541 12686 24091 12688
rect 21541 12683 21607 12686
rect 24025 12683 24091 12686
rect 26233 12746 26299 12749
rect 29729 12746 29795 12749
rect 26233 12744 29795 12746
rect 26233 12688 26238 12744
rect 26294 12688 29734 12744
rect 29790 12688 29795 12744
rect 26233 12686 29795 12688
rect 26233 12683 26299 12686
rect 29729 12683 29795 12686
rect 41689 12746 41755 12749
rect 46289 12746 46355 12749
rect 41689 12744 46355 12746
rect 41689 12688 41694 12744
rect 41750 12688 46294 12744
rect 46350 12688 46355 12744
rect 41689 12686 46355 12688
rect 41689 12683 41755 12686
rect 46289 12683 46355 12686
rect 66161 12746 66227 12749
rect 93393 12746 93459 12749
rect 66161 12744 93459 12746
rect 66161 12688 66166 12744
rect 66222 12688 93398 12744
rect 93454 12688 93459 12744
rect 66161 12686 93459 12688
rect 66161 12683 66227 12686
rect 93393 12683 93459 12686
rect 103881 12746 103947 12749
rect 133137 12746 133203 12749
rect 103881 12744 133203 12746
rect 103881 12688 103886 12744
rect 103942 12688 133142 12744
rect 133198 12688 133203 12744
rect 103881 12686 133203 12688
rect 133830 12746 133890 12822
rect 134885 12880 156755 12882
rect 134885 12824 134890 12880
rect 134946 12824 156694 12880
rect 156750 12824 156755 12880
rect 134885 12822 156755 12824
rect 134885 12819 134951 12822
rect 156689 12819 156755 12822
rect 134333 12746 134399 12749
rect 135713 12746 135779 12749
rect 133830 12744 135779 12746
rect 133830 12688 134338 12744
rect 134394 12688 135718 12744
rect 135774 12688 135779 12744
rect 133830 12686 135779 12688
rect 103881 12683 103947 12686
rect 133137 12683 133203 12686
rect 134333 12683 134399 12686
rect 135713 12683 135779 12686
rect 146293 12746 146359 12749
rect 150801 12746 150867 12749
rect 146293 12744 150867 12746
rect 146293 12688 146298 12744
rect 146354 12688 150806 12744
rect 150862 12688 150867 12744
rect 146293 12686 150867 12688
rect 146293 12683 146359 12686
rect 150801 12683 150867 12686
rect 153377 12746 153443 12749
rect 154297 12746 154363 12749
rect 153377 12744 154363 12746
rect 153377 12688 153382 12744
rect 153438 12688 154302 12744
rect 154358 12688 154363 12744
rect 153377 12686 154363 12688
rect 153377 12683 153443 12686
rect 154297 12683 154363 12686
rect 74809 12610 74875 12613
rect 88977 12610 89043 12613
rect 74809 12608 89043 12610
rect 74809 12552 74814 12608
rect 74870 12552 88982 12608
rect 89038 12552 89043 12608
rect 74809 12550 89043 12552
rect 74809 12547 74875 12550
rect 88977 12547 89043 12550
rect 116117 12610 116183 12613
rect 136725 12610 136791 12613
rect 116117 12608 136791 12610
rect 116117 12552 116122 12608
rect 116178 12552 136730 12608
rect 136786 12552 136791 12608
rect 116117 12550 136791 12552
rect 116117 12547 116183 12550
rect 136725 12547 136791 12550
rect 145097 12610 145163 12613
rect 152917 12610 152983 12613
rect 145097 12608 152983 12610
rect 145097 12552 145102 12608
rect 145158 12552 152922 12608
rect 152978 12552 152983 12608
rect 145097 12550 152983 12552
rect 145097 12547 145163 12550
rect 152917 12547 152983 12550
rect 20668 12544 20984 12545
rect 20668 12480 20674 12544
rect 20738 12480 20754 12544
rect 20818 12480 20834 12544
rect 20898 12480 20914 12544
rect 20978 12480 20984 12544
rect 20668 12479 20984 12480
rect 60113 12544 60429 12545
rect 60113 12480 60119 12544
rect 60183 12480 60199 12544
rect 60263 12480 60279 12544
rect 60343 12480 60359 12544
rect 60423 12480 60429 12544
rect 60113 12479 60429 12480
rect 99558 12544 99874 12545
rect 99558 12480 99564 12544
rect 99628 12480 99644 12544
rect 99708 12480 99724 12544
rect 99788 12480 99804 12544
rect 99868 12480 99874 12544
rect 99558 12479 99874 12480
rect 139003 12544 139319 12545
rect 139003 12480 139009 12544
rect 139073 12480 139089 12544
rect 139153 12480 139169 12544
rect 139233 12480 139249 12544
rect 139313 12480 139319 12544
rect 139003 12479 139319 12480
rect 45553 12474 45619 12477
rect 46933 12474 46999 12477
rect 45553 12472 46999 12474
rect 45553 12416 45558 12472
rect 45614 12416 46938 12472
rect 46994 12416 46999 12472
rect 45553 12414 46999 12416
rect 45553 12411 45619 12414
rect 46933 12411 46999 12414
rect 77293 12474 77359 12477
rect 80237 12474 80303 12477
rect 77293 12472 80303 12474
rect 77293 12416 77298 12472
rect 77354 12416 80242 12472
rect 80298 12416 80303 12472
rect 77293 12414 80303 12416
rect 77293 12411 77359 12414
rect 80237 12411 80303 12414
rect 81341 12474 81407 12477
rect 83181 12474 83247 12477
rect 81341 12472 83247 12474
rect 81341 12416 81346 12472
rect 81402 12416 83186 12472
rect 83242 12416 83247 12472
rect 81341 12414 83247 12416
rect 81341 12411 81407 12414
rect 83181 12411 83247 12414
rect 110413 12474 110479 12477
rect 120257 12474 120323 12477
rect 110413 12472 120323 12474
rect 110413 12416 110418 12472
rect 110474 12416 120262 12472
rect 120318 12416 120323 12472
rect 110413 12414 120323 12416
rect 110413 12411 110479 12414
rect 120257 12411 120323 12414
rect 123293 12474 123359 12477
rect 136633 12474 136699 12477
rect 123293 12472 136699 12474
rect 123293 12416 123298 12472
rect 123354 12416 136638 12472
rect 136694 12416 136699 12472
rect 123293 12414 136699 12416
rect 123293 12411 123359 12414
rect 136633 12411 136699 12414
rect 139945 12474 140011 12477
rect 153101 12474 153167 12477
rect 139945 12472 153167 12474
rect 139945 12416 139950 12472
rect 140006 12416 153106 12472
rect 153162 12416 153167 12472
rect 139945 12414 153167 12416
rect 139945 12411 140011 12414
rect 153101 12411 153167 12414
rect 12065 12338 12131 12341
rect 12433 12338 12499 12341
rect 12065 12336 12499 12338
rect 12065 12280 12070 12336
rect 12126 12280 12438 12336
rect 12494 12280 12499 12336
rect 12065 12278 12499 12280
rect 12065 12275 12131 12278
rect 12433 12275 12499 12278
rect 40217 12338 40283 12341
rect 40861 12338 40927 12341
rect 40217 12336 40927 12338
rect 40217 12280 40222 12336
rect 40278 12280 40866 12336
rect 40922 12280 40927 12336
rect 40217 12278 40927 12280
rect 40217 12275 40283 12278
rect 40861 12275 40927 12278
rect 42149 12338 42215 12341
rect 46749 12338 46815 12341
rect 42149 12336 46815 12338
rect 42149 12280 42154 12336
rect 42210 12280 46754 12336
rect 46810 12280 46815 12336
rect 42149 12278 46815 12280
rect 42149 12275 42215 12278
rect 46749 12275 46815 12278
rect 50889 12338 50955 12341
rect 55949 12338 56015 12341
rect 50889 12336 56015 12338
rect 50889 12280 50894 12336
rect 50950 12280 55954 12336
rect 56010 12280 56015 12336
rect 50889 12278 56015 12280
rect 50889 12275 50955 12278
rect 55949 12275 56015 12278
rect 57145 12338 57211 12341
rect 58801 12338 58867 12341
rect 57145 12336 58867 12338
rect 57145 12280 57150 12336
rect 57206 12280 58806 12336
rect 58862 12280 58867 12336
rect 57145 12278 58867 12280
rect 57145 12275 57211 12278
rect 58801 12275 58867 12278
rect 78581 12338 78647 12341
rect 81893 12338 81959 12341
rect 78581 12336 81959 12338
rect 78581 12280 78586 12336
rect 78642 12280 81898 12336
rect 81954 12280 81959 12336
rect 78581 12278 81959 12280
rect 78581 12275 78647 12278
rect 81893 12275 81959 12278
rect 82077 12338 82143 12341
rect 85481 12338 85547 12341
rect 82077 12336 85547 12338
rect 82077 12280 82082 12336
rect 82138 12280 85486 12336
rect 85542 12280 85547 12336
rect 82077 12278 85547 12280
rect 82077 12275 82143 12278
rect 85481 12275 85547 12278
rect 96797 12338 96863 12341
rect 127157 12338 127223 12341
rect 130193 12338 130259 12341
rect 96797 12336 130259 12338
rect 96797 12280 96802 12336
rect 96858 12280 127162 12336
rect 127218 12280 130198 12336
rect 130254 12280 130259 12336
rect 96797 12278 130259 12280
rect 96797 12275 96863 12278
rect 127157 12275 127223 12278
rect 130193 12275 130259 12278
rect 136909 12338 136975 12341
rect 140589 12338 140655 12341
rect 136909 12336 140655 12338
rect 136909 12280 136914 12336
rect 136970 12280 140594 12336
rect 140650 12280 140655 12336
rect 136909 12278 140655 12280
rect 136909 12275 136975 12278
rect 140589 12275 140655 12278
rect 144177 12338 144243 12341
rect 147305 12338 147371 12341
rect 156321 12338 156387 12341
rect 144177 12336 147371 12338
rect 144177 12280 144182 12336
rect 144238 12280 147310 12336
rect 147366 12280 147371 12336
rect 144177 12278 147371 12280
rect 144177 12275 144243 12278
rect 147305 12275 147371 12278
rect 147630 12336 156387 12338
rect 147630 12280 156326 12336
rect 156382 12280 156387 12336
rect 147630 12278 156387 12280
rect 9857 12202 9923 12205
rect 14825 12202 14891 12205
rect 17953 12202 18019 12205
rect 9857 12200 18019 12202
rect 9857 12144 9862 12200
rect 9918 12144 14830 12200
rect 14886 12144 17958 12200
rect 18014 12144 18019 12200
rect 9857 12142 18019 12144
rect 9857 12139 9923 12142
rect 14825 12139 14891 12142
rect 17953 12139 18019 12142
rect 45461 12202 45527 12205
rect 55121 12202 55187 12205
rect 45461 12200 55187 12202
rect 45461 12144 45466 12200
rect 45522 12144 55126 12200
rect 55182 12144 55187 12200
rect 45461 12142 55187 12144
rect 45461 12139 45527 12142
rect 55121 12139 55187 12142
rect 77293 12202 77359 12205
rect 122833 12202 122899 12205
rect 77293 12200 122899 12202
rect 77293 12144 77298 12200
rect 77354 12144 122838 12200
rect 122894 12144 122899 12200
rect 77293 12142 122899 12144
rect 77293 12139 77359 12142
rect 122833 12139 122899 12142
rect 123845 12202 123911 12205
rect 125317 12202 125383 12205
rect 123845 12200 125383 12202
rect 123845 12144 123850 12200
rect 123906 12144 125322 12200
rect 125378 12144 125383 12200
rect 123845 12142 125383 12144
rect 123845 12139 123911 12142
rect 125317 12139 125383 12142
rect 127709 12202 127775 12205
rect 130653 12202 130719 12205
rect 127709 12200 130719 12202
rect 127709 12144 127714 12200
rect 127770 12144 130658 12200
rect 130714 12144 130719 12200
rect 127709 12142 130719 12144
rect 127709 12139 127775 12142
rect 130653 12139 130719 12142
rect 133965 12202 134031 12205
rect 147630 12202 147690 12278
rect 156321 12275 156387 12278
rect 133965 12200 147690 12202
rect 133965 12144 133970 12200
rect 134026 12144 147690 12200
rect 133965 12142 147690 12144
rect 133965 12139 134031 12142
rect 104341 12066 104407 12069
rect 105813 12066 105879 12069
rect 104341 12064 105879 12066
rect 104341 12008 104346 12064
rect 104402 12008 105818 12064
rect 105874 12008 105879 12064
rect 104341 12006 105879 12008
rect 104341 12003 104407 12006
rect 105813 12003 105879 12006
rect 116485 12066 116551 12069
rect 119061 12066 119127 12069
rect 116485 12064 119127 12066
rect 116485 12008 116490 12064
rect 116546 12008 119066 12064
rect 119122 12008 119127 12064
rect 116485 12006 119127 12008
rect 116485 12003 116551 12006
rect 119061 12003 119127 12006
rect 120809 12066 120875 12069
rect 127198 12066 127204 12068
rect 120809 12064 127204 12066
rect 120809 12008 120814 12064
rect 120870 12008 127204 12064
rect 120809 12006 127204 12008
rect 120809 12003 120875 12006
rect 127198 12004 127204 12006
rect 127268 12004 127274 12068
rect 130009 12066 130075 12069
rect 143073 12066 143139 12069
rect 153469 12066 153535 12069
rect 130009 12064 143139 12066
rect 130009 12008 130014 12064
rect 130070 12008 143078 12064
rect 143134 12008 143139 12064
rect 130009 12006 143139 12008
rect 130009 12003 130075 12006
rect 143073 12003 143139 12006
rect 143214 12064 153535 12066
rect 143214 12008 153474 12064
rect 153530 12008 153535 12064
rect 143214 12006 153535 12008
rect 40390 12000 40706 12001
rect 40390 11936 40396 12000
rect 40460 11936 40476 12000
rect 40540 11936 40556 12000
rect 40620 11936 40636 12000
rect 40700 11936 40706 12000
rect 40390 11935 40706 11936
rect 79835 12000 80151 12001
rect 79835 11936 79841 12000
rect 79905 11936 79921 12000
rect 79985 11936 80001 12000
rect 80065 11936 80081 12000
rect 80145 11936 80151 12000
rect 79835 11935 80151 11936
rect 119280 12000 119596 12001
rect 119280 11936 119286 12000
rect 119350 11936 119366 12000
rect 119430 11936 119446 12000
rect 119510 11936 119526 12000
rect 119590 11936 119596 12000
rect 119280 11935 119596 11936
rect 48773 11930 48839 11933
rect 52821 11930 52887 11933
rect 118877 11930 118943 11933
rect 48773 11928 52887 11930
rect 48773 11872 48778 11928
rect 48834 11872 52826 11928
rect 52882 11872 52887 11928
rect 48773 11870 52887 11872
rect 48773 11867 48839 11870
rect 52821 11867 52887 11870
rect 99330 11928 118943 11930
rect 99330 11872 118882 11928
rect 118938 11872 118943 11928
rect 99330 11870 118943 11872
rect 11881 11794 11947 11797
rect 15929 11794 15995 11797
rect 11881 11792 15995 11794
rect 11881 11736 11886 11792
rect 11942 11736 15934 11792
rect 15990 11736 15995 11792
rect 11881 11734 15995 11736
rect 11881 11731 11947 11734
rect 15929 11731 15995 11734
rect 61561 11794 61627 11797
rect 96797 11794 96863 11797
rect 61561 11792 96863 11794
rect 61561 11736 61566 11792
rect 61622 11736 96802 11792
rect 96858 11736 96863 11792
rect 61561 11734 96863 11736
rect 61561 11731 61627 11734
rect 96797 11731 96863 11734
rect 98453 11794 98519 11797
rect 99330 11794 99390 11870
rect 118877 11867 118943 11870
rect 120165 11930 120231 11933
rect 125501 11930 125567 11933
rect 120165 11928 125567 11930
rect 120165 11872 120170 11928
rect 120226 11872 125506 11928
rect 125562 11872 125567 11928
rect 120165 11870 125567 11872
rect 120165 11867 120231 11870
rect 125501 11867 125567 11870
rect 127341 11930 127407 11933
rect 131062 11930 131068 11932
rect 127341 11928 131068 11930
rect 127341 11872 127346 11928
rect 127402 11872 131068 11928
rect 127341 11870 131068 11872
rect 127341 11867 127407 11870
rect 131062 11868 131068 11870
rect 131132 11930 131138 11932
rect 131205 11930 131271 11933
rect 131132 11928 131271 11930
rect 131132 11872 131210 11928
rect 131266 11872 131271 11928
rect 131132 11870 131271 11872
rect 131132 11868 131138 11870
rect 131205 11867 131271 11870
rect 142613 11930 142679 11933
rect 143214 11930 143274 12006
rect 153469 12003 153535 12006
rect 158725 12000 159041 12001
rect 158725 11936 158731 12000
rect 158795 11936 158811 12000
rect 158875 11936 158891 12000
rect 158955 11936 158971 12000
rect 159035 11936 159041 12000
rect 158725 11935 159041 11936
rect 142613 11928 143274 11930
rect 142613 11872 142618 11928
rect 142674 11872 143274 11928
rect 142613 11870 143274 11872
rect 145005 11930 145071 11933
rect 147990 11930 147996 11932
rect 145005 11928 147996 11930
rect 145005 11872 145010 11928
rect 145066 11872 147996 11928
rect 145005 11870 147996 11872
rect 142613 11867 142679 11870
rect 145005 11867 145071 11870
rect 147990 11868 147996 11870
rect 148060 11868 148066 11932
rect 148501 11930 148567 11933
rect 150617 11930 150683 11933
rect 148501 11928 150683 11930
rect 148501 11872 148506 11928
rect 148562 11872 150622 11928
rect 150678 11872 150683 11928
rect 148501 11870 150683 11872
rect 148501 11867 148567 11870
rect 150617 11867 150683 11870
rect 98453 11792 99390 11794
rect 98453 11736 98458 11792
rect 98514 11736 99390 11792
rect 98453 11734 99390 11736
rect 117313 11794 117379 11797
rect 121637 11794 121703 11797
rect 117313 11792 121703 11794
rect 117313 11736 117318 11792
rect 117374 11736 121642 11792
rect 121698 11736 121703 11792
rect 117313 11734 121703 11736
rect 98453 11731 98519 11734
rect 117313 11731 117379 11734
rect 121637 11731 121703 11734
rect 124305 11794 124371 11797
rect 124949 11794 125015 11797
rect 124305 11792 125015 11794
rect 124305 11736 124310 11792
rect 124366 11736 124954 11792
rect 125010 11736 125015 11792
rect 124305 11734 125015 11736
rect 124305 11731 124371 11734
rect 124949 11731 125015 11734
rect 133454 11732 133460 11796
rect 133524 11794 133530 11796
rect 150433 11794 150499 11797
rect 133524 11792 150499 11794
rect 133524 11736 150438 11792
rect 150494 11736 150499 11792
rect 133524 11734 150499 11736
rect 133524 11732 133530 11734
rect 150433 11731 150499 11734
rect 155309 11794 155375 11797
rect 156137 11794 156203 11797
rect 155309 11792 156203 11794
rect 155309 11736 155314 11792
rect 155370 11736 156142 11792
rect 156198 11736 156203 11792
rect 155309 11734 156203 11736
rect 155309 11731 155375 11734
rect 156137 11731 156203 11734
rect 10685 11658 10751 11661
rect 12893 11658 12959 11661
rect 10685 11656 12959 11658
rect 10685 11600 10690 11656
rect 10746 11600 12898 11656
rect 12954 11600 12959 11656
rect 10685 11598 12959 11600
rect 10685 11595 10751 11598
rect 12893 11595 12959 11598
rect 20621 11658 20687 11661
rect 22461 11658 22527 11661
rect 20621 11656 22527 11658
rect 20621 11600 20626 11656
rect 20682 11600 22466 11656
rect 22522 11600 22527 11656
rect 20621 11598 22527 11600
rect 20621 11595 20687 11598
rect 22461 11595 22527 11598
rect 34789 11658 34855 11661
rect 53925 11658 53991 11661
rect 34789 11656 53991 11658
rect 34789 11600 34794 11656
rect 34850 11600 53930 11656
rect 53986 11600 53991 11656
rect 34789 11598 53991 11600
rect 34789 11595 34855 11598
rect 53925 11595 53991 11598
rect 78765 11658 78831 11661
rect 86677 11658 86743 11661
rect 78765 11656 86743 11658
rect 78765 11600 78770 11656
rect 78826 11600 86682 11656
rect 86738 11600 86743 11656
rect 78765 11598 86743 11600
rect 78765 11595 78831 11598
rect 86677 11595 86743 11598
rect 99373 11658 99439 11661
rect 143165 11658 143231 11661
rect 99373 11656 143231 11658
rect 99373 11600 99378 11656
rect 99434 11600 143170 11656
rect 143226 11600 143231 11656
rect 99373 11598 143231 11600
rect 99373 11595 99439 11598
rect 143165 11595 143231 11598
rect 145833 11658 145899 11661
rect 149237 11658 149303 11661
rect 145833 11656 149303 11658
rect 145833 11600 145838 11656
rect 145894 11600 149242 11656
rect 149298 11600 149303 11656
rect 145833 11598 149303 11600
rect 145833 11595 145899 11598
rect 149237 11595 149303 11598
rect 149421 11658 149487 11661
rect 151445 11658 151511 11661
rect 149421 11656 151511 11658
rect 149421 11600 149426 11656
rect 149482 11600 151450 11656
rect 151506 11600 151511 11656
rect 149421 11598 151511 11600
rect 149421 11595 149487 11598
rect 151445 11595 151511 11598
rect 42609 11522 42675 11525
rect 43069 11522 43135 11525
rect 42609 11520 43135 11522
rect 42609 11464 42614 11520
rect 42670 11464 43074 11520
rect 43130 11464 43135 11520
rect 42609 11462 43135 11464
rect 42609 11459 42675 11462
rect 43069 11459 43135 11462
rect 50705 11522 50771 11525
rect 52545 11522 52611 11525
rect 50705 11520 52611 11522
rect 50705 11464 50710 11520
rect 50766 11464 52550 11520
rect 52606 11464 52611 11520
rect 50705 11462 52611 11464
rect 50705 11459 50771 11462
rect 52545 11459 52611 11462
rect 88149 11522 88215 11525
rect 90357 11522 90423 11525
rect 88149 11520 90423 11522
rect 88149 11464 88154 11520
rect 88210 11464 90362 11520
rect 90418 11464 90423 11520
rect 88149 11462 90423 11464
rect 88149 11459 88215 11462
rect 90357 11459 90423 11462
rect 123937 11522 124003 11525
rect 133045 11522 133111 11525
rect 123937 11520 133111 11522
rect 123937 11464 123942 11520
rect 123998 11464 133050 11520
rect 133106 11464 133111 11520
rect 123937 11462 133111 11464
rect 123937 11459 124003 11462
rect 133045 11459 133111 11462
rect 143257 11522 143323 11525
rect 152641 11522 152707 11525
rect 143257 11520 152707 11522
rect 143257 11464 143262 11520
rect 143318 11464 152646 11520
rect 152702 11464 152707 11520
rect 143257 11462 152707 11464
rect 143257 11459 143323 11462
rect 152641 11459 152707 11462
rect 20668 11456 20984 11457
rect 20668 11392 20674 11456
rect 20738 11392 20754 11456
rect 20818 11392 20834 11456
rect 20898 11392 20914 11456
rect 20978 11392 20984 11456
rect 20668 11391 20984 11392
rect 60113 11456 60429 11457
rect 60113 11392 60119 11456
rect 60183 11392 60199 11456
rect 60263 11392 60279 11456
rect 60343 11392 60359 11456
rect 60423 11392 60429 11456
rect 60113 11391 60429 11392
rect 99558 11456 99874 11457
rect 99558 11392 99564 11456
rect 99628 11392 99644 11456
rect 99708 11392 99724 11456
rect 99788 11392 99804 11456
rect 99868 11392 99874 11456
rect 99558 11391 99874 11392
rect 139003 11456 139319 11457
rect 139003 11392 139009 11456
rect 139073 11392 139089 11456
rect 139153 11392 139169 11456
rect 139233 11392 139249 11456
rect 139313 11392 139319 11456
rect 139003 11391 139319 11392
rect 42057 11386 42123 11389
rect 45369 11386 45435 11389
rect 42057 11384 45435 11386
rect 42057 11328 42062 11384
rect 42118 11328 45374 11384
rect 45430 11328 45435 11384
rect 42057 11326 45435 11328
rect 42057 11323 42123 11326
rect 45369 11323 45435 11326
rect 86217 11386 86283 11389
rect 93669 11386 93735 11389
rect 86217 11384 93735 11386
rect 86217 11328 86222 11384
rect 86278 11328 93674 11384
rect 93730 11328 93735 11384
rect 86217 11326 93735 11328
rect 86217 11323 86283 11326
rect 93669 11323 93735 11326
rect 121361 11386 121427 11389
rect 124213 11386 124279 11389
rect 121361 11384 124279 11386
rect 121361 11328 121366 11384
rect 121422 11328 124218 11384
rect 124274 11328 124279 11384
rect 121361 11326 124279 11328
rect 121361 11323 121427 11326
rect 124213 11323 124279 11326
rect 124949 11386 125015 11389
rect 139485 11386 139551 11389
rect 141325 11386 141391 11389
rect 124949 11384 128370 11386
rect 124949 11328 124954 11384
rect 125010 11328 128370 11384
rect 124949 11326 128370 11328
rect 124949 11323 125015 11326
rect 10501 11250 10567 11253
rect 14089 11250 14155 11253
rect 10501 11248 14155 11250
rect 10501 11192 10506 11248
rect 10562 11192 14094 11248
rect 14150 11192 14155 11248
rect 10501 11190 14155 11192
rect 10501 11187 10567 11190
rect 14089 11187 14155 11190
rect 51625 11250 51691 11253
rect 58617 11250 58683 11253
rect 51625 11248 58683 11250
rect 51625 11192 51630 11248
rect 51686 11192 58622 11248
rect 58678 11192 58683 11248
rect 51625 11190 58683 11192
rect 51625 11187 51691 11190
rect 58617 11187 58683 11190
rect 92841 11250 92907 11253
rect 121177 11250 121243 11253
rect 123661 11250 123727 11253
rect 92841 11248 123727 11250
rect 92841 11192 92846 11248
rect 92902 11192 121182 11248
rect 121238 11192 123666 11248
rect 123722 11192 123727 11248
rect 92841 11190 123727 11192
rect 92841 11187 92907 11190
rect 121177 11187 121243 11190
rect 123661 11187 123727 11190
rect 124305 11250 124371 11253
rect 127893 11250 127959 11253
rect 124305 11248 127959 11250
rect 124305 11192 124310 11248
rect 124366 11192 127898 11248
rect 127954 11192 127959 11248
rect 124305 11190 127959 11192
rect 128310 11250 128370 11326
rect 139485 11384 141391 11386
rect 139485 11328 139490 11384
rect 139546 11328 141330 11384
rect 141386 11328 141391 11384
rect 139485 11326 141391 11328
rect 139485 11323 139551 11326
rect 141325 11323 141391 11326
rect 145281 11386 145347 11389
rect 147673 11386 147739 11389
rect 145281 11384 147739 11386
rect 145281 11328 145286 11384
rect 145342 11328 147678 11384
rect 147734 11328 147739 11384
rect 145281 11326 147739 11328
rect 145281 11323 145347 11326
rect 147673 11323 147739 11326
rect 148041 11386 148107 11389
rect 154665 11386 154731 11389
rect 148041 11384 154731 11386
rect 148041 11328 148046 11384
rect 148102 11328 154670 11384
rect 154726 11328 154731 11384
rect 148041 11326 154731 11328
rect 148041 11323 148107 11326
rect 154665 11323 154731 11326
rect 141509 11250 141575 11253
rect 128310 11248 141575 11250
rect 128310 11192 141514 11248
rect 141570 11192 141575 11248
rect 128310 11190 141575 11192
rect 124305 11187 124371 11190
rect 127893 11187 127959 11190
rect 141509 11187 141575 11190
rect 144637 11250 144703 11253
rect 157057 11250 157123 11253
rect 144637 11248 157123 11250
rect 144637 11192 144642 11248
rect 144698 11192 157062 11248
rect 157118 11192 157123 11248
rect 144637 11190 157123 11192
rect 144637 11187 144703 11190
rect 157057 11187 157123 11190
rect 19333 11114 19399 11117
rect 28901 11114 28967 11117
rect 19333 11112 28967 11114
rect 19333 11056 19338 11112
rect 19394 11056 28906 11112
rect 28962 11056 28967 11112
rect 19333 11054 28967 11056
rect 19333 11051 19399 11054
rect 28901 11051 28967 11054
rect 72969 11114 73035 11117
rect 100661 11114 100727 11117
rect 72969 11112 100727 11114
rect 72969 11056 72974 11112
rect 73030 11056 100666 11112
rect 100722 11056 100727 11112
rect 72969 11054 100727 11056
rect 72969 11051 73035 11054
rect 100661 11051 100727 11054
rect 116945 11114 117011 11117
rect 128077 11114 128143 11117
rect 116945 11112 128143 11114
rect 116945 11056 116950 11112
rect 117006 11056 128082 11112
rect 128138 11056 128143 11112
rect 116945 11054 128143 11056
rect 116945 11051 117011 11054
rect 128077 11051 128143 11054
rect 130653 11114 130719 11117
rect 140405 11114 140471 11117
rect 130653 11112 140471 11114
rect 130653 11056 130658 11112
rect 130714 11056 140410 11112
rect 140466 11056 140471 11112
rect 130653 11054 140471 11056
rect 130653 11051 130719 11054
rect 140405 11051 140471 11054
rect 143441 11114 143507 11117
rect 147438 11114 147444 11116
rect 143441 11112 147444 11114
rect 143441 11056 143446 11112
rect 143502 11056 147444 11112
rect 143441 11054 147444 11056
rect 143441 11051 143507 11054
rect 147438 11052 147444 11054
rect 147508 11052 147514 11116
rect 147765 11114 147831 11117
rect 152365 11114 152431 11117
rect 152825 11116 152891 11117
rect 152774 11114 152780 11116
rect 147765 11112 152431 11114
rect 147765 11056 147770 11112
rect 147826 11056 152370 11112
rect 152426 11056 152431 11112
rect 147765 11054 152431 11056
rect 152734 11054 152780 11114
rect 152844 11112 152891 11116
rect 152886 11056 152891 11112
rect 147765 11051 147831 11054
rect 152365 11051 152431 11054
rect 152774 11052 152780 11054
rect 152844 11052 152891 11056
rect 152825 11051 152891 11052
rect 26877 10978 26943 10981
rect 30373 10978 30439 10981
rect 26877 10976 30439 10978
rect 26877 10920 26882 10976
rect 26938 10920 30378 10976
rect 30434 10920 30439 10976
rect 26877 10918 30439 10920
rect 26877 10915 26943 10918
rect 30373 10915 30439 10918
rect 49141 10978 49207 10981
rect 51165 10978 51231 10981
rect 49141 10976 51231 10978
rect 49141 10920 49146 10976
rect 49202 10920 51170 10976
rect 51226 10920 51231 10976
rect 49141 10918 51231 10920
rect 49141 10915 49207 10918
rect 51165 10915 51231 10918
rect 67725 10978 67791 10981
rect 74625 10978 74691 10981
rect 67725 10976 74691 10978
rect 67725 10920 67730 10976
rect 67786 10920 74630 10976
rect 74686 10920 74691 10976
rect 67725 10918 74691 10920
rect 67725 10915 67791 10918
rect 74625 10915 74691 10918
rect 81249 10978 81315 10981
rect 86861 10978 86927 10981
rect 81249 10976 86927 10978
rect 81249 10920 81254 10976
rect 81310 10920 86866 10976
rect 86922 10920 86927 10976
rect 81249 10918 86927 10920
rect 81249 10915 81315 10918
rect 86861 10915 86927 10918
rect 124765 10978 124831 10981
rect 128629 10978 128695 10981
rect 124765 10976 128695 10978
rect 124765 10920 124770 10976
rect 124826 10920 128634 10976
rect 128690 10920 128695 10976
rect 124765 10918 128695 10920
rect 124765 10915 124831 10918
rect 128629 10915 128695 10918
rect 135161 10978 135227 10981
rect 141233 10978 141299 10981
rect 135161 10976 141299 10978
rect 135161 10920 135166 10976
rect 135222 10920 141238 10976
rect 141294 10920 141299 10976
rect 135161 10918 141299 10920
rect 135161 10915 135227 10918
rect 141233 10915 141299 10918
rect 146334 10916 146340 10980
rect 146404 10978 146410 10980
rect 156965 10978 157031 10981
rect 146404 10976 157031 10978
rect 146404 10920 156970 10976
rect 157026 10920 157031 10976
rect 146404 10918 157031 10920
rect 146404 10916 146410 10918
rect 156965 10915 157031 10918
rect 40390 10912 40706 10913
rect 40390 10848 40396 10912
rect 40460 10848 40476 10912
rect 40540 10848 40556 10912
rect 40620 10848 40636 10912
rect 40700 10848 40706 10912
rect 40390 10847 40706 10848
rect 79835 10912 80151 10913
rect 79835 10848 79841 10912
rect 79905 10848 79921 10912
rect 79985 10848 80001 10912
rect 80065 10848 80081 10912
rect 80145 10848 80151 10912
rect 79835 10847 80151 10848
rect 119280 10912 119596 10913
rect 119280 10848 119286 10912
rect 119350 10848 119366 10912
rect 119430 10848 119446 10912
rect 119510 10848 119526 10912
rect 119590 10848 119596 10912
rect 119280 10847 119596 10848
rect 158725 10912 159041 10913
rect 158725 10848 158731 10912
rect 158795 10848 158811 10912
rect 158875 10848 158891 10912
rect 158955 10848 158971 10912
rect 159035 10848 159041 10912
rect 158725 10847 159041 10848
rect 50153 10842 50219 10845
rect 53833 10842 53899 10845
rect 50153 10840 53899 10842
rect 50153 10784 50158 10840
rect 50214 10784 53838 10840
rect 53894 10784 53899 10840
rect 50153 10782 53899 10784
rect 50153 10779 50219 10782
rect 53833 10779 53899 10782
rect 58341 10842 58407 10845
rect 63861 10842 63927 10845
rect 107837 10842 107903 10845
rect 109033 10842 109099 10845
rect 58341 10840 63927 10842
rect 58341 10784 58346 10840
rect 58402 10784 63866 10840
rect 63922 10784 63927 10840
rect 58341 10782 63927 10784
rect 58341 10779 58407 10782
rect 63861 10779 63927 10782
rect 89670 10840 107903 10842
rect 89670 10784 107842 10840
rect 107898 10784 107903 10840
rect 89670 10782 107903 10784
rect 17217 10706 17283 10709
rect 27797 10706 27863 10709
rect 17217 10704 27863 10706
rect 17217 10648 17222 10704
rect 17278 10648 27802 10704
rect 27858 10648 27863 10704
rect 17217 10646 27863 10648
rect 17217 10643 17283 10646
rect 27797 10643 27863 10646
rect 52545 10706 52611 10709
rect 53097 10706 53163 10709
rect 63861 10706 63927 10709
rect 52545 10704 63927 10706
rect 52545 10648 52550 10704
rect 52606 10648 53102 10704
rect 53158 10648 63866 10704
rect 63922 10648 63927 10704
rect 52545 10646 63927 10648
rect 52545 10643 52611 10646
rect 53097 10643 53163 10646
rect 63861 10643 63927 10646
rect 79869 10706 79935 10709
rect 89670 10706 89730 10782
rect 107837 10779 107903 10782
rect 108990 10840 109099 10842
rect 108990 10784 109038 10840
rect 109094 10784 109099 10840
rect 108990 10779 109099 10784
rect 116025 10842 116091 10845
rect 118969 10842 119035 10845
rect 116025 10840 119035 10842
rect 116025 10784 116030 10840
rect 116086 10784 118974 10840
rect 119030 10784 119035 10840
rect 116025 10782 119035 10784
rect 116025 10779 116091 10782
rect 118969 10779 119035 10782
rect 125685 10842 125751 10845
rect 126145 10842 126211 10845
rect 125685 10840 126211 10842
rect 125685 10784 125690 10840
rect 125746 10784 126150 10840
rect 126206 10784 126211 10840
rect 125685 10782 126211 10784
rect 125685 10779 125751 10782
rect 126145 10779 126211 10782
rect 138013 10842 138079 10845
rect 138749 10842 138815 10845
rect 138013 10840 138815 10842
rect 138013 10784 138018 10840
rect 138074 10784 138754 10840
rect 138810 10784 138815 10840
rect 138013 10782 138815 10784
rect 138013 10779 138079 10782
rect 138749 10779 138815 10782
rect 144729 10842 144795 10845
rect 148317 10842 148383 10845
rect 144729 10840 148383 10842
rect 144729 10784 144734 10840
rect 144790 10784 148322 10840
rect 148378 10784 148383 10840
rect 144729 10782 148383 10784
rect 144729 10779 144795 10782
rect 148317 10779 148383 10782
rect 148777 10842 148843 10845
rect 155217 10842 155283 10845
rect 148777 10840 155283 10842
rect 148777 10784 148782 10840
rect 148838 10784 155222 10840
rect 155278 10784 155283 10840
rect 148777 10782 155283 10784
rect 148777 10779 148843 10782
rect 155217 10779 155283 10782
rect 79869 10704 89730 10706
rect 79869 10648 79874 10704
rect 79930 10648 89730 10704
rect 79869 10646 89730 10648
rect 107745 10706 107811 10709
rect 108990 10706 109050 10779
rect 107745 10704 109050 10706
rect 107745 10648 107750 10704
rect 107806 10648 109050 10704
rect 107745 10646 109050 10648
rect 113449 10706 113515 10709
rect 118509 10706 118575 10709
rect 113449 10704 118575 10706
rect 113449 10648 113454 10704
rect 113510 10648 118514 10704
rect 118570 10648 118575 10704
rect 113449 10646 118575 10648
rect 79869 10643 79935 10646
rect 107745 10643 107811 10646
rect 113449 10643 113515 10646
rect 118509 10643 118575 10646
rect 123201 10706 123267 10709
rect 152641 10706 152707 10709
rect 123201 10704 152707 10706
rect 123201 10648 123206 10704
rect 123262 10648 152646 10704
rect 152702 10648 152707 10704
rect 123201 10646 152707 10648
rect 123201 10643 123267 10646
rect 152641 10643 152707 10646
rect 12433 10570 12499 10573
rect 13353 10570 13419 10573
rect 34421 10570 34487 10573
rect 12433 10568 34487 10570
rect 12433 10512 12438 10568
rect 12494 10512 13358 10568
rect 13414 10512 34426 10568
rect 34482 10512 34487 10568
rect 12433 10510 34487 10512
rect 12433 10507 12499 10510
rect 13353 10507 13419 10510
rect 34421 10507 34487 10510
rect 87229 10570 87295 10573
rect 127065 10570 127131 10573
rect 87229 10568 127131 10570
rect 87229 10512 87234 10568
rect 87290 10512 127070 10568
rect 127126 10512 127131 10568
rect 87229 10510 127131 10512
rect 87229 10507 87295 10510
rect 127065 10507 127131 10510
rect 127985 10570 128051 10573
rect 135529 10570 135595 10573
rect 127985 10568 135595 10570
rect 127985 10512 127990 10568
rect 128046 10512 135534 10568
rect 135590 10512 135595 10568
rect 127985 10510 135595 10512
rect 127985 10507 128051 10510
rect 135529 10507 135595 10510
rect 136633 10570 136699 10573
rect 156137 10570 156203 10573
rect 136633 10568 156203 10570
rect 136633 10512 136638 10568
rect 136694 10512 156142 10568
rect 156198 10512 156203 10568
rect 136633 10510 156203 10512
rect 136633 10507 136699 10510
rect 156137 10507 156203 10510
rect 48773 10434 48839 10437
rect 56501 10434 56567 10437
rect 48773 10432 56567 10434
rect 48773 10376 48778 10432
rect 48834 10376 56506 10432
rect 56562 10376 56567 10432
rect 48773 10374 56567 10376
rect 48773 10371 48839 10374
rect 56501 10371 56567 10374
rect 104157 10434 104223 10437
rect 120349 10434 120415 10437
rect 104157 10432 120415 10434
rect 104157 10376 104162 10432
rect 104218 10376 120354 10432
rect 120410 10376 120415 10432
rect 104157 10374 120415 10376
rect 104157 10371 104223 10374
rect 120349 10371 120415 10374
rect 121729 10434 121795 10437
rect 134517 10434 134583 10437
rect 121729 10432 134583 10434
rect 121729 10376 121734 10432
rect 121790 10376 134522 10432
rect 134578 10376 134583 10432
rect 121729 10374 134583 10376
rect 121729 10371 121795 10374
rect 134517 10371 134583 10374
rect 139761 10434 139827 10437
rect 151721 10434 151787 10437
rect 139761 10432 151787 10434
rect 139761 10376 139766 10432
rect 139822 10376 151726 10432
rect 151782 10376 151787 10432
rect 139761 10374 151787 10376
rect 139761 10371 139827 10374
rect 151721 10371 151787 10374
rect 20668 10368 20984 10369
rect 20668 10304 20674 10368
rect 20738 10304 20754 10368
rect 20818 10304 20834 10368
rect 20898 10304 20914 10368
rect 20978 10304 20984 10368
rect 20668 10303 20984 10304
rect 60113 10368 60429 10369
rect 60113 10304 60119 10368
rect 60183 10304 60199 10368
rect 60263 10304 60279 10368
rect 60343 10304 60359 10368
rect 60423 10304 60429 10368
rect 60113 10303 60429 10304
rect 99558 10368 99874 10369
rect 99558 10304 99564 10368
rect 99628 10304 99644 10368
rect 99708 10304 99724 10368
rect 99788 10304 99804 10368
rect 99868 10304 99874 10368
rect 99558 10303 99874 10304
rect 139003 10368 139319 10369
rect 139003 10304 139009 10368
rect 139073 10304 139089 10368
rect 139153 10304 139169 10368
rect 139233 10304 139249 10368
rect 139313 10304 139319 10368
rect 139003 10303 139319 10304
rect 49141 10298 49207 10301
rect 57513 10298 57579 10301
rect 49141 10296 57579 10298
rect 49141 10240 49146 10296
rect 49202 10240 57518 10296
rect 57574 10240 57579 10296
rect 49141 10238 57579 10240
rect 49141 10235 49207 10238
rect 57513 10235 57579 10238
rect 93209 10298 93275 10301
rect 95509 10298 95575 10301
rect 93209 10296 95575 10298
rect 93209 10240 93214 10296
rect 93270 10240 95514 10296
rect 95570 10240 95575 10296
rect 93209 10238 95575 10240
rect 93209 10235 93275 10238
rect 95509 10235 95575 10238
rect 101857 10298 101923 10301
rect 104985 10298 105051 10301
rect 101857 10296 105051 10298
rect 101857 10240 101862 10296
rect 101918 10240 104990 10296
rect 105046 10240 105051 10296
rect 101857 10238 105051 10240
rect 101857 10235 101923 10238
rect 104985 10235 105051 10238
rect 105169 10298 105235 10301
rect 129641 10298 129707 10301
rect 105169 10296 129707 10298
rect 105169 10240 105174 10296
rect 105230 10240 129646 10296
rect 129702 10240 129707 10296
rect 105169 10238 129707 10240
rect 105169 10235 105235 10238
rect 129641 10235 129707 10238
rect 131757 10298 131823 10301
rect 137185 10298 137251 10301
rect 131757 10296 137251 10298
rect 131757 10240 131762 10296
rect 131818 10240 137190 10296
rect 137246 10240 137251 10296
rect 131757 10238 137251 10240
rect 131757 10235 131823 10238
rect 137185 10235 137251 10238
rect 139853 10298 139919 10301
rect 149421 10298 149487 10301
rect 150249 10298 150315 10301
rect 139853 10296 150315 10298
rect 139853 10240 139858 10296
rect 139914 10240 149426 10296
rect 149482 10240 150254 10296
rect 150310 10240 150315 10296
rect 139853 10238 150315 10240
rect 139853 10235 139919 10238
rect 149421 10235 149487 10238
rect 150249 10235 150315 10238
rect 150382 10236 150388 10300
rect 150452 10298 150458 10300
rect 154665 10298 154731 10301
rect 159265 10298 159331 10301
rect 150452 10296 159331 10298
rect 150452 10240 154670 10296
rect 154726 10240 159270 10296
rect 159326 10240 159331 10296
rect 150452 10238 159331 10240
rect 150452 10236 150458 10238
rect 154665 10235 154731 10238
rect 159265 10235 159331 10238
rect 51533 10162 51599 10165
rect 52177 10162 52243 10165
rect 54385 10162 54451 10165
rect 55949 10162 56015 10165
rect 58985 10162 59051 10165
rect 51533 10160 59051 10162
rect 51533 10104 51538 10160
rect 51594 10104 52182 10160
rect 52238 10104 54390 10160
rect 54446 10104 55954 10160
rect 56010 10104 58990 10160
rect 59046 10104 59051 10160
rect 51533 10102 59051 10104
rect 51533 10099 51599 10102
rect 52177 10099 52243 10102
rect 54385 10099 54451 10102
rect 55949 10099 56015 10102
rect 58985 10099 59051 10102
rect 59997 10162 60063 10165
rect 60825 10162 60891 10165
rect 59997 10160 60891 10162
rect 59997 10104 60002 10160
rect 60058 10104 60830 10160
rect 60886 10104 60891 10160
rect 59997 10102 60891 10104
rect 59997 10099 60063 10102
rect 60825 10099 60891 10102
rect 70485 10162 70551 10165
rect 71221 10162 71287 10165
rect 104709 10162 104775 10165
rect 70485 10160 104775 10162
rect 70485 10104 70490 10160
rect 70546 10104 71226 10160
rect 71282 10104 104714 10160
rect 104770 10104 104775 10160
rect 70485 10102 104775 10104
rect 70485 10099 70551 10102
rect 71221 10099 71287 10102
rect 104709 10099 104775 10102
rect 107745 10162 107811 10165
rect 111609 10162 111675 10165
rect 107745 10160 111675 10162
rect 107745 10104 107750 10160
rect 107806 10104 111614 10160
rect 111670 10104 111675 10160
rect 107745 10102 111675 10104
rect 107745 10099 107811 10102
rect 111609 10099 111675 10102
rect 113541 10162 113607 10165
rect 153837 10162 153903 10165
rect 113541 10160 153903 10162
rect 113541 10104 113546 10160
rect 113602 10104 153842 10160
rect 153898 10104 153903 10160
rect 113541 10102 153903 10104
rect 113541 10099 113607 10102
rect 153837 10099 153903 10102
rect 54201 10026 54267 10029
rect 57053 10026 57119 10029
rect 67633 10026 67699 10029
rect 54201 10024 57119 10026
rect 54201 9968 54206 10024
rect 54262 9968 57058 10024
rect 57114 9968 57119 10024
rect 54201 9966 57119 9968
rect 54201 9963 54267 9966
rect 57053 9963 57119 9966
rect 67590 10024 67699 10026
rect 67590 9968 67638 10024
rect 67694 9968 67699 10024
rect 67590 9963 67699 9968
rect 74717 10026 74783 10029
rect 118233 10026 118299 10029
rect 120717 10026 120783 10029
rect 122925 10026 122991 10029
rect 74717 10024 118299 10026
rect 74717 9968 74722 10024
rect 74778 9968 118238 10024
rect 118294 9968 118299 10024
rect 74717 9966 118299 9968
rect 74717 9963 74783 9966
rect 118233 9963 118299 9966
rect 118650 9966 119722 10026
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 54109 9890 54175 9893
rect 57789 9890 57855 9893
rect 54109 9888 57855 9890
rect 54109 9832 54114 9888
rect 54170 9832 57794 9888
rect 57850 9832 57855 9888
rect 54109 9830 57855 9832
rect 54109 9827 54175 9830
rect 57789 9827 57855 9830
rect 40390 9824 40706 9825
rect 40390 9760 40396 9824
rect 40460 9760 40476 9824
rect 40540 9760 40556 9824
rect 40620 9760 40636 9824
rect 40700 9760 40706 9824
rect 40390 9759 40706 9760
rect 67590 9757 67650 9963
rect 81249 9890 81315 9893
rect 84837 9890 84903 9893
rect 81249 9888 84903 9890
rect 81249 9832 81254 9888
rect 81310 9832 84842 9888
rect 84898 9832 84903 9888
rect 81249 9830 84903 9832
rect 81249 9827 81315 9830
rect 84837 9827 84903 9830
rect 95325 9890 95391 9893
rect 104157 9890 104223 9893
rect 95325 9888 104223 9890
rect 95325 9832 95330 9888
rect 95386 9832 104162 9888
rect 104218 9832 104223 9888
rect 95325 9830 104223 9832
rect 95325 9827 95391 9830
rect 104157 9827 104223 9830
rect 113081 9890 113147 9893
rect 118650 9890 118710 9966
rect 113081 9888 118710 9890
rect 113081 9832 113086 9888
rect 113142 9832 118710 9888
rect 113081 9830 118710 9832
rect 119662 9890 119722 9966
rect 120717 10024 122991 10026
rect 120717 9968 120722 10024
rect 120778 9968 122930 10024
rect 122986 9968 122991 10024
rect 120717 9966 122991 9968
rect 120717 9963 120783 9966
rect 122925 9963 122991 9966
rect 125593 10026 125659 10029
rect 126145 10026 126211 10029
rect 125593 10024 126211 10026
rect 125593 9968 125598 10024
rect 125654 9968 126150 10024
rect 126206 9968 126211 10024
rect 125593 9966 126211 9968
rect 125593 9963 125659 9966
rect 126145 9963 126211 9966
rect 126329 10026 126395 10029
rect 150065 10026 150131 10029
rect 126329 10024 150131 10026
rect 126329 9968 126334 10024
rect 126390 9968 150070 10024
rect 150126 9968 150131 10024
rect 126329 9966 150131 9968
rect 126329 9963 126395 9966
rect 150065 9963 150131 9966
rect 150433 10026 150499 10029
rect 151261 10026 151327 10029
rect 150433 10024 151327 10026
rect 150433 9968 150438 10024
rect 150494 9968 151266 10024
rect 151322 9968 151327 10024
rect 150433 9966 151327 9968
rect 150433 9963 150499 9966
rect 151261 9963 151327 9966
rect 154665 10026 154731 10029
rect 157517 10026 157583 10029
rect 154665 10024 157583 10026
rect 154665 9968 154670 10024
rect 154726 9968 157522 10024
rect 157578 9968 157583 10024
rect 154665 9966 157583 9968
rect 154665 9963 154731 9966
rect 157517 9963 157583 9966
rect 142797 9890 142863 9893
rect 119662 9888 142863 9890
rect 119662 9832 142802 9888
rect 142858 9832 142863 9888
rect 119662 9830 142863 9832
rect 113081 9827 113147 9830
rect 142797 9827 142863 9830
rect 148593 9890 148659 9893
rect 152181 9890 152247 9893
rect 148593 9888 152247 9890
rect 148593 9832 148598 9888
rect 148654 9832 152186 9888
rect 152242 9832 152247 9888
rect 148593 9830 152247 9832
rect 148593 9827 148659 9830
rect 152181 9827 152247 9830
rect 79835 9824 80151 9825
rect 79835 9760 79841 9824
rect 79905 9760 79921 9824
rect 79985 9760 80001 9824
rect 80065 9760 80081 9824
rect 80145 9760 80151 9824
rect 79835 9759 80151 9760
rect 119280 9824 119596 9825
rect 119280 9760 119286 9824
rect 119350 9760 119366 9824
rect 119430 9760 119446 9824
rect 119510 9760 119526 9824
rect 119590 9760 119596 9824
rect 119280 9759 119596 9760
rect 158725 9824 159041 9825
rect 158725 9760 158731 9824
rect 158795 9760 158811 9824
rect 158875 9760 158891 9824
rect 158955 9760 158971 9824
rect 159035 9760 159041 9824
rect 158725 9759 159041 9760
rect 32029 9754 32095 9757
rect 37181 9754 37247 9757
rect 32029 9752 37247 9754
rect 32029 9696 32034 9752
rect 32090 9696 37186 9752
rect 37242 9696 37247 9752
rect 32029 9694 37247 9696
rect 32029 9691 32095 9694
rect 37181 9691 37247 9694
rect 60457 9754 60523 9757
rect 62573 9754 62639 9757
rect 60457 9752 62639 9754
rect 60457 9696 60462 9752
rect 60518 9696 62578 9752
rect 62634 9696 62639 9752
rect 60457 9694 62639 9696
rect 67590 9752 67699 9757
rect 67590 9696 67638 9752
rect 67694 9696 67699 9752
rect 67590 9694 67699 9696
rect 60457 9691 60523 9694
rect 62573 9691 62639 9694
rect 67633 9691 67699 9694
rect 88241 9754 88307 9757
rect 90081 9754 90147 9757
rect 88241 9752 90147 9754
rect 88241 9696 88246 9752
rect 88302 9696 90086 9752
rect 90142 9696 90147 9752
rect 88241 9694 90147 9696
rect 88241 9691 88307 9694
rect 90081 9691 90147 9694
rect 107837 9754 107903 9757
rect 115841 9754 115907 9757
rect 107837 9752 115907 9754
rect 107837 9696 107842 9752
rect 107898 9696 115846 9752
rect 115902 9696 115907 9752
rect 107837 9694 115907 9696
rect 107837 9691 107903 9694
rect 115841 9691 115907 9694
rect 116945 9754 117011 9757
rect 119153 9754 119219 9757
rect 124397 9756 124463 9757
rect 124397 9754 124444 9756
rect 116945 9752 119219 9754
rect 116945 9696 116950 9752
rect 117006 9696 119158 9752
rect 119214 9696 119219 9752
rect 116945 9694 119219 9696
rect 124352 9752 124444 9754
rect 124352 9696 124402 9752
rect 124352 9694 124444 9696
rect 116945 9691 117011 9694
rect 119153 9691 119219 9694
rect 124397 9692 124444 9694
rect 124508 9692 124514 9756
rect 126145 9754 126211 9757
rect 133873 9754 133939 9757
rect 126145 9752 133939 9754
rect 126145 9696 126150 9752
rect 126206 9696 133878 9752
rect 133934 9696 133939 9752
rect 126145 9694 133939 9696
rect 124397 9691 124463 9692
rect 126145 9691 126211 9694
rect 133873 9691 133939 9694
rect 135621 9754 135687 9757
rect 139761 9754 139827 9757
rect 135621 9752 139827 9754
rect 135621 9696 135626 9752
rect 135682 9696 139766 9752
rect 139822 9696 139827 9752
rect 135621 9694 139827 9696
rect 135621 9691 135687 9694
rect 139761 9691 139827 9694
rect 143993 9754 144059 9757
rect 144637 9754 144703 9757
rect 143993 9752 144703 9754
rect 143993 9696 143998 9752
rect 144054 9696 144642 9752
rect 144698 9696 144703 9752
rect 143993 9694 144703 9696
rect 143993 9691 144059 9694
rect 144637 9691 144703 9694
rect 144913 9754 144979 9757
rect 157609 9754 157675 9757
rect 144913 9752 157675 9754
rect 144913 9696 144918 9752
rect 144974 9696 157614 9752
rect 157670 9696 157675 9752
rect 144913 9694 157675 9696
rect 144913 9691 144979 9694
rect 157609 9691 157675 9694
rect 56225 9618 56291 9621
rect 57145 9618 57211 9621
rect 56225 9616 57211 9618
rect 56225 9560 56230 9616
rect 56286 9560 57150 9616
rect 57206 9560 57211 9616
rect 56225 9558 57211 9560
rect 56225 9555 56291 9558
rect 57145 9555 57211 9558
rect 77845 9618 77911 9621
rect 112621 9618 112687 9621
rect 77845 9616 112687 9618
rect 77845 9560 77850 9616
rect 77906 9560 112626 9616
rect 112682 9560 112687 9616
rect 77845 9558 112687 9560
rect 77845 9555 77911 9558
rect 112621 9555 112687 9558
rect 114921 9618 114987 9621
rect 138565 9618 138631 9621
rect 139301 9618 139367 9621
rect 114921 9616 139367 9618
rect 114921 9560 114926 9616
rect 114982 9560 138570 9616
rect 138626 9560 139306 9616
rect 139362 9560 139367 9616
rect 114921 9558 139367 9560
rect 114921 9555 114987 9558
rect 138565 9555 138631 9558
rect 139301 9555 139367 9558
rect 140037 9618 140103 9621
rect 145557 9618 145623 9621
rect 151997 9618 152063 9621
rect 152549 9620 152615 9621
rect 152549 9618 152596 9620
rect 140037 9616 152063 9618
rect 140037 9560 140042 9616
rect 140098 9560 145562 9616
rect 145618 9560 152002 9616
rect 152058 9560 152063 9616
rect 140037 9558 152063 9560
rect 152504 9616 152596 9618
rect 152504 9560 152554 9616
rect 152504 9558 152596 9560
rect 140037 9555 140103 9558
rect 145557 9555 145623 9558
rect 151997 9555 152063 9558
rect 152549 9556 152596 9558
rect 152660 9556 152666 9620
rect 152549 9555 152615 9556
rect 19793 9482 19859 9485
rect 28625 9482 28691 9485
rect 19793 9480 28691 9482
rect 19793 9424 19798 9480
rect 19854 9424 28630 9480
rect 28686 9424 28691 9480
rect 19793 9422 28691 9424
rect 19793 9419 19859 9422
rect 28625 9419 28691 9422
rect 92749 9482 92815 9485
rect 124397 9482 124463 9485
rect 135161 9482 135227 9485
rect 92749 9480 135227 9482
rect 92749 9424 92754 9480
rect 92810 9424 124402 9480
rect 124458 9424 135166 9480
rect 135222 9424 135227 9480
rect 92749 9422 135227 9424
rect 92749 9419 92815 9422
rect 124397 9419 124463 9422
rect 135161 9419 135227 9422
rect 138013 9482 138079 9485
rect 148685 9482 148751 9485
rect 138013 9480 148751 9482
rect 138013 9424 138018 9480
rect 138074 9424 148690 9480
rect 148746 9424 148751 9480
rect 138013 9422 148751 9424
rect 138013 9419 138079 9422
rect 148685 9419 148751 9422
rect 148869 9482 148935 9485
rect 153285 9482 153351 9485
rect 148869 9480 153351 9482
rect 148869 9424 148874 9480
rect 148930 9424 153290 9480
rect 153346 9424 153351 9480
rect 148869 9422 153351 9424
rect 148869 9419 148935 9422
rect 153285 9419 153351 9422
rect 153653 9482 153719 9485
rect 156873 9482 156939 9485
rect 153653 9480 156939 9482
rect 153653 9424 153658 9480
rect 153714 9424 156878 9480
rect 156934 9424 156939 9480
rect 153653 9422 156939 9424
rect 153653 9419 153719 9422
rect 156873 9419 156939 9422
rect 42057 9346 42123 9349
rect 46289 9346 46355 9349
rect 47669 9346 47735 9349
rect 42057 9344 47735 9346
rect 42057 9288 42062 9344
rect 42118 9288 46294 9344
rect 46350 9288 47674 9344
rect 47730 9288 47735 9344
rect 42057 9286 47735 9288
rect 42057 9283 42123 9286
rect 46289 9283 46355 9286
rect 47669 9283 47735 9286
rect 87781 9346 87847 9349
rect 90449 9346 90515 9349
rect 87781 9344 90515 9346
rect 87781 9288 87786 9344
rect 87842 9288 90454 9344
rect 90510 9288 90515 9344
rect 87781 9286 90515 9288
rect 87781 9283 87847 9286
rect 90449 9283 90515 9286
rect 115565 9346 115631 9349
rect 129089 9346 129155 9349
rect 115565 9344 129155 9346
rect 115565 9288 115570 9344
rect 115626 9288 129094 9344
rect 129150 9288 129155 9344
rect 115565 9286 129155 9288
rect 115565 9283 115631 9286
rect 129089 9283 129155 9286
rect 137461 9346 137527 9349
rect 138841 9346 138907 9349
rect 137461 9344 138907 9346
rect 137461 9288 137466 9344
rect 137522 9288 138846 9344
rect 138902 9288 138907 9344
rect 137461 9286 138907 9288
rect 137461 9283 137527 9286
rect 138841 9283 138907 9286
rect 139853 9346 139919 9349
rect 142337 9346 142403 9349
rect 139853 9344 142403 9346
rect 139853 9288 139858 9344
rect 139914 9288 142342 9344
rect 142398 9288 142403 9344
rect 139853 9286 142403 9288
rect 139853 9283 139919 9286
rect 142337 9283 142403 9286
rect 143717 9346 143783 9349
rect 156045 9346 156111 9349
rect 143717 9344 156111 9346
rect 143717 9288 143722 9344
rect 143778 9288 156050 9344
rect 156106 9288 156111 9344
rect 143717 9286 156111 9288
rect 143717 9283 143783 9286
rect 156045 9283 156111 9286
rect 20668 9280 20984 9281
rect 20668 9216 20674 9280
rect 20738 9216 20754 9280
rect 20818 9216 20834 9280
rect 20898 9216 20914 9280
rect 20978 9216 20984 9280
rect 20668 9215 20984 9216
rect 60113 9280 60429 9281
rect 60113 9216 60119 9280
rect 60183 9216 60199 9280
rect 60263 9216 60279 9280
rect 60343 9216 60359 9280
rect 60423 9216 60429 9280
rect 60113 9215 60429 9216
rect 99558 9280 99874 9281
rect 99558 9216 99564 9280
rect 99628 9216 99644 9280
rect 99708 9216 99724 9280
rect 99788 9216 99804 9280
rect 99868 9216 99874 9280
rect 99558 9215 99874 9216
rect 139003 9280 139319 9281
rect 139003 9216 139009 9280
rect 139073 9216 139089 9280
rect 139153 9216 139169 9280
rect 139233 9216 139249 9280
rect 139313 9216 139319 9280
rect 139003 9215 139319 9216
rect 115289 9210 115355 9213
rect 130837 9210 130903 9213
rect 115289 9208 130903 9210
rect 115289 9152 115294 9208
rect 115350 9152 130842 9208
rect 130898 9152 130903 9208
rect 115289 9150 130903 9152
rect 115289 9147 115355 9150
rect 130837 9147 130903 9150
rect 137921 9210 137987 9213
rect 138197 9210 138263 9213
rect 137921 9208 138263 9210
rect 137921 9152 137926 9208
rect 137982 9152 138202 9208
rect 138258 9152 138263 9208
rect 137921 9150 138263 9152
rect 137921 9147 137987 9150
rect 138197 9147 138263 9150
rect 142797 9210 142863 9213
rect 148777 9210 148843 9213
rect 142797 9208 148843 9210
rect 142797 9152 142802 9208
rect 142858 9152 148782 9208
rect 148838 9152 148843 9208
rect 142797 9150 148843 9152
rect 142797 9147 142863 9150
rect 148777 9147 148843 9150
rect 149237 9210 149303 9213
rect 155861 9210 155927 9213
rect 149237 9208 155927 9210
rect 149237 9152 149242 9208
rect 149298 9152 155866 9208
rect 155922 9152 155927 9208
rect 149237 9150 155927 9152
rect 149237 9147 149303 9150
rect 155861 9147 155927 9150
rect 14273 9074 14339 9077
rect 16941 9074 17007 9077
rect 14273 9072 17007 9074
rect 14273 9016 14278 9072
rect 14334 9016 16946 9072
rect 17002 9016 17007 9072
rect 14273 9014 17007 9016
rect 14273 9011 14339 9014
rect 16941 9011 17007 9014
rect 41229 9074 41295 9077
rect 47945 9074 48011 9077
rect 41229 9072 48011 9074
rect 41229 9016 41234 9072
rect 41290 9016 47950 9072
rect 48006 9016 48011 9072
rect 41229 9014 48011 9016
rect 41229 9011 41295 9014
rect 47945 9011 48011 9014
rect 89713 9074 89779 9077
rect 90909 9074 90975 9077
rect 89713 9072 90975 9074
rect 89713 9016 89718 9072
rect 89774 9016 90914 9072
rect 90970 9016 90975 9072
rect 89713 9014 90975 9016
rect 89713 9011 89779 9014
rect 90909 9011 90975 9014
rect 93853 9074 93919 9077
rect 121821 9074 121887 9077
rect 93853 9072 121887 9074
rect 93853 9016 93858 9072
rect 93914 9016 121826 9072
rect 121882 9016 121887 9072
rect 93853 9014 121887 9016
rect 93853 9011 93919 9014
rect 121821 9011 121887 9014
rect 128261 9074 128327 9077
rect 128813 9074 128879 9077
rect 128261 9072 128879 9074
rect 128261 9016 128266 9072
rect 128322 9016 128818 9072
rect 128874 9016 128879 9072
rect 128261 9014 128879 9016
rect 128261 9011 128327 9014
rect 128813 9011 128879 9014
rect 131113 9074 131179 9077
rect 146201 9074 146267 9077
rect 148133 9074 148199 9077
rect 156137 9074 156203 9077
rect 131113 9072 146267 9074
rect 131113 9016 131118 9072
rect 131174 9016 146206 9072
rect 146262 9016 146267 9072
rect 131113 9014 146267 9016
rect 131113 9011 131179 9014
rect 146201 9011 146267 9014
rect 147262 9014 148058 9074
rect 39757 8938 39823 8941
rect 41597 8938 41663 8941
rect 39757 8936 41663 8938
rect 39757 8880 39762 8936
rect 39818 8880 41602 8936
rect 41658 8880 41663 8936
rect 39757 8878 41663 8880
rect 39757 8875 39823 8878
rect 41597 8875 41663 8878
rect 62665 8938 62731 8941
rect 95325 8938 95391 8941
rect 62665 8936 95391 8938
rect 62665 8880 62670 8936
rect 62726 8880 95330 8936
rect 95386 8880 95391 8936
rect 62665 8878 95391 8880
rect 62665 8875 62731 8878
rect 95325 8875 95391 8878
rect 100661 8938 100727 8941
rect 132125 8938 132191 8941
rect 100661 8936 132191 8938
rect 100661 8880 100666 8936
rect 100722 8880 132130 8936
rect 132186 8880 132191 8936
rect 100661 8878 132191 8880
rect 100661 8875 100727 8878
rect 132125 8875 132191 8878
rect 137369 8938 137435 8941
rect 139485 8938 139551 8941
rect 137369 8936 139551 8938
rect 137369 8880 137374 8936
rect 137430 8880 139490 8936
rect 139546 8880 139551 8936
rect 137369 8878 139551 8880
rect 137369 8875 137435 8878
rect 139485 8875 139551 8878
rect 139710 8876 139716 8940
rect 139780 8938 139786 8940
rect 145281 8938 145347 8941
rect 139780 8936 145347 8938
rect 139780 8880 145286 8936
rect 145342 8880 145347 8936
rect 139780 8878 145347 8880
rect 139780 8876 139786 8878
rect 145281 8875 145347 8878
rect 145557 8938 145623 8941
rect 147262 8938 147322 9014
rect 145557 8936 147322 8938
rect 145557 8880 145562 8936
rect 145618 8880 147322 8936
rect 145557 8878 147322 8880
rect 147397 8938 147463 8941
rect 147765 8938 147831 8941
rect 147397 8936 147831 8938
rect 147397 8880 147402 8936
rect 147458 8880 147770 8936
rect 147826 8880 147831 8936
rect 147397 8878 147831 8880
rect 147998 8938 148058 9014
rect 148133 9072 153210 9074
rect 148133 9016 148138 9072
rect 148194 9016 153210 9072
rect 148133 9014 153210 9016
rect 148133 9011 148199 9014
rect 148542 8938 148548 8940
rect 147998 8878 148548 8938
rect 145557 8875 145623 8878
rect 147397 8875 147463 8878
rect 147765 8875 147831 8878
rect 148542 8876 148548 8878
rect 148612 8876 148618 8940
rect 148685 8938 148751 8941
rect 151169 8938 151235 8941
rect 148685 8936 151235 8938
rect 148685 8880 148690 8936
rect 148746 8880 151174 8936
rect 151230 8880 151235 8936
rect 148685 8878 151235 8880
rect 153150 8938 153210 9014
rect 156094 9072 156203 9074
rect 156094 9016 156142 9072
rect 156198 9016 156203 9072
rect 156094 9011 156203 9016
rect 154798 8938 154804 8940
rect 153150 8878 154804 8938
rect 148685 8875 148751 8878
rect 151169 8875 151235 8878
rect 154798 8876 154804 8878
rect 154868 8938 154874 8940
rect 156094 8938 156154 9011
rect 154868 8878 156154 8938
rect 154868 8876 154874 8878
rect 88333 8802 88399 8805
rect 92473 8802 92539 8805
rect 93209 8802 93275 8805
rect 88333 8800 93275 8802
rect 88333 8744 88338 8800
rect 88394 8744 92478 8800
rect 92534 8744 93214 8800
rect 93270 8744 93275 8800
rect 88333 8742 93275 8744
rect 88333 8739 88399 8742
rect 92473 8739 92539 8742
rect 93209 8739 93275 8742
rect 114461 8802 114527 8805
rect 116853 8802 116919 8805
rect 114461 8800 116919 8802
rect 114461 8744 114466 8800
rect 114522 8744 116858 8800
rect 116914 8744 116919 8800
rect 114461 8742 116919 8744
rect 114461 8739 114527 8742
rect 116853 8739 116919 8742
rect 117221 8802 117287 8805
rect 119153 8802 119219 8805
rect 117221 8800 119219 8802
rect 117221 8744 117226 8800
rect 117282 8744 119158 8800
rect 119214 8744 119219 8800
rect 117221 8742 119219 8744
rect 117221 8739 117287 8742
rect 119153 8739 119219 8742
rect 122373 8802 122439 8805
rect 123753 8802 123819 8805
rect 122373 8800 123819 8802
rect 122373 8744 122378 8800
rect 122434 8744 123758 8800
rect 123814 8744 123819 8800
rect 122373 8742 123819 8744
rect 122373 8739 122439 8742
rect 123753 8739 123819 8742
rect 127198 8740 127204 8804
rect 127268 8802 127274 8804
rect 143717 8802 143783 8805
rect 127268 8800 143783 8802
rect 127268 8744 143722 8800
rect 143778 8744 143783 8800
rect 127268 8742 143783 8744
rect 127268 8740 127274 8742
rect 143717 8739 143783 8742
rect 144085 8802 144151 8805
rect 148777 8802 148843 8805
rect 144085 8800 148843 8802
rect 144085 8744 144090 8800
rect 144146 8744 148782 8800
rect 148838 8744 148843 8800
rect 144085 8742 148843 8744
rect 144085 8739 144151 8742
rect 148777 8739 148843 8742
rect 149145 8802 149211 8805
rect 150382 8802 150388 8804
rect 149145 8800 150388 8802
rect 149145 8744 149150 8800
rect 149206 8744 150388 8800
rect 149145 8742 150388 8744
rect 149145 8739 149211 8742
rect 150382 8740 150388 8742
rect 150452 8802 150458 8804
rect 150893 8802 150959 8805
rect 150452 8800 150959 8802
rect 150452 8744 150898 8800
rect 150954 8744 150959 8800
rect 150452 8742 150959 8744
rect 150452 8740 150458 8742
rect 150893 8739 150959 8742
rect 152365 8802 152431 8805
rect 155217 8802 155283 8805
rect 152365 8800 155283 8802
rect 152365 8744 152370 8800
rect 152426 8744 155222 8800
rect 155278 8744 155283 8800
rect 152365 8742 155283 8744
rect 152365 8739 152431 8742
rect 155217 8739 155283 8742
rect 40390 8736 40706 8737
rect 40390 8672 40396 8736
rect 40460 8672 40476 8736
rect 40540 8672 40556 8736
rect 40620 8672 40636 8736
rect 40700 8672 40706 8736
rect 40390 8671 40706 8672
rect 79835 8736 80151 8737
rect 79835 8672 79841 8736
rect 79905 8672 79921 8736
rect 79985 8672 80001 8736
rect 80065 8672 80081 8736
rect 80145 8672 80151 8736
rect 79835 8671 80151 8672
rect 119280 8736 119596 8737
rect 119280 8672 119286 8736
rect 119350 8672 119366 8736
rect 119430 8672 119446 8736
rect 119510 8672 119526 8736
rect 119590 8672 119596 8736
rect 119280 8671 119596 8672
rect 158725 8736 159041 8737
rect 158725 8672 158731 8736
rect 158795 8672 158811 8736
rect 158875 8672 158891 8736
rect 158955 8672 158971 8736
rect 159035 8672 159041 8736
rect 158725 8671 159041 8672
rect 91093 8666 91159 8669
rect 107653 8666 107719 8669
rect 91093 8664 107719 8666
rect 91093 8608 91098 8664
rect 91154 8608 107658 8664
rect 107714 8608 107719 8664
rect 91093 8606 107719 8608
rect 91093 8603 91159 8606
rect 107653 8603 107719 8606
rect 107837 8666 107903 8669
rect 115565 8666 115631 8669
rect 107837 8664 115631 8666
rect 107837 8608 107842 8664
rect 107898 8608 115570 8664
rect 115626 8608 115631 8664
rect 107837 8606 115631 8608
rect 107837 8603 107903 8606
rect 115565 8603 115631 8606
rect 120717 8666 120783 8669
rect 123569 8666 123635 8669
rect 120717 8664 123635 8666
rect 120717 8608 120722 8664
rect 120778 8608 123574 8664
rect 123630 8608 123635 8664
rect 120717 8606 123635 8608
rect 120717 8603 120783 8606
rect 123569 8603 123635 8606
rect 128077 8666 128143 8669
rect 136357 8666 136423 8669
rect 128077 8664 136423 8666
rect 128077 8608 128082 8664
rect 128138 8608 136362 8664
rect 136418 8608 136423 8664
rect 128077 8606 136423 8608
rect 128077 8603 128143 8606
rect 136357 8603 136423 8606
rect 141785 8666 141851 8669
rect 144821 8666 144887 8669
rect 141785 8664 144887 8666
rect 141785 8608 141790 8664
rect 141846 8608 144826 8664
rect 144882 8608 144887 8664
rect 141785 8606 144887 8608
rect 141785 8603 141851 8606
rect 144821 8603 144887 8606
rect 147070 8604 147076 8668
rect 147140 8666 147146 8668
rect 149053 8666 149119 8669
rect 149605 8668 149671 8669
rect 150157 8668 150223 8669
rect 149605 8666 149652 8668
rect 147140 8664 149119 8666
rect 147140 8608 149058 8664
rect 149114 8608 149119 8664
rect 147140 8606 149119 8608
rect 149560 8664 149652 8666
rect 149560 8608 149610 8664
rect 149560 8606 149652 8608
rect 147140 8604 147146 8606
rect 149053 8603 149119 8606
rect 149605 8604 149652 8606
rect 149716 8604 149722 8668
rect 150157 8664 150204 8668
rect 150268 8666 150274 8668
rect 150525 8666 150591 8669
rect 153561 8666 153627 8669
rect 150157 8608 150162 8664
rect 150157 8604 150204 8608
rect 150268 8606 150314 8666
rect 150525 8664 153627 8666
rect 150525 8608 150530 8664
rect 150586 8608 153566 8664
rect 153622 8608 153627 8664
rect 150525 8606 153627 8608
rect 150268 8604 150274 8606
rect 149605 8603 149671 8604
rect 150157 8603 150223 8604
rect 150525 8603 150591 8606
rect 153561 8603 153627 8606
rect 154573 8666 154639 8669
rect 156689 8666 156755 8669
rect 154573 8664 156755 8666
rect 154573 8608 154578 8664
rect 154634 8608 156694 8664
rect 156750 8608 156755 8664
rect 154573 8606 156755 8608
rect 154573 8603 154639 8606
rect 156689 8603 156755 8606
rect 21909 8530 21975 8533
rect 27705 8530 27771 8533
rect 21909 8528 27771 8530
rect 21909 8472 21914 8528
rect 21970 8472 27710 8528
rect 27766 8472 27771 8528
rect 21909 8470 27771 8472
rect 21909 8467 21975 8470
rect 27705 8467 27771 8470
rect 41045 8530 41111 8533
rect 44725 8530 44791 8533
rect 41045 8528 44791 8530
rect 41045 8472 41050 8528
rect 41106 8472 44730 8528
rect 44786 8472 44791 8528
rect 41045 8470 44791 8472
rect 41045 8467 41111 8470
rect 44725 8467 44791 8470
rect 48865 8530 48931 8533
rect 83365 8530 83431 8533
rect 48865 8528 83431 8530
rect 48865 8472 48870 8528
rect 48926 8472 83370 8528
rect 83426 8472 83431 8528
rect 48865 8470 83431 8472
rect 48865 8467 48931 8470
rect 83365 8467 83431 8470
rect 115933 8530 115999 8533
rect 118969 8530 119035 8533
rect 115933 8528 119035 8530
rect 115933 8472 115938 8528
rect 115994 8472 118974 8528
rect 119030 8472 119035 8528
rect 115933 8470 119035 8472
rect 115933 8467 115999 8470
rect 118969 8467 119035 8470
rect 120165 8530 120231 8533
rect 122925 8530 122991 8533
rect 124397 8530 124463 8533
rect 120165 8528 124463 8530
rect 120165 8472 120170 8528
rect 120226 8472 122930 8528
rect 122986 8472 124402 8528
rect 124458 8472 124463 8528
rect 120165 8470 124463 8472
rect 120165 8467 120231 8470
rect 122925 8467 122991 8470
rect 124397 8467 124463 8470
rect 126421 8530 126487 8533
rect 156965 8530 157031 8533
rect 126421 8528 157031 8530
rect 126421 8472 126426 8528
rect 126482 8472 156970 8528
rect 157026 8472 157031 8528
rect 126421 8470 157031 8472
rect 126421 8467 126487 8470
rect 156965 8467 157031 8470
rect 16757 8394 16823 8397
rect 19425 8394 19491 8397
rect 16757 8392 19491 8394
rect 16757 8336 16762 8392
rect 16818 8336 19430 8392
rect 19486 8336 19491 8392
rect 16757 8334 19491 8336
rect 16757 8331 16823 8334
rect 19425 8331 19491 8334
rect 27061 8394 27127 8397
rect 28165 8394 28231 8397
rect 27061 8392 28231 8394
rect 27061 8336 27066 8392
rect 27122 8336 28170 8392
rect 28226 8336 28231 8392
rect 27061 8334 28231 8336
rect 27061 8331 27127 8334
rect 28165 8331 28231 8334
rect 70209 8394 70275 8397
rect 115289 8394 115355 8397
rect 70209 8392 115355 8394
rect 70209 8336 70214 8392
rect 70270 8336 115294 8392
rect 115350 8336 115355 8392
rect 70209 8334 115355 8336
rect 70209 8331 70275 8334
rect 115289 8331 115355 8334
rect 116761 8394 116827 8397
rect 118417 8394 118483 8397
rect 116761 8392 118483 8394
rect 116761 8336 116766 8392
rect 116822 8336 118422 8392
rect 118478 8336 118483 8392
rect 116761 8334 118483 8336
rect 116761 8331 116827 8334
rect 118417 8331 118483 8334
rect 124254 8332 124260 8396
rect 124324 8394 124330 8396
rect 151997 8394 152063 8397
rect 124324 8392 152063 8394
rect 124324 8336 152002 8392
rect 152058 8336 152063 8392
rect 124324 8334 152063 8336
rect 124324 8332 124330 8334
rect 151997 8331 152063 8334
rect 153142 8332 153148 8396
rect 153212 8394 153218 8396
rect 154297 8394 154363 8397
rect 155401 8394 155467 8397
rect 153212 8392 154363 8394
rect 153212 8336 154302 8392
rect 154358 8336 154363 8392
rect 153212 8334 154363 8336
rect 153212 8332 153218 8334
rect 154297 8331 154363 8334
rect 154438 8392 155467 8394
rect 154438 8336 155406 8392
rect 155462 8336 155467 8392
rect 154438 8334 155467 8336
rect 110045 8258 110111 8261
rect 110045 8256 138030 8258
rect 110045 8200 110050 8256
rect 110106 8200 138030 8256
rect 110045 8198 138030 8200
rect 110045 8195 110111 8198
rect 20668 8192 20984 8193
rect 20668 8128 20674 8192
rect 20738 8128 20754 8192
rect 20818 8128 20834 8192
rect 20898 8128 20914 8192
rect 20978 8128 20984 8192
rect 20668 8127 20984 8128
rect 60113 8192 60429 8193
rect 60113 8128 60119 8192
rect 60183 8128 60199 8192
rect 60263 8128 60279 8192
rect 60343 8128 60359 8192
rect 60423 8128 60429 8192
rect 60113 8127 60429 8128
rect 99558 8192 99874 8193
rect 99558 8128 99564 8192
rect 99628 8128 99644 8192
rect 99708 8128 99724 8192
rect 99788 8128 99804 8192
rect 99868 8128 99874 8192
rect 99558 8127 99874 8128
rect 107929 8122 107995 8125
rect 112529 8122 112595 8125
rect 107929 8120 112595 8122
rect 107929 8064 107934 8120
rect 107990 8064 112534 8120
rect 112590 8064 112595 8120
rect 107929 8062 112595 8064
rect 107929 8059 107995 8062
rect 112529 8059 112595 8062
rect 113357 8122 113423 8125
rect 121361 8122 121427 8125
rect 113357 8120 121427 8122
rect 113357 8064 113362 8120
rect 113418 8064 121366 8120
rect 121422 8064 121427 8120
rect 113357 8062 121427 8064
rect 113357 8059 113423 8062
rect 121361 8059 121427 8062
rect 128905 8122 128971 8125
rect 135989 8122 136055 8125
rect 128905 8120 136055 8122
rect 128905 8064 128910 8120
rect 128966 8064 135994 8120
rect 136050 8064 136055 8120
rect 128905 8062 136055 8064
rect 128905 8059 128971 8062
rect 135989 8059 136055 8062
rect 104709 7986 104775 7989
rect 129917 7986 129983 7989
rect 104709 7984 129983 7986
rect 104709 7928 104714 7984
rect 104770 7928 129922 7984
rect 129978 7928 129983 7984
rect 104709 7926 129983 7928
rect 137970 7986 138030 8198
rect 145046 8196 145052 8260
rect 145116 8258 145122 8260
rect 148041 8258 148107 8261
rect 148910 8258 148916 8260
rect 145116 8198 147920 8258
rect 145116 8196 145122 8198
rect 139003 8192 139319 8193
rect 139003 8128 139009 8192
rect 139073 8128 139089 8192
rect 139153 8128 139169 8192
rect 139233 8128 139249 8192
rect 139313 8128 139319 8192
rect 139003 8127 139319 8128
rect 145833 8122 145899 8125
rect 147213 8124 147279 8125
rect 146886 8122 146892 8124
rect 145833 8120 146892 8122
rect 145833 8064 145838 8120
rect 145894 8064 146892 8120
rect 145833 8062 146892 8064
rect 145833 8059 145899 8062
rect 146886 8060 146892 8062
rect 146956 8060 146962 8124
rect 147213 8122 147260 8124
rect 147168 8120 147260 8122
rect 147168 8064 147218 8120
rect 147168 8062 147260 8064
rect 147213 8060 147260 8062
rect 147324 8060 147330 8124
rect 147860 8122 147920 8198
rect 148041 8256 148916 8258
rect 148041 8200 148046 8256
rect 148102 8200 148916 8256
rect 148041 8198 148916 8200
rect 148041 8195 148107 8198
rect 148910 8196 148916 8198
rect 148980 8196 148986 8260
rect 149053 8258 149119 8261
rect 150157 8258 150223 8261
rect 149053 8256 150223 8258
rect 149053 8200 149058 8256
rect 149114 8200 150162 8256
rect 150218 8200 150223 8256
rect 149053 8198 150223 8200
rect 149053 8195 149119 8198
rect 150157 8195 150223 8198
rect 150382 8196 150388 8260
rect 150452 8258 150458 8260
rect 151670 8258 151676 8260
rect 150452 8198 151676 8258
rect 150452 8196 150458 8198
rect 151670 8196 151676 8198
rect 151740 8258 151746 8260
rect 154438 8258 154498 8334
rect 155401 8331 155467 8334
rect 151740 8198 154498 8258
rect 151740 8196 151746 8198
rect 151077 8122 151143 8125
rect 147860 8120 151143 8122
rect 147860 8064 151082 8120
rect 151138 8064 151143 8120
rect 147860 8062 151143 8064
rect 147213 8059 147279 8060
rect 151077 8059 151143 8062
rect 151261 8122 151327 8125
rect 153101 8122 153167 8125
rect 151261 8120 153167 8122
rect 151261 8064 151266 8120
rect 151322 8064 153106 8120
rect 153162 8064 153167 8120
rect 151261 8062 153167 8064
rect 151261 8059 151327 8062
rect 153101 8059 153167 8062
rect 142061 7986 142127 7989
rect 137970 7984 142127 7986
rect 137970 7928 142066 7984
rect 142122 7928 142127 7984
rect 137970 7926 142127 7928
rect 104709 7923 104775 7926
rect 129917 7923 129983 7926
rect 142061 7923 142127 7926
rect 143809 7986 143875 7989
rect 156597 7986 156663 7989
rect 143809 7984 156663 7986
rect 143809 7928 143814 7984
rect 143870 7928 156602 7984
rect 156658 7928 156663 7984
rect 143809 7926 156663 7928
rect 143809 7923 143875 7926
rect 156597 7923 156663 7926
rect 158253 7986 158319 7989
rect 159200 7986 160000 8016
rect 158253 7984 160000 7986
rect 158253 7928 158258 7984
rect 158314 7928 160000 7984
rect 158253 7926 160000 7928
rect 158253 7923 158319 7926
rect 159200 7896 160000 7926
rect 90725 7850 90791 7853
rect 93761 7850 93827 7853
rect 90725 7848 93827 7850
rect 90725 7792 90730 7848
rect 90786 7792 93766 7848
rect 93822 7792 93827 7848
rect 90725 7790 93827 7792
rect 90725 7787 90791 7790
rect 93761 7787 93827 7790
rect 108849 7850 108915 7853
rect 113265 7850 113331 7853
rect 108849 7848 113331 7850
rect 108849 7792 108854 7848
rect 108910 7792 113270 7848
rect 113326 7792 113331 7848
rect 108849 7790 113331 7792
rect 108849 7787 108915 7790
rect 113265 7787 113331 7790
rect 116209 7850 116275 7853
rect 131021 7850 131087 7853
rect 116209 7848 131087 7850
rect 116209 7792 116214 7848
rect 116270 7792 131026 7848
rect 131082 7792 131087 7848
rect 116209 7790 131087 7792
rect 116209 7787 116275 7790
rect 131021 7787 131087 7790
rect 136357 7850 136423 7853
rect 154246 7850 154252 7852
rect 136357 7848 154252 7850
rect 136357 7792 136362 7848
rect 136418 7792 154252 7848
rect 136357 7790 154252 7792
rect 136357 7787 136423 7790
rect 154246 7788 154252 7790
rect 154316 7788 154322 7852
rect 90817 7714 90883 7717
rect 95141 7714 95207 7717
rect 90817 7712 95207 7714
rect 90817 7656 90822 7712
rect 90878 7656 95146 7712
rect 95202 7656 95207 7712
rect 90817 7654 95207 7656
rect 90817 7651 90883 7654
rect 95141 7651 95207 7654
rect 100385 7714 100451 7717
rect 114737 7714 114803 7717
rect 100385 7712 114803 7714
rect 100385 7656 100390 7712
rect 100446 7656 114742 7712
rect 114798 7656 114803 7712
rect 100385 7654 114803 7656
rect 100385 7651 100451 7654
rect 114737 7651 114803 7654
rect 124857 7714 124923 7717
rect 128905 7714 128971 7717
rect 124857 7712 128971 7714
rect 124857 7656 124862 7712
rect 124918 7656 128910 7712
rect 128966 7656 128971 7712
rect 124857 7654 128971 7656
rect 124857 7651 124923 7654
rect 128905 7651 128971 7654
rect 129181 7714 129247 7717
rect 141141 7714 141207 7717
rect 142061 7714 142127 7717
rect 129181 7712 142127 7714
rect 129181 7656 129186 7712
rect 129242 7656 141146 7712
rect 141202 7656 142066 7712
rect 142122 7656 142127 7712
rect 129181 7654 142127 7656
rect 129181 7651 129247 7654
rect 141141 7651 141207 7654
rect 142061 7651 142127 7654
rect 144913 7714 144979 7717
rect 155861 7714 155927 7717
rect 144913 7712 155927 7714
rect 144913 7656 144918 7712
rect 144974 7656 155866 7712
rect 155922 7656 155927 7712
rect 144913 7654 155927 7656
rect 144913 7651 144979 7654
rect 155861 7651 155927 7654
rect 40390 7648 40706 7649
rect 40390 7584 40396 7648
rect 40460 7584 40476 7648
rect 40540 7584 40556 7648
rect 40620 7584 40636 7648
rect 40700 7584 40706 7648
rect 40390 7583 40706 7584
rect 79835 7648 80151 7649
rect 79835 7584 79841 7648
rect 79905 7584 79921 7648
rect 79985 7584 80001 7648
rect 80065 7584 80081 7648
rect 80145 7584 80151 7648
rect 79835 7583 80151 7584
rect 119280 7648 119596 7649
rect 119280 7584 119286 7648
rect 119350 7584 119366 7648
rect 119430 7584 119446 7648
rect 119510 7584 119526 7648
rect 119590 7584 119596 7648
rect 119280 7583 119596 7584
rect 158725 7648 159041 7649
rect 158725 7584 158731 7648
rect 158795 7584 158811 7648
rect 158875 7584 158891 7648
rect 158955 7584 158971 7648
rect 159035 7584 159041 7648
rect 158725 7583 159041 7584
rect 89345 7578 89411 7581
rect 89805 7578 89871 7581
rect 89345 7576 89871 7578
rect 89345 7520 89350 7576
rect 89406 7520 89810 7576
rect 89866 7520 89871 7576
rect 89345 7518 89871 7520
rect 89345 7515 89411 7518
rect 89805 7515 89871 7518
rect 90817 7578 90883 7581
rect 93485 7578 93551 7581
rect 90817 7576 93551 7578
rect 90817 7520 90822 7576
rect 90878 7520 93490 7576
rect 93546 7520 93551 7576
rect 90817 7518 93551 7520
rect 90817 7515 90883 7518
rect 93485 7515 93551 7518
rect 93945 7578 94011 7581
rect 129641 7578 129707 7581
rect 93945 7576 118710 7578
rect 93945 7520 93950 7576
rect 94006 7520 118710 7576
rect 93945 7518 118710 7520
rect 93945 7515 94011 7518
rect 72877 7442 72943 7445
rect 118650 7442 118710 7518
rect 119662 7576 129707 7578
rect 119662 7520 129646 7576
rect 129702 7520 129707 7576
rect 119662 7518 129707 7520
rect 119662 7442 119722 7518
rect 129641 7515 129707 7518
rect 133873 7578 133939 7581
rect 145649 7578 145715 7581
rect 133873 7576 145715 7578
rect 133873 7520 133878 7576
rect 133934 7520 145654 7576
rect 145710 7520 145715 7576
rect 133873 7518 145715 7520
rect 133873 7515 133939 7518
rect 145649 7515 145715 7518
rect 145833 7578 145899 7581
rect 150801 7580 150867 7581
rect 145833 7576 150634 7578
rect 145833 7520 145838 7576
rect 145894 7520 150634 7576
rect 145833 7518 150634 7520
rect 145833 7515 145899 7518
rect 136633 7442 136699 7445
rect 72877 7440 109050 7442
rect 72877 7384 72882 7440
rect 72938 7384 109050 7440
rect 72877 7382 109050 7384
rect 118650 7382 119722 7442
rect 128310 7440 136699 7442
rect 128310 7384 136638 7440
rect 136694 7384 136699 7440
rect 128310 7382 136699 7384
rect 72877 7379 72943 7382
rect 91369 7306 91435 7309
rect 93853 7306 93919 7309
rect 91369 7304 93919 7306
rect 91369 7248 91374 7304
rect 91430 7248 93858 7304
rect 93914 7248 93919 7304
rect 91369 7246 93919 7248
rect 91369 7243 91435 7246
rect 93853 7243 93919 7246
rect 108990 7170 109050 7382
rect 110321 7306 110387 7309
rect 112437 7306 112503 7309
rect 110321 7304 112503 7306
rect 110321 7248 110326 7304
rect 110382 7248 112442 7304
rect 112498 7248 112503 7304
rect 110321 7246 112503 7248
rect 110321 7243 110387 7246
rect 112437 7243 112503 7246
rect 112621 7306 112687 7309
rect 126605 7306 126671 7309
rect 128310 7306 128370 7382
rect 136633 7379 136699 7382
rect 137093 7442 137159 7445
rect 141325 7442 141391 7445
rect 137093 7440 141391 7442
rect 137093 7384 137098 7440
rect 137154 7384 141330 7440
rect 141386 7384 141391 7440
rect 137093 7382 141391 7384
rect 137093 7379 137159 7382
rect 141325 7379 141391 7382
rect 141969 7442 142035 7445
rect 150382 7442 150388 7444
rect 141969 7440 150388 7442
rect 141969 7384 141974 7440
rect 142030 7384 150388 7440
rect 141969 7382 150388 7384
rect 141969 7379 142035 7382
rect 150382 7380 150388 7382
rect 150452 7380 150458 7444
rect 150574 7442 150634 7518
rect 150750 7516 150756 7580
rect 150820 7578 150867 7580
rect 151997 7578 152063 7581
rect 156965 7578 157031 7581
rect 150820 7576 150912 7578
rect 150862 7520 150912 7576
rect 150820 7518 150912 7520
rect 151997 7576 157031 7578
rect 151997 7520 152002 7576
rect 152058 7520 156970 7576
rect 157026 7520 157031 7576
rect 151997 7518 157031 7520
rect 150820 7516 150867 7518
rect 150801 7515 150867 7516
rect 151997 7515 152063 7518
rect 156965 7515 157031 7518
rect 154297 7442 154363 7445
rect 150574 7440 154363 7442
rect 150574 7384 154302 7440
rect 154358 7384 154363 7440
rect 150574 7382 154363 7384
rect 154297 7379 154363 7382
rect 112621 7304 128370 7306
rect 112621 7248 112626 7304
rect 112682 7248 126610 7304
rect 126666 7248 128370 7304
rect 112621 7246 128370 7248
rect 128537 7306 128603 7309
rect 130285 7306 130351 7309
rect 128537 7304 130351 7306
rect 128537 7248 128542 7304
rect 128598 7248 130290 7304
rect 130346 7248 130351 7304
rect 128537 7246 130351 7248
rect 112621 7243 112687 7246
rect 126605 7243 126671 7246
rect 128537 7243 128603 7246
rect 130285 7243 130351 7246
rect 130837 7306 130903 7309
rect 155953 7306 156019 7309
rect 130837 7304 156019 7306
rect 130837 7248 130842 7304
rect 130898 7248 155958 7304
rect 156014 7248 156019 7304
rect 130837 7246 156019 7248
rect 130837 7243 130903 7246
rect 155953 7243 156019 7246
rect 121821 7170 121887 7173
rect 124121 7170 124187 7173
rect 108990 7168 121887 7170
rect 108990 7112 121826 7168
rect 121882 7112 121887 7168
rect 108990 7110 121887 7112
rect 121821 7107 121887 7110
rect 122606 7168 124187 7170
rect 122606 7112 124126 7168
rect 124182 7112 124187 7168
rect 122606 7110 124187 7112
rect 20668 7104 20984 7105
rect 20668 7040 20674 7104
rect 20738 7040 20754 7104
rect 20818 7040 20834 7104
rect 20898 7040 20914 7104
rect 20978 7040 20984 7104
rect 20668 7039 20984 7040
rect 60113 7104 60429 7105
rect 60113 7040 60119 7104
rect 60183 7040 60199 7104
rect 60263 7040 60279 7104
rect 60343 7040 60359 7104
rect 60423 7040 60429 7104
rect 60113 7039 60429 7040
rect 99558 7104 99874 7105
rect 99558 7040 99564 7104
rect 99628 7040 99644 7104
rect 99708 7040 99724 7104
rect 99788 7040 99804 7104
rect 99868 7040 99874 7104
rect 99558 7039 99874 7040
rect 110597 7034 110663 7037
rect 114461 7034 114527 7037
rect 110597 7032 114527 7034
rect 110597 6976 110602 7032
rect 110658 6976 114466 7032
rect 114522 6976 114527 7032
rect 110597 6974 114527 6976
rect 110597 6971 110663 6974
rect 114461 6971 114527 6974
rect 117405 7034 117471 7037
rect 122606 7034 122666 7110
rect 124121 7107 124187 7110
rect 125501 7170 125567 7173
rect 131062 7170 131068 7172
rect 125501 7168 131068 7170
rect 125501 7112 125506 7168
rect 125562 7112 131068 7168
rect 125501 7110 131068 7112
rect 125501 7107 125567 7110
rect 131062 7108 131068 7110
rect 131132 7108 131138 7172
rect 131757 7170 131823 7173
rect 137093 7170 137159 7173
rect 131757 7168 137159 7170
rect 131757 7112 131762 7168
rect 131818 7112 137098 7168
rect 137154 7112 137159 7168
rect 131757 7110 137159 7112
rect 131757 7107 131823 7110
rect 137093 7107 137159 7110
rect 139669 7170 139735 7173
rect 140773 7170 140839 7173
rect 139669 7168 140839 7170
rect 139669 7112 139674 7168
rect 139730 7112 140778 7168
rect 140834 7112 140839 7168
rect 139669 7110 140839 7112
rect 139669 7107 139735 7110
rect 140773 7107 140839 7110
rect 142061 7170 142127 7173
rect 145833 7170 145899 7173
rect 142061 7168 145899 7170
rect 142061 7112 142066 7168
rect 142122 7112 145838 7168
rect 145894 7112 145899 7168
rect 142061 7110 145899 7112
rect 142061 7107 142127 7110
rect 145833 7107 145899 7110
rect 146886 7108 146892 7172
rect 146956 7170 146962 7172
rect 147121 7170 147187 7173
rect 146956 7168 147187 7170
rect 146956 7112 147126 7168
rect 147182 7112 147187 7168
rect 146956 7110 147187 7112
rect 146956 7108 146962 7110
rect 147121 7107 147187 7110
rect 147438 7108 147444 7172
rect 147508 7170 147514 7172
rect 147806 7170 147812 7172
rect 147508 7110 147812 7170
rect 147508 7108 147514 7110
rect 147806 7108 147812 7110
rect 147876 7108 147882 7172
rect 148041 7170 148107 7173
rect 151077 7170 151143 7173
rect 157241 7170 157307 7173
rect 148041 7168 151143 7170
rect 148041 7112 148046 7168
rect 148102 7112 151082 7168
rect 151138 7112 151143 7168
rect 148041 7110 151143 7112
rect 148041 7107 148107 7110
rect 151077 7107 151143 7110
rect 152414 7168 157307 7170
rect 152414 7112 157246 7168
rect 157302 7112 157307 7168
rect 152414 7110 157307 7112
rect 139003 7104 139319 7105
rect 139003 7040 139009 7104
rect 139073 7040 139089 7104
rect 139153 7040 139169 7104
rect 139233 7040 139249 7104
rect 139313 7040 139319 7104
rect 139003 7039 139319 7040
rect 117405 7032 122666 7034
rect 117405 6976 117410 7032
rect 117466 6976 122666 7032
rect 117405 6974 122666 6976
rect 122833 7034 122899 7037
rect 137277 7034 137343 7037
rect 122833 7032 137343 7034
rect 122833 6976 122838 7032
rect 122894 6976 137282 7032
rect 137338 6976 137343 7032
rect 122833 6974 137343 6976
rect 117405 6971 117471 6974
rect 122833 6971 122899 6974
rect 137277 6971 137343 6974
rect 142337 7034 142403 7037
rect 144821 7034 144887 7037
rect 142337 7032 144887 7034
rect 142337 6976 142342 7032
rect 142398 6976 144826 7032
rect 144882 6976 144887 7032
rect 142337 6974 144887 6976
rect 142337 6971 142403 6974
rect 144821 6971 144887 6974
rect 145005 7036 145071 7037
rect 145005 7032 145052 7036
rect 145116 7034 145122 7036
rect 145281 7034 145347 7037
rect 152414 7034 152474 7110
rect 157241 7107 157307 7110
rect 145005 6976 145010 7032
rect 145005 6972 145052 6976
rect 145116 6974 145162 7034
rect 145281 7032 152474 7034
rect 145281 6976 145286 7032
rect 145342 6976 152474 7032
rect 145281 6974 152474 6976
rect 145116 6972 145122 6974
rect 145005 6971 145071 6972
rect 145281 6971 145347 6974
rect 153326 6972 153332 7036
rect 153396 7034 153402 7036
rect 154113 7034 154179 7037
rect 153396 7032 154179 7034
rect 153396 6976 154118 7032
rect 154174 6976 154179 7032
rect 153396 6974 154179 6976
rect 153396 6972 153402 6974
rect 154113 6971 154179 6974
rect 100753 6898 100819 6901
rect 102501 6898 102567 6901
rect 133413 6900 133479 6901
rect 133413 6898 133460 6900
rect 100753 6896 133460 6898
rect 100753 6840 100758 6896
rect 100814 6840 102506 6896
rect 102562 6840 133418 6896
rect 100753 6838 133460 6840
rect 100753 6835 100819 6838
rect 102501 6835 102567 6838
rect 133413 6836 133460 6838
rect 133524 6836 133530 6900
rect 137921 6898 137987 6901
rect 141417 6898 141483 6901
rect 137921 6896 141483 6898
rect 137921 6840 137926 6896
rect 137982 6840 141422 6896
rect 141478 6840 141483 6896
rect 137921 6838 141483 6840
rect 133413 6835 133479 6836
rect 137921 6835 137987 6838
rect 141417 6835 141483 6838
rect 144177 6898 144243 6901
rect 147673 6898 147739 6901
rect 144177 6896 147739 6898
rect 144177 6840 144182 6896
rect 144238 6840 147678 6896
rect 147734 6840 147739 6896
rect 144177 6838 147739 6840
rect 144177 6835 144243 6838
rect 147673 6835 147739 6838
rect 147806 6836 147812 6900
rect 147876 6898 147882 6900
rect 153193 6898 153259 6901
rect 147876 6896 153259 6898
rect 147876 6840 153198 6896
rect 153254 6840 153259 6896
rect 147876 6838 153259 6840
rect 147876 6836 147882 6838
rect 153193 6835 153259 6838
rect 106457 6762 106523 6765
rect 114001 6762 114067 6765
rect 106457 6760 114067 6762
rect 106457 6704 106462 6760
rect 106518 6704 114006 6760
rect 114062 6704 114067 6760
rect 106457 6702 114067 6704
rect 106457 6699 106523 6702
rect 114001 6699 114067 6702
rect 114737 6762 114803 6765
rect 153469 6762 153535 6765
rect 114737 6760 153535 6762
rect 114737 6704 114742 6760
rect 114798 6704 153474 6760
rect 153530 6704 153535 6760
rect 114737 6702 153535 6704
rect 114737 6699 114803 6702
rect 153469 6699 153535 6702
rect 110597 6626 110663 6629
rect 115473 6626 115539 6629
rect 110597 6624 115539 6626
rect 110597 6568 110602 6624
rect 110658 6568 115478 6624
rect 115534 6568 115539 6624
rect 110597 6566 115539 6568
rect 110597 6563 110663 6566
rect 115473 6563 115539 6566
rect 127065 6626 127131 6629
rect 127198 6626 127204 6628
rect 127065 6624 127204 6626
rect 127065 6568 127070 6624
rect 127126 6568 127204 6624
rect 127065 6566 127204 6568
rect 127065 6563 127131 6566
rect 127198 6564 127204 6566
rect 127268 6564 127274 6628
rect 138381 6626 138447 6629
rect 140773 6626 140839 6629
rect 128310 6566 138030 6626
rect 40390 6560 40706 6561
rect 40390 6496 40396 6560
rect 40460 6496 40476 6560
rect 40540 6496 40556 6560
rect 40620 6496 40636 6560
rect 40700 6496 40706 6560
rect 40390 6495 40706 6496
rect 79835 6560 80151 6561
rect 79835 6496 79841 6560
rect 79905 6496 79921 6560
rect 79985 6496 80001 6560
rect 80065 6496 80081 6560
rect 80145 6496 80151 6560
rect 79835 6495 80151 6496
rect 119280 6560 119596 6561
rect 119280 6496 119286 6560
rect 119350 6496 119366 6560
rect 119430 6496 119446 6560
rect 119510 6496 119526 6560
rect 119590 6496 119596 6560
rect 119280 6495 119596 6496
rect 107101 6490 107167 6493
rect 115381 6490 115447 6493
rect 107101 6488 115447 6490
rect 107101 6432 107106 6488
rect 107162 6432 115386 6488
rect 115442 6432 115447 6488
rect 107101 6430 115447 6432
rect 107101 6427 107167 6430
rect 115381 6427 115447 6430
rect 120073 6490 120139 6493
rect 125961 6490 126027 6493
rect 128310 6490 128370 6566
rect 120073 6488 128370 6490
rect 120073 6432 120078 6488
rect 120134 6432 125966 6488
rect 126022 6432 128370 6488
rect 120073 6430 128370 6432
rect 137970 6490 138030 6566
rect 138381 6624 140839 6626
rect 138381 6568 138386 6624
rect 138442 6568 140778 6624
rect 140834 6568 140839 6624
rect 138381 6566 140839 6568
rect 138381 6563 138447 6566
rect 140773 6563 140839 6566
rect 142245 6626 142311 6629
rect 146477 6626 146543 6629
rect 142245 6624 146543 6626
rect 142245 6568 142250 6624
rect 142306 6568 146482 6624
rect 146538 6568 146543 6624
rect 142245 6566 146543 6568
rect 142245 6563 142311 6566
rect 146477 6563 146543 6566
rect 146753 6626 146819 6629
rect 151537 6626 151603 6629
rect 152365 6626 152431 6629
rect 146753 6624 152431 6626
rect 146753 6568 146758 6624
rect 146814 6568 151542 6624
rect 151598 6568 152370 6624
rect 152426 6568 152431 6624
rect 146753 6566 152431 6568
rect 146753 6563 146819 6566
rect 151537 6563 151603 6566
rect 152365 6563 152431 6566
rect 152549 6626 152615 6629
rect 154757 6626 154823 6629
rect 152549 6624 154823 6626
rect 152549 6568 152554 6624
rect 152610 6568 154762 6624
rect 154818 6568 154823 6624
rect 152549 6566 154823 6568
rect 152549 6563 152615 6566
rect 154757 6563 154823 6566
rect 158725 6560 159041 6561
rect 158725 6496 158731 6560
rect 158795 6496 158811 6560
rect 158875 6496 158891 6560
rect 158955 6496 158971 6560
rect 159035 6496 159041 6560
rect 158725 6495 159041 6496
rect 146334 6490 146340 6492
rect 137970 6430 146340 6490
rect 120073 6427 120139 6430
rect 125961 6427 126027 6430
rect 146334 6428 146340 6430
rect 146404 6428 146410 6492
rect 146937 6490 147003 6493
rect 152457 6490 152523 6493
rect 146937 6488 152523 6490
rect 146937 6432 146942 6488
rect 146998 6432 152462 6488
rect 152518 6432 152523 6488
rect 146937 6430 152523 6432
rect 146937 6427 147003 6430
rect 152457 6427 152523 6430
rect 91461 6354 91527 6357
rect 115381 6354 115447 6357
rect 91461 6352 115447 6354
rect 91461 6296 91466 6352
rect 91522 6296 115386 6352
rect 115442 6296 115447 6352
rect 91461 6294 115447 6296
rect 91461 6291 91527 6294
rect 115381 6291 115447 6294
rect 126513 6354 126579 6357
rect 129089 6354 129155 6357
rect 126513 6352 129155 6354
rect 126513 6296 126518 6352
rect 126574 6296 129094 6352
rect 129150 6296 129155 6352
rect 126513 6294 129155 6296
rect 126513 6291 126579 6294
rect 129089 6291 129155 6294
rect 135345 6354 135411 6357
rect 139710 6354 139716 6356
rect 135345 6352 139716 6354
rect 135345 6296 135350 6352
rect 135406 6296 139716 6352
rect 135345 6294 139716 6296
rect 135345 6291 135411 6294
rect 139710 6292 139716 6294
rect 139780 6292 139786 6356
rect 141141 6354 141207 6357
rect 143809 6354 143875 6357
rect 141141 6352 143875 6354
rect 141141 6296 141146 6352
rect 141202 6296 143814 6352
rect 143870 6296 143875 6352
rect 141141 6294 143875 6296
rect 141141 6291 141207 6294
rect 143809 6291 143875 6294
rect 144545 6354 144611 6357
rect 150433 6354 150499 6357
rect 144545 6352 150499 6354
rect 144545 6296 144550 6352
rect 144606 6296 150438 6352
rect 150494 6296 150499 6352
rect 144545 6294 150499 6296
rect 144545 6291 144611 6294
rect 150433 6291 150499 6294
rect 153561 6354 153627 6357
rect 154849 6354 154915 6357
rect 153561 6352 154915 6354
rect 153561 6296 153566 6352
rect 153622 6296 154854 6352
rect 154910 6296 154915 6352
rect 153561 6294 154915 6296
rect 153561 6291 153627 6294
rect 154849 6291 154915 6294
rect 10317 6218 10383 6221
rect 29361 6218 29427 6221
rect 10317 6216 29427 6218
rect 10317 6160 10322 6216
rect 10378 6160 29366 6216
rect 29422 6160 29427 6216
rect 10317 6158 29427 6160
rect 10317 6155 10383 6158
rect 29361 6155 29427 6158
rect 100293 6218 100359 6221
rect 124397 6218 124463 6221
rect 133873 6218 133939 6221
rect 100293 6216 133939 6218
rect 100293 6160 100298 6216
rect 100354 6160 124402 6216
rect 124458 6160 133878 6216
rect 133934 6160 133939 6216
rect 100293 6158 133939 6160
rect 100293 6155 100359 6158
rect 124397 6155 124463 6158
rect 133873 6155 133939 6158
rect 134425 6218 134491 6221
rect 147857 6218 147923 6221
rect 134425 6216 147923 6218
rect 134425 6160 134430 6216
rect 134486 6160 147862 6216
rect 147918 6160 147923 6216
rect 134425 6158 147923 6160
rect 134425 6155 134491 6158
rect 147857 6155 147923 6158
rect 149278 6156 149284 6220
rect 149348 6218 149354 6220
rect 149881 6218 149947 6221
rect 149348 6216 149947 6218
rect 149348 6160 149886 6216
rect 149942 6160 149947 6216
rect 149348 6158 149947 6160
rect 149348 6156 149354 6158
rect 149881 6155 149947 6158
rect 150249 6218 150315 6221
rect 150985 6218 151051 6221
rect 150249 6216 151051 6218
rect 150249 6160 150254 6216
rect 150310 6160 150990 6216
rect 151046 6160 151051 6216
rect 150249 6158 151051 6160
rect 150249 6155 150315 6158
rect 150985 6155 151051 6158
rect 153929 6218 153995 6221
rect 155217 6218 155283 6221
rect 153929 6216 155283 6218
rect 153929 6160 153934 6216
rect 153990 6160 155222 6216
rect 155278 6160 155283 6216
rect 153929 6158 155283 6160
rect 153929 6155 153995 6158
rect 155217 6155 155283 6158
rect 101857 6082 101923 6085
rect 122741 6082 122807 6085
rect 129733 6082 129799 6085
rect 101857 6080 122807 6082
rect 101857 6024 101862 6080
rect 101918 6024 122746 6080
rect 122802 6024 122807 6080
rect 101857 6022 122807 6024
rect 101857 6019 101923 6022
rect 122741 6019 122807 6022
rect 125550 6080 129799 6082
rect 125550 6024 129738 6080
rect 129794 6024 129799 6080
rect 125550 6022 129799 6024
rect 20668 6016 20984 6017
rect 0 5946 800 5976
rect 20668 5952 20674 6016
rect 20738 5952 20754 6016
rect 20818 5952 20834 6016
rect 20898 5952 20914 6016
rect 20978 5952 20984 6016
rect 20668 5951 20984 5952
rect 60113 6016 60429 6017
rect 60113 5952 60119 6016
rect 60183 5952 60199 6016
rect 60263 5952 60279 6016
rect 60343 5952 60359 6016
rect 60423 5952 60429 6016
rect 60113 5951 60429 5952
rect 99558 6016 99874 6017
rect 99558 5952 99564 6016
rect 99628 5952 99644 6016
rect 99708 5952 99724 6016
rect 99788 5952 99804 6016
rect 99868 5952 99874 6016
rect 99558 5951 99874 5952
rect 1577 5946 1643 5949
rect 0 5944 1643 5946
rect 0 5888 1582 5944
rect 1638 5888 1643 5944
rect 0 5886 1643 5888
rect 0 5856 800 5886
rect 1577 5883 1643 5886
rect 106917 5946 106983 5949
rect 111977 5946 112043 5949
rect 106917 5944 112043 5946
rect 106917 5888 106922 5944
rect 106978 5888 111982 5944
rect 112038 5888 112043 5944
rect 106917 5886 112043 5888
rect 106917 5883 106983 5886
rect 111977 5883 112043 5886
rect 117405 5946 117471 5949
rect 124254 5946 124260 5948
rect 117405 5944 124260 5946
rect 117405 5888 117410 5944
rect 117466 5888 124260 5944
rect 117405 5886 124260 5888
rect 117405 5883 117471 5886
rect 124254 5884 124260 5886
rect 124324 5884 124330 5948
rect 125550 5946 125610 6022
rect 129733 6019 129799 6022
rect 129917 6082 129983 6085
rect 134428 6082 134488 6155
rect 129917 6080 134488 6082
rect 129917 6024 129922 6080
rect 129978 6024 134488 6080
rect 129917 6022 134488 6024
rect 139577 6082 139643 6085
rect 156689 6082 156755 6085
rect 139577 6080 156755 6082
rect 139577 6024 139582 6080
rect 139638 6024 156694 6080
rect 156750 6024 156755 6080
rect 139577 6022 156755 6024
rect 129917 6019 129983 6022
rect 139577 6019 139643 6022
rect 156689 6019 156755 6022
rect 139003 6016 139319 6017
rect 139003 5952 139009 6016
rect 139073 5952 139089 6016
rect 139153 5952 139169 6016
rect 139233 5952 139249 6016
rect 139313 5952 139319 6016
rect 139003 5951 139319 5952
rect 124400 5886 125610 5946
rect 128169 5946 128235 5949
rect 131297 5946 131363 5949
rect 128169 5944 131363 5946
rect 128169 5888 128174 5944
rect 128230 5888 131302 5944
rect 131358 5888 131363 5944
rect 128169 5886 131363 5888
rect 116945 5810 117011 5813
rect 124400 5810 124460 5886
rect 128169 5883 128235 5886
rect 131297 5883 131363 5886
rect 142153 5946 142219 5949
rect 145189 5946 145255 5949
rect 142153 5944 145255 5946
rect 142153 5888 142158 5944
rect 142214 5888 145194 5944
rect 145250 5888 145255 5944
rect 142153 5886 145255 5888
rect 142153 5883 142219 5886
rect 145189 5883 145255 5886
rect 145649 5946 145715 5949
rect 147029 5946 147095 5949
rect 145649 5944 147095 5946
rect 145649 5888 145654 5944
rect 145710 5888 147034 5944
rect 147090 5888 147095 5944
rect 145649 5886 147095 5888
rect 145649 5883 145715 5886
rect 147029 5883 147095 5886
rect 148317 5946 148383 5949
rect 155309 5946 155375 5949
rect 148317 5944 155375 5946
rect 148317 5888 148322 5944
rect 148378 5888 155314 5944
rect 155370 5888 155375 5944
rect 148317 5886 155375 5888
rect 148317 5883 148383 5886
rect 155309 5883 155375 5886
rect 116945 5808 124460 5810
rect 116945 5752 116950 5808
rect 117006 5752 124460 5808
rect 116945 5750 124460 5752
rect 124581 5810 124647 5813
rect 125685 5810 125751 5813
rect 124581 5808 125751 5810
rect 124581 5752 124586 5808
rect 124642 5752 125690 5808
rect 125746 5752 125751 5808
rect 124581 5750 125751 5752
rect 116945 5747 117011 5750
rect 124581 5747 124647 5750
rect 125685 5747 125751 5750
rect 137737 5810 137803 5813
rect 154665 5810 154731 5813
rect 137737 5808 154731 5810
rect 137737 5752 137742 5808
rect 137798 5752 154670 5808
rect 154726 5752 154731 5808
rect 137737 5750 154731 5752
rect 137737 5747 137803 5750
rect 154665 5747 154731 5750
rect 22093 5674 22159 5677
rect 30373 5674 30439 5677
rect 22093 5672 30439 5674
rect 22093 5616 22098 5672
rect 22154 5616 30378 5672
rect 30434 5616 30439 5672
rect 22093 5614 30439 5616
rect 22093 5611 22159 5614
rect 30373 5611 30439 5614
rect 107377 5674 107443 5677
rect 113725 5674 113791 5677
rect 107377 5672 113791 5674
rect 107377 5616 107382 5672
rect 107438 5616 113730 5672
rect 113786 5616 113791 5672
rect 107377 5614 113791 5616
rect 107377 5611 107443 5614
rect 113725 5611 113791 5614
rect 115381 5674 115447 5677
rect 134517 5674 134583 5677
rect 146937 5674 147003 5677
rect 115381 5672 147003 5674
rect 115381 5616 115386 5672
rect 115442 5616 134522 5672
rect 134578 5616 146942 5672
rect 146998 5616 147003 5672
rect 115381 5614 147003 5616
rect 115381 5611 115447 5614
rect 134517 5611 134583 5614
rect 146937 5611 147003 5614
rect 147305 5674 147371 5677
rect 149513 5674 149579 5677
rect 147305 5672 149579 5674
rect 147305 5616 147310 5672
rect 147366 5616 149518 5672
rect 149574 5616 149579 5672
rect 147305 5614 149579 5616
rect 147305 5611 147371 5614
rect 149513 5611 149579 5614
rect 149697 5674 149763 5677
rect 150198 5674 150204 5676
rect 149697 5672 150204 5674
rect 149697 5616 149702 5672
rect 149758 5616 150204 5672
rect 149697 5614 150204 5616
rect 149697 5611 149763 5614
rect 150198 5612 150204 5614
rect 150268 5612 150274 5676
rect 151854 5612 151860 5676
rect 151924 5674 151930 5676
rect 155493 5674 155559 5677
rect 155953 5676 156019 5677
rect 155902 5674 155908 5676
rect 151924 5672 155559 5674
rect 151924 5616 155498 5672
rect 155554 5616 155559 5672
rect 151924 5614 155559 5616
rect 155862 5614 155908 5674
rect 155972 5672 156019 5676
rect 156014 5616 156019 5672
rect 151924 5612 151930 5614
rect 155493 5611 155559 5614
rect 155902 5612 155908 5614
rect 155972 5612 156019 5616
rect 155953 5611 156019 5612
rect 123109 5538 123175 5541
rect 125869 5538 125935 5541
rect 123109 5536 125935 5538
rect 123109 5480 123114 5536
rect 123170 5480 125874 5536
rect 125930 5480 125935 5536
rect 123109 5478 125935 5480
rect 123109 5475 123175 5478
rect 125869 5475 125935 5478
rect 129733 5538 129799 5541
rect 141969 5538 142035 5541
rect 129733 5536 142035 5538
rect 129733 5480 129738 5536
rect 129794 5480 141974 5536
rect 142030 5480 142035 5536
rect 129733 5478 142035 5480
rect 129733 5475 129799 5478
rect 141969 5475 142035 5478
rect 145281 5538 145347 5541
rect 147254 5538 147260 5540
rect 145281 5536 147260 5538
rect 145281 5480 145286 5536
rect 145342 5480 147260 5536
rect 145281 5478 147260 5480
rect 145281 5475 145347 5478
rect 147254 5476 147260 5478
rect 147324 5538 147330 5540
rect 152457 5538 152523 5541
rect 147324 5536 152523 5538
rect 147324 5480 152462 5536
rect 152518 5480 152523 5536
rect 147324 5478 152523 5480
rect 147324 5476 147330 5478
rect 152457 5475 152523 5478
rect 154297 5538 154363 5541
rect 157057 5538 157123 5541
rect 154297 5536 157123 5538
rect 154297 5480 154302 5536
rect 154358 5480 157062 5536
rect 157118 5480 157123 5536
rect 154297 5478 157123 5480
rect 154297 5475 154363 5478
rect 157057 5475 157123 5478
rect 40390 5472 40706 5473
rect 40390 5408 40396 5472
rect 40460 5408 40476 5472
rect 40540 5408 40556 5472
rect 40620 5408 40636 5472
rect 40700 5408 40706 5472
rect 40390 5407 40706 5408
rect 79835 5472 80151 5473
rect 79835 5408 79841 5472
rect 79905 5408 79921 5472
rect 79985 5408 80001 5472
rect 80065 5408 80081 5472
rect 80145 5408 80151 5472
rect 79835 5407 80151 5408
rect 119280 5472 119596 5473
rect 119280 5408 119286 5472
rect 119350 5408 119366 5472
rect 119430 5408 119446 5472
rect 119510 5408 119526 5472
rect 119590 5408 119596 5472
rect 119280 5407 119596 5408
rect 158725 5472 159041 5473
rect 158725 5408 158731 5472
rect 158795 5408 158811 5472
rect 158875 5408 158891 5472
rect 158955 5408 158971 5472
rect 159035 5408 159041 5472
rect 158725 5407 159041 5408
rect 16297 5402 16363 5405
rect 17309 5402 17375 5405
rect 16297 5400 17375 5402
rect 16297 5344 16302 5400
rect 16358 5344 17314 5400
rect 17370 5344 17375 5400
rect 16297 5342 17375 5344
rect 16297 5339 16363 5342
rect 17309 5339 17375 5342
rect 126973 5402 127039 5405
rect 147990 5402 147996 5404
rect 126973 5400 147996 5402
rect 126973 5344 126978 5400
rect 127034 5344 147996 5400
rect 126973 5342 147996 5344
rect 126973 5339 127039 5342
rect 147990 5340 147996 5342
rect 148060 5402 148066 5404
rect 151997 5402 152063 5405
rect 156781 5404 156847 5405
rect 156781 5402 156828 5404
rect 148060 5400 152063 5402
rect 148060 5344 152002 5400
rect 152058 5344 152063 5400
rect 148060 5342 152063 5344
rect 156736 5400 156828 5402
rect 156736 5344 156786 5400
rect 156736 5342 156828 5344
rect 148060 5340 148066 5342
rect 151997 5339 152063 5342
rect 156781 5340 156828 5342
rect 156892 5340 156898 5404
rect 156781 5339 156847 5340
rect 99925 5266 99991 5269
rect 127157 5266 127223 5269
rect 99925 5264 127223 5266
rect 99925 5208 99930 5264
rect 99986 5208 127162 5264
rect 127218 5208 127223 5264
rect 99925 5206 127223 5208
rect 99925 5203 99991 5206
rect 127157 5203 127223 5206
rect 139485 5266 139551 5269
rect 148225 5266 148291 5269
rect 139485 5264 148291 5266
rect 139485 5208 139490 5264
rect 139546 5208 148230 5264
rect 148286 5208 148291 5264
rect 139485 5206 148291 5208
rect 139485 5203 139551 5206
rect 148225 5203 148291 5206
rect 148910 5204 148916 5268
rect 148980 5266 148986 5268
rect 151077 5266 151143 5269
rect 148980 5264 151143 5266
rect 148980 5208 151082 5264
rect 151138 5208 151143 5264
rect 148980 5206 151143 5208
rect 148980 5204 148986 5206
rect 151077 5203 151143 5206
rect 151353 5266 151419 5269
rect 155493 5266 155559 5269
rect 151353 5264 155559 5266
rect 151353 5208 151358 5264
rect 151414 5208 155498 5264
rect 155554 5208 155559 5264
rect 151353 5206 155559 5208
rect 151353 5203 151419 5206
rect 155493 5203 155559 5206
rect 100017 5130 100083 5133
rect 140589 5130 140655 5133
rect 100017 5128 140655 5130
rect 100017 5072 100022 5128
rect 100078 5072 140594 5128
rect 140650 5072 140655 5128
rect 100017 5070 140655 5072
rect 100017 5067 100083 5070
rect 140589 5067 140655 5070
rect 146937 5130 147003 5133
rect 147070 5130 147076 5132
rect 146937 5128 147076 5130
rect 146937 5072 146942 5128
rect 146998 5072 147076 5128
rect 146937 5070 147076 5072
rect 146937 5067 147003 5070
rect 147070 5068 147076 5070
rect 147140 5068 147146 5132
rect 147305 5130 147371 5133
rect 152273 5130 152339 5133
rect 154297 5132 154363 5133
rect 147305 5128 152339 5130
rect 147305 5072 147310 5128
rect 147366 5072 152278 5128
rect 152334 5072 152339 5128
rect 147305 5070 152339 5072
rect 147305 5067 147371 5070
rect 152273 5067 152339 5070
rect 154246 5068 154252 5132
rect 154316 5130 154363 5132
rect 154316 5128 154408 5130
rect 154358 5072 154408 5128
rect 154316 5070 154408 5072
rect 154316 5068 154363 5070
rect 154297 5067 154363 5068
rect 139577 4994 139643 4997
rect 146293 4994 146359 4997
rect 139577 4992 146359 4994
rect 139577 4936 139582 4992
rect 139638 4936 146298 4992
rect 146354 4936 146359 4992
rect 139577 4934 146359 4936
rect 139577 4931 139643 4934
rect 146293 4931 146359 4934
rect 146477 4994 146543 4997
rect 157609 4994 157675 4997
rect 146477 4992 157675 4994
rect 146477 4936 146482 4992
rect 146538 4936 157614 4992
rect 157670 4936 157675 4992
rect 146477 4934 157675 4936
rect 146477 4931 146543 4934
rect 157609 4931 157675 4934
rect 20668 4928 20984 4929
rect 20668 4864 20674 4928
rect 20738 4864 20754 4928
rect 20818 4864 20834 4928
rect 20898 4864 20914 4928
rect 20978 4864 20984 4928
rect 20668 4863 20984 4864
rect 60113 4928 60429 4929
rect 60113 4864 60119 4928
rect 60183 4864 60199 4928
rect 60263 4864 60279 4928
rect 60343 4864 60359 4928
rect 60423 4864 60429 4928
rect 60113 4863 60429 4864
rect 99558 4928 99874 4929
rect 99558 4864 99564 4928
rect 99628 4864 99644 4928
rect 99708 4864 99724 4928
rect 99788 4864 99804 4928
rect 99868 4864 99874 4928
rect 99558 4863 99874 4864
rect 139003 4928 139319 4929
rect 139003 4864 139009 4928
rect 139073 4864 139089 4928
rect 139153 4864 139169 4928
rect 139233 4864 139249 4928
rect 139313 4864 139319 4928
rect 139003 4863 139319 4864
rect 117221 4858 117287 4861
rect 118693 4858 118759 4861
rect 117221 4856 118759 4858
rect 117221 4800 117226 4856
rect 117282 4800 118698 4856
rect 118754 4800 118759 4856
rect 117221 4798 118759 4800
rect 117221 4795 117287 4798
rect 118693 4795 118759 4798
rect 146017 4858 146083 4861
rect 156045 4858 156111 4861
rect 146017 4856 156111 4858
rect 146017 4800 146022 4856
rect 146078 4800 156050 4856
rect 156106 4800 156111 4856
rect 146017 4798 156111 4800
rect 146017 4795 146083 4798
rect 156045 4795 156111 4798
rect 117773 4722 117839 4725
rect 122741 4722 122807 4725
rect 117773 4720 122807 4722
rect 117773 4664 117778 4720
rect 117834 4664 122746 4720
rect 122802 4664 122807 4720
rect 117773 4662 122807 4664
rect 117773 4659 117839 4662
rect 122741 4659 122807 4662
rect 128905 4722 128971 4725
rect 152089 4722 152155 4725
rect 128905 4720 152155 4722
rect 128905 4664 128910 4720
rect 128966 4664 152094 4720
rect 152150 4664 152155 4720
rect 128905 4662 152155 4664
rect 128905 4659 128971 4662
rect 152089 4659 152155 4662
rect 76373 4586 76439 4589
rect 130193 4586 130259 4589
rect 76373 4584 130259 4586
rect 76373 4528 76378 4584
rect 76434 4528 130198 4584
rect 130254 4528 130259 4584
rect 76373 4526 130259 4528
rect 76373 4523 76439 4526
rect 130193 4523 130259 4526
rect 137829 4586 137895 4589
rect 140037 4586 140103 4589
rect 137829 4584 140103 4586
rect 137829 4528 137834 4584
rect 137890 4528 140042 4584
rect 140098 4528 140103 4584
rect 137829 4526 140103 4528
rect 137829 4523 137895 4526
rect 140037 4523 140103 4526
rect 141049 4586 141115 4589
rect 151261 4586 151327 4589
rect 152917 4586 152983 4589
rect 141049 4584 150266 4586
rect 141049 4528 141054 4584
rect 141110 4528 150266 4584
rect 141049 4526 150266 4528
rect 141049 4523 141115 4526
rect 109217 4450 109283 4453
rect 115381 4450 115447 4453
rect 109217 4448 115447 4450
rect 109217 4392 109222 4448
rect 109278 4392 115386 4448
rect 115442 4392 115447 4448
rect 109217 4390 115447 4392
rect 109217 4387 109283 4390
rect 115381 4387 115447 4390
rect 120349 4450 120415 4453
rect 140681 4450 140747 4453
rect 120349 4448 140747 4450
rect 120349 4392 120354 4448
rect 120410 4392 140686 4448
rect 140742 4392 140747 4448
rect 120349 4390 140747 4392
rect 120349 4387 120415 4390
rect 140681 4387 140747 4390
rect 145557 4450 145623 4453
rect 146937 4450 147003 4453
rect 149789 4450 149855 4453
rect 145557 4448 147003 4450
rect 145557 4392 145562 4448
rect 145618 4392 146942 4448
rect 146998 4392 147003 4448
rect 145557 4390 147003 4392
rect 145557 4387 145623 4390
rect 146937 4387 147003 4390
rect 147078 4448 149855 4450
rect 147078 4392 149794 4448
rect 149850 4392 149855 4448
rect 147078 4390 149855 4392
rect 150206 4450 150266 4526
rect 151261 4584 152983 4586
rect 151261 4528 151266 4584
rect 151322 4528 152922 4584
rect 152978 4528 152983 4584
rect 151261 4526 152983 4528
rect 151261 4523 151327 4526
rect 152917 4523 152983 4526
rect 150893 4450 150959 4453
rect 150206 4448 150959 4450
rect 150206 4392 150898 4448
rect 150954 4392 150959 4448
rect 150206 4390 150959 4392
rect 40390 4384 40706 4385
rect 40390 4320 40396 4384
rect 40460 4320 40476 4384
rect 40540 4320 40556 4384
rect 40620 4320 40636 4384
rect 40700 4320 40706 4384
rect 40390 4319 40706 4320
rect 79835 4384 80151 4385
rect 79835 4320 79841 4384
rect 79905 4320 79921 4384
rect 79985 4320 80001 4384
rect 80065 4320 80081 4384
rect 80145 4320 80151 4384
rect 79835 4319 80151 4320
rect 119280 4384 119596 4385
rect 119280 4320 119286 4384
rect 119350 4320 119366 4384
rect 119430 4320 119446 4384
rect 119510 4320 119526 4384
rect 119590 4320 119596 4384
rect 119280 4319 119596 4320
rect 126605 4314 126671 4317
rect 127985 4314 128051 4317
rect 126605 4312 128051 4314
rect 126605 4256 126610 4312
rect 126666 4256 127990 4312
rect 128046 4256 128051 4312
rect 126605 4254 128051 4256
rect 126605 4251 126671 4254
rect 127985 4251 128051 4254
rect 130837 4314 130903 4317
rect 133965 4314 134031 4317
rect 130837 4312 134031 4314
rect 130837 4256 130842 4312
rect 130898 4256 133970 4312
rect 134026 4256 134031 4312
rect 130837 4254 134031 4256
rect 130837 4251 130903 4254
rect 133965 4251 134031 4254
rect 137921 4314 137987 4317
rect 143073 4314 143139 4317
rect 137921 4312 143139 4314
rect 137921 4256 137926 4312
rect 137982 4256 143078 4312
rect 143134 4256 143139 4312
rect 137921 4254 143139 4256
rect 137921 4251 137987 4254
rect 143073 4251 143139 4254
rect 143625 4314 143691 4317
rect 145557 4314 145623 4317
rect 143625 4312 145623 4314
rect 143625 4256 143630 4312
rect 143686 4256 145562 4312
rect 145618 4256 145623 4312
rect 143625 4254 145623 4256
rect 143625 4251 143691 4254
rect 145557 4251 145623 4254
rect 145925 4314 145991 4317
rect 147078 4314 147138 4390
rect 149789 4387 149855 4390
rect 150893 4387 150959 4390
rect 158725 4384 159041 4385
rect 158725 4320 158731 4384
rect 158795 4320 158811 4384
rect 158875 4320 158891 4384
rect 158955 4320 158971 4384
rect 159035 4320 159041 4384
rect 158725 4319 159041 4320
rect 145925 4312 147138 4314
rect 145925 4256 145930 4312
rect 145986 4256 147138 4312
rect 145925 4254 147138 4256
rect 147949 4314 148015 4317
rect 153142 4314 153148 4316
rect 147949 4312 153148 4314
rect 147949 4256 147954 4312
rect 148010 4256 153148 4312
rect 147949 4254 153148 4256
rect 145925 4251 145991 4254
rect 147949 4251 148015 4254
rect 153142 4252 153148 4254
rect 153212 4252 153218 4316
rect 155217 4314 155283 4317
rect 155174 4312 155283 4314
rect 155174 4256 155222 4312
rect 155278 4256 155283 4312
rect 155174 4251 155283 4256
rect 112713 4178 112779 4181
rect 131113 4178 131179 4181
rect 112713 4176 131179 4178
rect 112713 4120 112718 4176
rect 112774 4120 131118 4176
rect 131174 4120 131179 4176
rect 112713 4118 131179 4120
rect 112713 4115 112779 4118
rect 131113 4115 131179 4118
rect 132033 4178 132099 4181
rect 133137 4178 133203 4181
rect 133597 4178 133663 4181
rect 132033 4176 133663 4178
rect 132033 4120 132038 4176
rect 132094 4120 133142 4176
rect 133198 4120 133602 4176
rect 133658 4120 133663 4176
rect 132033 4118 133663 4120
rect 132033 4115 132099 4118
rect 133137 4115 133203 4118
rect 133597 4115 133663 4118
rect 138289 4178 138355 4181
rect 139945 4178 140011 4181
rect 138289 4176 140011 4178
rect 138289 4120 138294 4176
rect 138350 4120 139950 4176
rect 140006 4120 140011 4176
rect 138289 4118 140011 4120
rect 138289 4115 138355 4118
rect 139945 4115 140011 4118
rect 140129 4178 140195 4181
rect 144729 4178 144795 4181
rect 140129 4176 144795 4178
rect 140129 4120 140134 4176
rect 140190 4120 144734 4176
rect 144790 4120 144795 4176
rect 140129 4118 144795 4120
rect 140129 4115 140195 4118
rect 144729 4115 144795 4118
rect 144913 4178 144979 4181
rect 145649 4178 145715 4181
rect 144913 4176 145715 4178
rect 144913 4120 144918 4176
rect 144974 4120 145654 4176
rect 145710 4120 145715 4176
rect 144913 4118 145715 4120
rect 144913 4115 144979 4118
rect 145649 4115 145715 4118
rect 147029 4178 147095 4181
rect 152590 4178 152596 4180
rect 147029 4176 152596 4178
rect 147029 4120 147034 4176
rect 147090 4120 152596 4176
rect 147029 4118 152596 4120
rect 147029 4115 147095 4118
rect 152590 4116 152596 4118
rect 152660 4178 152666 4180
rect 155174 4178 155234 4251
rect 152660 4118 155234 4178
rect 152660 4116 152666 4118
rect 115289 4042 115355 4045
rect 125225 4042 125291 4045
rect 115289 4040 125291 4042
rect 115289 3984 115294 4040
rect 115350 3984 125230 4040
rect 125286 3984 125291 4040
rect 115289 3982 125291 3984
rect 115289 3979 115355 3982
rect 125225 3979 125291 3982
rect 128629 4042 128695 4045
rect 141785 4042 141851 4045
rect 149053 4042 149119 4045
rect 128629 4040 149119 4042
rect 128629 3984 128634 4040
rect 128690 3984 141790 4040
rect 141846 3984 149058 4040
rect 149114 3984 149119 4040
rect 128629 3982 149119 3984
rect 128629 3979 128695 3982
rect 141785 3979 141851 3982
rect 149053 3979 149119 3982
rect 149237 4042 149303 4045
rect 153561 4042 153627 4045
rect 155125 4044 155191 4045
rect 155769 4044 155835 4045
rect 155125 4042 155172 4044
rect 149237 4040 153627 4042
rect 149237 3984 149242 4040
rect 149298 3984 153566 4040
rect 153622 3984 153627 4040
rect 149237 3982 153627 3984
rect 155080 4040 155172 4042
rect 155080 3984 155130 4040
rect 155080 3982 155172 3984
rect 149237 3979 149303 3982
rect 153561 3979 153627 3982
rect 155125 3980 155172 3982
rect 155236 3980 155242 4044
rect 155718 4042 155724 4044
rect 155678 3982 155724 4042
rect 155788 4040 155835 4044
rect 155830 3984 155835 4040
rect 155718 3980 155724 3982
rect 155788 3980 155835 3984
rect 155125 3979 155191 3980
rect 155769 3979 155835 3980
rect 105997 3906 106063 3909
rect 133689 3906 133755 3909
rect 105997 3904 133755 3906
rect 105997 3848 106002 3904
rect 106058 3848 133694 3904
rect 133750 3848 133755 3904
rect 105997 3846 133755 3848
rect 105997 3843 106063 3846
rect 133689 3843 133755 3846
rect 146201 3906 146267 3909
rect 156781 3906 156847 3909
rect 146201 3904 156847 3906
rect 146201 3848 146206 3904
rect 146262 3848 156786 3904
rect 156842 3848 156847 3904
rect 146201 3846 156847 3848
rect 146201 3843 146267 3846
rect 156781 3843 156847 3846
rect 20668 3840 20984 3841
rect 20668 3776 20674 3840
rect 20738 3776 20754 3840
rect 20818 3776 20834 3840
rect 20898 3776 20914 3840
rect 20978 3776 20984 3840
rect 20668 3775 20984 3776
rect 60113 3840 60429 3841
rect 60113 3776 60119 3840
rect 60183 3776 60199 3840
rect 60263 3776 60279 3840
rect 60343 3776 60359 3840
rect 60423 3776 60429 3840
rect 60113 3775 60429 3776
rect 99558 3840 99874 3841
rect 99558 3776 99564 3840
rect 99628 3776 99644 3840
rect 99708 3776 99724 3840
rect 99788 3776 99804 3840
rect 99868 3776 99874 3840
rect 99558 3775 99874 3776
rect 139003 3840 139319 3841
rect 139003 3776 139009 3840
rect 139073 3776 139089 3840
rect 139153 3776 139169 3840
rect 139233 3776 139249 3840
rect 139313 3776 139319 3840
rect 139003 3775 139319 3776
rect 118233 3770 118299 3773
rect 119245 3770 119311 3773
rect 118233 3768 119311 3770
rect 118233 3712 118238 3768
rect 118294 3712 119250 3768
rect 119306 3712 119311 3768
rect 118233 3710 119311 3712
rect 118233 3707 118299 3710
rect 119245 3707 119311 3710
rect 128353 3770 128419 3773
rect 132769 3770 132835 3773
rect 128353 3768 132835 3770
rect 128353 3712 128358 3768
rect 128414 3712 132774 3768
rect 132830 3712 132835 3768
rect 128353 3710 132835 3712
rect 128353 3707 128419 3710
rect 132769 3707 132835 3710
rect 140681 3770 140747 3773
rect 146293 3770 146359 3773
rect 152825 3772 152891 3773
rect 151854 3770 151860 3772
rect 140681 3768 151860 3770
rect 140681 3712 140686 3768
rect 140742 3712 146298 3768
rect 146354 3712 151860 3768
rect 140681 3710 151860 3712
rect 140681 3707 140747 3710
rect 146293 3707 146359 3710
rect 151854 3708 151860 3710
rect 151924 3708 151930 3772
rect 152774 3708 152780 3772
rect 152844 3770 152891 3772
rect 153009 3770 153075 3773
rect 154665 3770 154731 3773
rect 152844 3768 152936 3770
rect 152886 3712 152936 3768
rect 152844 3710 152936 3712
rect 153009 3768 154731 3770
rect 153009 3712 153014 3768
rect 153070 3712 154670 3768
rect 154726 3712 154731 3768
rect 153009 3710 154731 3712
rect 152844 3708 152891 3710
rect 152825 3707 152891 3708
rect 153009 3707 153075 3710
rect 154665 3707 154731 3710
rect 154798 3708 154804 3772
rect 154868 3770 154874 3772
rect 155033 3770 155099 3773
rect 154868 3768 155099 3770
rect 154868 3712 155038 3768
rect 155094 3712 155099 3768
rect 154868 3710 155099 3712
rect 154868 3708 154874 3710
rect 155033 3707 155099 3710
rect 118785 3634 118851 3637
rect 132953 3634 133019 3637
rect 118785 3632 133019 3634
rect 118785 3576 118790 3632
rect 118846 3576 132958 3632
rect 133014 3576 133019 3632
rect 118785 3574 133019 3576
rect 118785 3571 118851 3574
rect 132953 3571 133019 3574
rect 137921 3634 137987 3637
rect 143625 3634 143691 3637
rect 137921 3632 143691 3634
rect 137921 3576 137926 3632
rect 137982 3576 143630 3632
rect 143686 3576 143691 3632
rect 137921 3574 143691 3576
rect 137921 3571 137987 3574
rect 143625 3571 143691 3574
rect 146937 3634 147003 3637
rect 147489 3634 147555 3637
rect 146937 3632 147555 3634
rect 146937 3576 146942 3632
rect 146998 3576 147494 3632
rect 147550 3576 147555 3632
rect 146937 3574 147555 3576
rect 146937 3571 147003 3574
rect 147489 3571 147555 3574
rect 147673 3634 147739 3637
rect 149697 3634 149763 3637
rect 147673 3632 149763 3634
rect 147673 3576 147678 3632
rect 147734 3576 149702 3632
rect 149758 3576 149763 3632
rect 147673 3574 149763 3576
rect 147673 3571 147739 3574
rect 149697 3571 149763 3574
rect 74809 3498 74875 3501
rect 130745 3498 130811 3501
rect 74809 3496 130811 3498
rect 74809 3440 74814 3496
rect 74870 3440 130750 3496
rect 130806 3440 130811 3496
rect 74809 3438 130811 3440
rect 74809 3435 74875 3438
rect 130745 3435 130811 3438
rect 131113 3498 131179 3501
rect 148225 3498 148291 3501
rect 131113 3496 148291 3498
rect 131113 3440 131118 3496
rect 131174 3440 148230 3496
rect 148286 3440 148291 3496
rect 131113 3438 148291 3440
rect 131113 3435 131179 3438
rect 148225 3435 148291 3438
rect 148869 3498 148935 3501
rect 150065 3498 150131 3501
rect 148869 3496 150131 3498
rect 148869 3440 148874 3496
rect 148930 3440 150070 3496
rect 150126 3440 150131 3496
rect 148869 3438 150131 3440
rect 148869 3435 148935 3438
rect 150065 3435 150131 3438
rect 151537 3498 151603 3501
rect 151670 3498 151676 3500
rect 151537 3496 151676 3498
rect 151537 3440 151542 3496
rect 151598 3440 151676 3496
rect 151537 3438 151676 3440
rect 151537 3435 151603 3438
rect 151670 3436 151676 3438
rect 151740 3436 151746 3500
rect 152457 3498 152523 3501
rect 152641 3498 152707 3501
rect 154481 3498 154547 3501
rect 152457 3496 154547 3498
rect 152457 3440 152462 3496
rect 152518 3440 152646 3496
rect 152702 3440 154486 3496
rect 154542 3440 154547 3496
rect 152457 3438 154547 3440
rect 152457 3435 152523 3438
rect 152641 3435 152707 3438
rect 154481 3435 154547 3438
rect 154665 3498 154731 3501
rect 155125 3498 155191 3501
rect 154665 3496 155191 3498
rect 154665 3440 154670 3496
rect 154726 3440 155130 3496
rect 155186 3440 155191 3496
rect 154665 3438 155191 3440
rect 154665 3435 154731 3438
rect 155125 3435 155191 3438
rect 49601 3362 49667 3365
rect 53557 3362 53623 3365
rect 49601 3360 53623 3362
rect 49601 3304 49606 3360
rect 49662 3304 53562 3360
rect 53618 3304 53623 3360
rect 49601 3302 53623 3304
rect 49601 3299 49667 3302
rect 53557 3299 53623 3302
rect 147305 3362 147371 3365
rect 147857 3362 147923 3365
rect 147305 3360 147923 3362
rect 147305 3304 147310 3360
rect 147366 3304 147862 3360
rect 147918 3304 147923 3360
rect 147305 3302 147923 3304
rect 147305 3299 147371 3302
rect 147857 3299 147923 3302
rect 148685 3362 148751 3365
rect 150433 3362 150499 3365
rect 148685 3360 150499 3362
rect 148685 3304 148690 3360
rect 148746 3304 150438 3360
rect 150494 3304 150499 3360
rect 148685 3302 150499 3304
rect 148685 3299 148751 3302
rect 150433 3299 150499 3302
rect 151077 3362 151143 3365
rect 153469 3362 153535 3365
rect 151077 3360 153535 3362
rect 151077 3304 151082 3360
rect 151138 3304 153474 3360
rect 153530 3304 153535 3360
rect 151077 3302 153535 3304
rect 151077 3299 151143 3302
rect 153469 3299 153535 3302
rect 154297 3362 154363 3365
rect 157609 3362 157675 3365
rect 154297 3360 157675 3362
rect 154297 3304 154302 3360
rect 154358 3304 157614 3360
rect 157670 3304 157675 3360
rect 154297 3302 157675 3304
rect 154297 3299 154363 3302
rect 157609 3299 157675 3302
rect 40390 3296 40706 3297
rect 40390 3232 40396 3296
rect 40460 3232 40476 3296
rect 40540 3232 40556 3296
rect 40620 3232 40636 3296
rect 40700 3232 40706 3296
rect 40390 3231 40706 3232
rect 79835 3296 80151 3297
rect 79835 3232 79841 3296
rect 79905 3232 79921 3296
rect 79985 3232 80001 3296
rect 80065 3232 80081 3296
rect 80145 3232 80151 3296
rect 79835 3231 80151 3232
rect 119280 3296 119596 3297
rect 119280 3232 119286 3296
rect 119350 3232 119366 3296
rect 119430 3232 119446 3296
rect 119510 3232 119526 3296
rect 119590 3232 119596 3296
rect 119280 3231 119596 3232
rect 158725 3296 159041 3297
rect 158725 3232 158731 3296
rect 158795 3232 158811 3296
rect 158875 3232 158891 3296
rect 158955 3232 158971 3296
rect 159035 3232 159041 3296
rect 158725 3231 159041 3232
rect 134149 3226 134215 3229
rect 153285 3226 153351 3229
rect 134149 3224 153351 3226
rect 134149 3168 134154 3224
rect 134210 3168 153290 3224
rect 153346 3168 153351 3224
rect 134149 3166 153351 3168
rect 134149 3163 134215 3166
rect 153285 3163 153351 3166
rect 20529 3090 20595 3093
rect 24761 3090 24827 3093
rect 20529 3088 24827 3090
rect 20529 3032 20534 3088
rect 20590 3032 24766 3088
rect 24822 3032 24827 3088
rect 20529 3030 24827 3032
rect 20529 3027 20595 3030
rect 24761 3027 24827 3030
rect 93485 3090 93551 3093
rect 123385 3090 123451 3093
rect 137737 3090 137803 3093
rect 93485 3088 137803 3090
rect 93485 3032 93490 3088
rect 93546 3032 123390 3088
rect 123446 3032 137742 3088
rect 137798 3032 137803 3088
rect 93485 3030 137803 3032
rect 93485 3027 93551 3030
rect 123385 3027 123451 3030
rect 137737 3027 137803 3030
rect 145465 3090 145531 3093
rect 147857 3090 147923 3093
rect 145465 3088 147923 3090
rect 145465 3032 145470 3088
rect 145526 3032 147862 3088
rect 147918 3032 147923 3088
rect 145465 3030 147923 3032
rect 145465 3027 145531 3030
rect 147857 3027 147923 3030
rect 148777 3090 148843 3093
rect 158069 3090 158135 3093
rect 148777 3088 158135 3090
rect 148777 3032 148782 3088
rect 148838 3032 158074 3088
rect 158130 3032 158135 3088
rect 148777 3030 158135 3032
rect 148777 3027 148843 3030
rect 158069 3027 158135 3030
rect 96705 2954 96771 2957
rect 130193 2954 130259 2957
rect 96705 2952 130259 2954
rect 96705 2896 96710 2952
rect 96766 2896 130198 2952
rect 130254 2896 130259 2952
rect 96705 2894 130259 2896
rect 96705 2891 96771 2894
rect 130193 2891 130259 2894
rect 135989 2954 136055 2957
rect 148501 2954 148567 2957
rect 135989 2952 148567 2954
rect 135989 2896 135994 2952
rect 136050 2896 148506 2952
rect 148562 2896 148567 2952
rect 135989 2894 148567 2896
rect 135989 2891 136055 2894
rect 148501 2891 148567 2894
rect 151813 2954 151879 2957
rect 154021 2954 154087 2957
rect 151813 2952 154087 2954
rect 151813 2896 151818 2952
rect 151874 2896 154026 2952
rect 154082 2896 154087 2952
rect 151813 2894 154087 2896
rect 151813 2891 151879 2894
rect 154021 2891 154087 2894
rect 117589 2818 117655 2821
rect 120165 2818 120231 2821
rect 117589 2816 120231 2818
rect 117589 2760 117594 2816
rect 117650 2760 120170 2816
rect 120226 2760 120231 2816
rect 117589 2758 120231 2760
rect 117589 2755 117655 2758
rect 120165 2755 120231 2758
rect 148685 2818 148751 2821
rect 155953 2818 156019 2821
rect 148685 2816 156019 2818
rect 148685 2760 148690 2816
rect 148746 2760 155958 2816
rect 156014 2760 156019 2816
rect 148685 2758 156019 2760
rect 148685 2755 148751 2758
rect 155953 2755 156019 2758
rect 20668 2752 20984 2753
rect 20668 2688 20674 2752
rect 20738 2688 20754 2752
rect 20818 2688 20834 2752
rect 20898 2688 20914 2752
rect 20978 2688 20984 2752
rect 20668 2687 20984 2688
rect 60113 2752 60429 2753
rect 60113 2688 60119 2752
rect 60183 2688 60199 2752
rect 60263 2688 60279 2752
rect 60343 2688 60359 2752
rect 60423 2688 60429 2752
rect 60113 2687 60429 2688
rect 99558 2752 99874 2753
rect 99558 2688 99564 2752
rect 99628 2688 99644 2752
rect 99708 2688 99724 2752
rect 99788 2688 99804 2752
rect 99868 2688 99874 2752
rect 99558 2687 99874 2688
rect 139003 2752 139319 2753
rect 139003 2688 139009 2752
rect 139073 2688 139089 2752
rect 139153 2688 139169 2752
rect 139233 2688 139249 2752
rect 139313 2688 139319 2752
rect 139003 2687 139319 2688
rect 118509 2682 118575 2685
rect 123017 2682 123083 2685
rect 118509 2680 123083 2682
rect 118509 2624 118514 2680
rect 118570 2624 123022 2680
rect 123078 2624 123083 2680
rect 118509 2622 123083 2624
rect 118509 2619 118575 2622
rect 123017 2619 123083 2622
rect 135069 2682 135135 2685
rect 136633 2682 136699 2685
rect 135069 2680 136699 2682
rect 135069 2624 135074 2680
rect 135130 2624 136638 2680
rect 136694 2624 136699 2680
rect 135069 2622 136699 2624
rect 135069 2619 135135 2622
rect 136633 2619 136699 2622
rect 141049 2682 141115 2685
rect 154297 2682 154363 2685
rect 141049 2680 154363 2682
rect 141049 2624 141054 2680
rect 141110 2624 154302 2680
rect 154358 2624 154363 2680
rect 141049 2622 154363 2624
rect 141049 2619 141115 2622
rect 154297 2619 154363 2622
rect 119981 2546 120047 2549
rect 129549 2546 129615 2549
rect 119981 2544 129615 2546
rect 119981 2488 119986 2544
rect 120042 2488 129554 2544
rect 129610 2488 129615 2544
rect 119981 2486 129615 2488
rect 119981 2483 120047 2486
rect 129549 2483 129615 2486
rect 131297 2546 131363 2549
rect 143717 2546 143783 2549
rect 131297 2544 143783 2546
rect 131297 2488 131302 2544
rect 131358 2488 143722 2544
rect 143778 2488 143783 2544
rect 131297 2486 143783 2488
rect 131297 2483 131363 2486
rect 143717 2483 143783 2486
rect 149605 2546 149671 2549
rect 152365 2546 152431 2549
rect 149605 2544 152431 2546
rect 149605 2488 149610 2544
rect 149666 2488 152370 2544
rect 152426 2488 152431 2544
rect 149605 2486 152431 2488
rect 149605 2483 149671 2486
rect 152365 2483 152431 2486
rect 95601 2410 95667 2413
rect 117405 2410 117471 2413
rect 138013 2410 138079 2413
rect 95601 2408 138079 2410
rect 95601 2352 95606 2408
rect 95662 2352 117410 2408
rect 117466 2352 138018 2408
rect 138074 2352 138079 2408
rect 95601 2350 138079 2352
rect 95601 2347 95667 2350
rect 117405 2347 117471 2350
rect 138013 2347 138079 2350
rect 140589 2410 140655 2413
rect 153653 2410 153719 2413
rect 140589 2408 153719 2410
rect 140589 2352 140594 2408
rect 140650 2352 153658 2408
rect 153714 2352 153719 2408
rect 140589 2350 153719 2352
rect 140589 2347 140655 2350
rect 153653 2347 153719 2350
rect 134057 2274 134123 2277
rect 141049 2274 141115 2277
rect 134057 2272 141115 2274
rect 134057 2216 134062 2272
rect 134118 2216 141054 2272
rect 141110 2216 141115 2272
rect 134057 2214 141115 2216
rect 134057 2211 134123 2214
rect 141049 2211 141115 2214
rect 145925 2274 145991 2277
rect 158161 2274 158227 2277
rect 145925 2272 158227 2274
rect 145925 2216 145930 2272
rect 145986 2216 158166 2272
rect 158222 2216 158227 2272
rect 145925 2214 158227 2216
rect 145925 2211 145991 2214
rect 158161 2211 158227 2214
rect 40390 2208 40706 2209
rect 40390 2144 40396 2208
rect 40460 2144 40476 2208
rect 40540 2144 40556 2208
rect 40620 2144 40636 2208
rect 40700 2144 40706 2208
rect 40390 2143 40706 2144
rect 79835 2208 80151 2209
rect 79835 2144 79841 2208
rect 79905 2144 79921 2208
rect 79985 2144 80001 2208
rect 80065 2144 80081 2208
rect 80145 2144 80151 2208
rect 79835 2143 80151 2144
rect 119280 2208 119596 2209
rect 119280 2144 119286 2208
rect 119350 2144 119366 2208
rect 119430 2144 119446 2208
rect 119510 2144 119526 2208
rect 119590 2144 119596 2208
rect 119280 2143 119596 2144
rect 158725 2208 159041 2209
rect 158725 2144 158731 2208
rect 158795 2144 158811 2208
rect 158875 2144 158891 2208
rect 158955 2144 158971 2208
rect 159035 2144 159041 2208
rect 158725 2143 159041 2144
rect 131062 2076 131068 2140
rect 131132 2138 131138 2140
rect 149605 2138 149671 2141
rect 131132 2136 149671 2138
rect 131132 2080 149610 2136
rect 149666 2080 149671 2136
rect 131132 2078 149671 2080
rect 131132 2076 131138 2078
rect 149605 2075 149671 2078
rect 150341 2138 150407 2141
rect 157793 2138 157859 2141
rect 150341 2136 157859 2138
rect 150341 2080 150346 2136
rect 150402 2080 157798 2136
rect 157854 2080 157859 2136
rect 150341 2078 157859 2080
rect 150341 2075 150407 2078
rect 157793 2075 157859 2078
rect 0 2002 800 2032
rect 1669 2002 1735 2005
rect 0 2000 1735 2002
rect 0 1944 1674 2000
rect 1730 1944 1735 2000
rect 0 1942 1735 1944
rect 0 1912 800 1942
rect 1669 1939 1735 1942
rect 108297 2002 108363 2005
rect 145005 2002 145071 2005
rect 108297 2000 145071 2002
rect 108297 1944 108302 2000
rect 108358 1944 145010 2000
rect 145066 1944 145071 2000
rect 108297 1942 145071 1944
rect 108297 1939 108363 1942
rect 145005 1939 145071 1942
rect 148133 2002 148199 2005
rect 155861 2002 155927 2005
rect 148133 2000 155927 2002
rect 148133 1944 148138 2000
rect 148194 1944 155866 2000
rect 155922 1944 155927 2000
rect 148133 1942 155927 1944
rect 148133 1939 148199 1942
rect 155861 1939 155927 1942
rect 143717 1866 143783 1869
rect 153326 1866 153332 1868
rect 143717 1864 153332 1866
rect 143717 1808 143722 1864
rect 143778 1808 153332 1864
rect 143717 1806 153332 1808
rect 143717 1803 143783 1806
rect 153326 1804 153332 1806
rect 153396 1804 153402 1868
rect 114277 1730 114343 1733
rect 149237 1730 149303 1733
rect 114277 1728 149303 1730
rect 114277 1672 114282 1728
rect 114338 1672 149242 1728
rect 149298 1672 149303 1728
rect 114277 1670 149303 1672
rect 114277 1667 114343 1670
rect 149237 1667 149303 1670
rect 123201 1322 123267 1325
rect 155902 1322 155908 1324
rect 123201 1320 155908 1322
rect 123201 1264 123206 1320
rect 123262 1264 155908 1320
rect 123201 1262 155908 1264
rect 123201 1259 123267 1262
rect 155902 1260 155908 1262
rect 155972 1260 155978 1324
rect 124438 1124 124444 1188
rect 124508 1186 124514 1188
rect 153745 1186 153811 1189
rect 124508 1184 153811 1186
rect 124508 1128 153750 1184
rect 153806 1128 153811 1184
rect 124508 1126 153811 1128
rect 124508 1124 124514 1126
rect 153745 1123 153811 1126
rect 145741 1050 145807 1053
rect 156413 1050 156479 1053
rect 145741 1048 156479 1050
rect 145741 992 145746 1048
rect 145802 992 156418 1048
rect 156474 992 156479 1048
rect 145741 990 156479 992
rect 145741 987 145807 990
rect 156413 987 156479 990
<< via3 >>
rect 150756 14452 150820 14516
rect 156828 14180 156892 14244
rect 155724 14044 155788 14108
rect 155172 13908 155236 13972
rect 20674 13628 20738 13632
rect 20674 13572 20678 13628
rect 20678 13572 20734 13628
rect 20734 13572 20738 13628
rect 20674 13568 20738 13572
rect 20754 13628 20818 13632
rect 20754 13572 20758 13628
rect 20758 13572 20814 13628
rect 20814 13572 20818 13628
rect 20754 13568 20818 13572
rect 20834 13628 20898 13632
rect 20834 13572 20838 13628
rect 20838 13572 20894 13628
rect 20894 13572 20898 13628
rect 20834 13568 20898 13572
rect 20914 13628 20978 13632
rect 20914 13572 20918 13628
rect 20918 13572 20974 13628
rect 20974 13572 20978 13628
rect 20914 13568 20978 13572
rect 60119 13628 60183 13632
rect 60119 13572 60123 13628
rect 60123 13572 60179 13628
rect 60179 13572 60183 13628
rect 60119 13568 60183 13572
rect 60199 13628 60263 13632
rect 60199 13572 60203 13628
rect 60203 13572 60259 13628
rect 60259 13572 60263 13628
rect 60199 13568 60263 13572
rect 60279 13628 60343 13632
rect 60279 13572 60283 13628
rect 60283 13572 60339 13628
rect 60339 13572 60343 13628
rect 60279 13568 60343 13572
rect 60359 13628 60423 13632
rect 60359 13572 60363 13628
rect 60363 13572 60419 13628
rect 60419 13572 60423 13628
rect 60359 13568 60423 13572
rect 99564 13628 99628 13632
rect 99564 13572 99568 13628
rect 99568 13572 99624 13628
rect 99624 13572 99628 13628
rect 99564 13568 99628 13572
rect 99644 13628 99708 13632
rect 99644 13572 99648 13628
rect 99648 13572 99704 13628
rect 99704 13572 99708 13628
rect 99644 13568 99708 13572
rect 99724 13628 99788 13632
rect 99724 13572 99728 13628
rect 99728 13572 99784 13628
rect 99784 13572 99788 13628
rect 99724 13568 99788 13572
rect 99804 13628 99868 13632
rect 99804 13572 99808 13628
rect 99808 13572 99864 13628
rect 99864 13572 99868 13628
rect 99804 13568 99868 13572
rect 139009 13628 139073 13632
rect 139009 13572 139013 13628
rect 139013 13572 139069 13628
rect 139069 13572 139073 13628
rect 139009 13568 139073 13572
rect 139089 13628 139153 13632
rect 139089 13572 139093 13628
rect 139093 13572 139149 13628
rect 139149 13572 139153 13628
rect 139089 13568 139153 13572
rect 139169 13628 139233 13632
rect 139169 13572 139173 13628
rect 139173 13572 139229 13628
rect 139229 13572 139233 13628
rect 139169 13568 139233 13572
rect 139249 13628 139313 13632
rect 139249 13572 139253 13628
rect 139253 13572 139309 13628
rect 139309 13572 139313 13628
rect 139249 13568 139313 13572
rect 40396 13084 40460 13088
rect 40396 13028 40400 13084
rect 40400 13028 40456 13084
rect 40456 13028 40460 13084
rect 40396 13024 40460 13028
rect 40476 13084 40540 13088
rect 40476 13028 40480 13084
rect 40480 13028 40536 13084
rect 40536 13028 40540 13084
rect 40476 13024 40540 13028
rect 40556 13084 40620 13088
rect 40556 13028 40560 13084
rect 40560 13028 40616 13084
rect 40616 13028 40620 13084
rect 40556 13024 40620 13028
rect 40636 13084 40700 13088
rect 40636 13028 40640 13084
rect 40640 13028 40696 13084
rect 40696 13028 40700 13084
rect 40636 13024 40700 13028
rect 79841 13084 79905 13088
rect 79841 13028 79845 13084
rect 79845 13028 79901 13084
rect 79901 13028 79905 13084
rect 79841 13024 79905 13028
rect 79921 13084 79985 13088
rect 79921 13028 79925 13084
rect 79925 13028 79981 13084
rect 79981 13028 79985 13084
rect 79921 13024 79985 13028
rect 80001 13084 80065 13088
rect 80001 13028 80005 13084
rect 80005 13028 80061 13084
rect 80061 13028 80065 13084
rect 80001 13024 80065 13028
rect 80081 13084 80145 13088
rect 80081 13028 80085 13084
rect 80085 13028 80141 13084
rect 80141 13028 80145 13084
rect 80081 13024 80145 13028
rect 119286 13084 119350 13088
rect 119286 13028 119290 13084
rect 119290 13028 119346 13084
rect 119346 13028 119350 13084
rect 119286 13024 119350 13028
rect 119366 13084 119430 13088
rect 119366 13028 119370 13084
rect 119370 13028 119426 13084
rect 119426 13028 119430 13084
rect 119366 13024 119430 13028
rect 119446 13084 119510 13088
rect 119446 13028 119450 13084
rect 119450 13028 119506 13084
rect 119506 13028 119510 13084
rect 119446 13024 119510 13028
rect 119526 13084 119590 13088
rect 119526 13028 119530 13084
rect 119530 13028 119586 13084
rect 119586 13028 119590 13084
rect 119526 13024 119590 13028
rect 158731 13084 158795 13088
rect 158731 13028 158735 13084
rect 158735 13028 158791 13084
rect 158791 13028 158795 13084
rect 158731 13024 158795 13028
rect 158811 13084 158875 13088
rect 158811 13028 158815 13084
rect 158815 13028 158871 13084
rect 158871 13028 158875 13084
rect 158811 13024 158875 13028
rect 158891 13084 158955 13088
rect 158891 13028 158895 13084
rect 158895 13028 158951 13084
rect 158951 13028 158955 13084
rect 158891 13024 158955 13028
rect 158971 13084 159035 13088
rect 158971 13028 158975 13084
rect 158975 13028 159031 13084
rect 159031 13028 159035 13084
rect 158971 13024 159035 13028
rect 149652 12956 149716 13020
rect 20674 12540 20738 12544
rect 20674 12484 20678 12540
rect 20678 12484 20734 12540
rect 20734 12484 20738 12540
rect 20674 12480 20738 12484
rect 20754 12540 20818 12544
rect 20754 12484 20758 12540
rect 20758 12484 20814 12540
rect 20814 12484 20818 12540
rect 20754 12480 20818 12484
rect 20834 12540 20898 12544
rect 20834 12484 20838 12540
rect 20838 12484 20894 12540
rect 20894 12484 20898 12540
rect 20834 12480 20898 12484
rect 20914 12540 20978 12544
rect 20914 12484 20918 12540
rect 20918 12484 20974 12540
rect 20974 12484 20978 12540
rect 20914 12480 20978 12484
rect 60119 12540 60183 12544
rect 60119 12484 60123 12540
rect 60123 12484 60179 12540
rect 60179 12484 60183 12540
rect 60119 12480 60183 12484
rect 60199 12540 60263 12544
rect 60199 12484 60203 12540
rect 60203 12484 60259 12540
rect 60259 12484 60263 12540
rect 60199 12480 60263 12484
rect 60279 12540 60343 12544
rect 60279 12484 60283 12540
rect 60283 12484 60339 12540
rect 60339 12484 60343 12540
rect 60279 12480 60343 12484
rect 60359 12540 60423 12544
rect 60359 12484 60363 12540
rect 60363 12484 60419 12540
rect 60419 12484 60423 12540
rect 60359 12480 60423 12484
rect 99564 12540 99628 12544
rect 99564 12484 99568 12540
rect 99568 12484 99624 12540
rect 99624 12484 99628 12540
rect 99564 12480 99628 12484
rect 99644 12540 99708 12544
rect 99644 12484 99648 12540
rect 99648 12484 99704 12540
rect 99704 12484 99708 12540
rect 99644 12480 99708 12484
rect 99724 12540 99788 12544
rect 99724 12484 99728 12540
rect 99728 12484 99784 12540
rect 99784 12484 99788 12540
rect 99724 12480 99788 12484
rect 99804 12540 99868 12544
rect 99804 12484 99808 12540
rect 99808 12484 99864 12540
rect 99864 12484 99868 12540
rect 99804 12480 99868 12484
rect 139009 12540 139073 12544
rect 139009 12484 139013 12540
rect 139013 12484 139069 12540
rect 139069 12484 139073 12540
rect 139009 12480 139073 12484
rect 139089 12540 139153 12544
rect 139089 12484 139093 12540
rect 139093 12484 139149 12540
rect 139149 12484 139153 12540
rect 139089 12480 139153 12484
rect 139169 12540 139233 12544
rect 139169 12484 139173 12540
rect 139173 12484 139229 12540
rect 139229 12484 139233 12540
rect 139169 12480 139233 12484
rect 139249 12540 139313 12544
rect 139249 12484 139253 12540
rect 139253 12484 139309 12540
rect 139309 12484 139313 12540
rect 139249 12480 139313 12484
rect 127204 12004 127268 12068
rect 40396 11996 40460 12000
rect 40396 11940 40400 11996
rect 40400 11940 40456 11996
rect 40456 11940 40460 11996
rect 40396 11936 40460 11940
rect 40476 11996 40540 12000
rect 40476 11940 40480 11996
rect 40480 11940 40536 11996
rect 40536 11940 40540 11996
rect 40476 11936 40540 11940
rect 40556 11996 40620 12000
rect 40556 11940 40560 11996
rect 40560 11940 40616 11996
rect 40616 11940 40620 11996
rect 40556 11936 40620 11940
rect 40636 11996 40700 12000
rect 40636 11940 40640 11996
rect 40640 11940 40696 11996
rect 40696 11940 40700 11996
rect 40636 11936 40700 11940
rect 79841 11996 79905 12000
rect 79841 11940 79845 11996
rect 79845 11940 79901 11996
rect 79901 11940 79905 11996
rect 79841 11936 79905 11940
rect 79921 11996 79985 12000
rect 79921 11940 79925 11996
rect 79925 11940 79981 11996
rect 79981 11940 79985 11996
rect 79921 11936 79985 11940
rect 80001 11996 80065 12000
rect 80001 11940 80005 11996
rect 80005 11940 80061 11996
rect 80061 11940 80065 11996
rect 80001 11936 80065 11940
rect 80081 11996 80145 12000
rect 80081 11940 80085 11996
rect 80085 11940 80141 11996
rect 80141 11940 80145 11996
rect 80081 11936 80145 11940
rect 119286 11996 119350 12000
rect 119286 11940 119290 11996
rect 119290 11940 119346 11996
rect 119346 11940 119350 11996
rect 119286 11936 119350 11940
rect 119366 11996 119430 12000
rect 119366 11940 119370 11996
rect 119370 11940 119426 11996
rect 119426 11940 119430 11996
rect 119366 11936 119430 11940
rect 119446 11996 119510 12000
rect 119446 11940 119450 11996
rect 119450 11940 119506 11996
rect 119506 11940 119510 11996
rect 119446 11936 119510 11940
rect 119526 11996 119590 12000
rect 119526 11940 119530 11996
rect 119530 11940 119586 11996
rect 119586 11940 119590 11996
rect 119526 11936 119590 11940
rect 131068 11868 131132 11932
rect 158731 11996 158795 12000
rect 158731 11940 158735 11996
rect 158735 11940 158791 11996
rect 158791 11940 158795 11996
rect 158731 11936 158795 11940
rect 158811 11996 158875 12000
rect 158811 11940 158815 11996
rect 158815 11940 158871 11996
rect 158871 11940 158875 11996
rect 158811 11936 158875 11940
rect 158891 11996 158955 12000
rect 158891 11940 158895 11996
rect 158895 11940 158951 11996
rect 158951 11940 158955 11996
rect 158891 11936 158955 11940
rect 158971 11996 159035 12000
rect 158971 11940 158975 11996
rect 158975 11940 159031 11996
rect 159031 11940 159035 11996
rect 158971 11936 159035 11940
rect 147996 11868 148060 11932
rect 133460 11732 133524 11796
rect 20674 11452 20738 11456
rect 20674 11396 20678 11452
rect 20678 11396 20734 11452
rect 20734 11396 20738 11452
rect 20674 11392 20738 11396
rect 20754 11452 20818 11456
rect 20754 11396 20758 11452
rect 20758 11396 20814 11452
rect 20814 11396 20818 11452
rect 20754 11392 20818 11396
rect 20834 11452 20898 11456
rect 20834 11396 20838 11452
rect 20838 11396 20894 11452
rect 20894 11396 20898 11452
rect 20834 11392 20898 11396
rect 20914 11452 20978 11456
rect 20914 11396 20918 11452
rect 20918 11396 20974 11452
rect 20974 11396 20978 11452
rect 20914 11392 20978 11396
rect 60119 11452 60183 11456
rect 60119 11396 60123 11452
rect 60123 11396 60179 11452
rect 60179 11396 60183 11452
rect 60119 11392 60183 11396
rect 60199 11452 60263 11456
rect 60199 11396 60203 11452
rect 60203 11396 60259 11452
rect 60259 11396 60263 11452
rect 60199 11392 60263 11396
rect 60279 11452 60343 11456
rect 60279 11396 60283 11452
rect 60283 11396 60339 11452
rect 60339 11396 60343 11452
rect 60279 11392 60343 11396
rect 60359 11452 60423 11456
rect 60359 11396 60363 11452
rect 60363 11396 60419 11452
rect 60419 11396 60423 11452
rect 60359 11392 60423 11396
rect 99564 11452 99628 11456
rect 99564 11396 99568 11452
rect 99568 11396 99624 11452
rect 99624 11396 99628 11452
rect 99564 11392 99628 11396
rect 99644 11452 99708 11456
rect 99644 11396 99648 11452
rect 99648 11396 99704 11452
rect 99704 11396 99708 11452
rect 99644 11392 99708 11396
rect 99724 11452 99788 11456
rect 99724 11396 99728 11452
rect 99728 11396 99784 11452
rect 99784 11396 99788 11452
rect 99724 11392 99788 11396
rect 99804 11452 99868 11456
rect 99804 11396 99808 11452
rect 99808 11396 99864 11452
rect 99864 11396 99868 11452
rect 99804 11392 99868 11396
rect 139009 11452 139073 11456
rect 139009 11396 139013 11452
rect 139013 11396 139069 11452
rect 139069 11396 139073 11452
rect 139009 11392 139073 11396
rect 139089 11452 139153 11456
rect 139089 11396 139093 11452
rect 139093 11396 139149 11452
rect 139149 11396 139153 11452
rect 139089 11392 139153 11396
rect 139169 11452 139233 11456
rect 139169 11396 139173 11452
rect 139173 11396 139229 11452
rect 139229 11396 139233 11452
rect 139169 11392 139233 11396
rect 139249 11452 139313 11456
rect 139249 11396 139253 11452
rect 139253 11396 139309 11452
rect 139309 11396 139313 11452
rect 139249 11392 139313 11396
rect 147444 11052 147508 11116
rect 152780 11112 152844 11116
rect 152780 11056 152830 11112
rect 152830 11056 152844 11112
rect 152780 11052 152844 11056
rect 146340 10916 146404 10980
rect 40396 10908 40460 10912
rect 40396 10852 40400 10908
rect 40400 10852 40456 10908
rect 40456 10852 40460 10908
rect 40396 10848 40460 10852
rect 40476 10908 40540 10912
rect 40476 10852 40480 10908
rect 40480 10852 40536 10908
rect 40536 10852 40540 10908
rect 40476 10848 40540 10852
rect 40556 10908 40620 10912
rect 40556 10852 40560 10908
rect 40560 10852 40616 10908
rect 40616 10852 40620 10908
rect 40556 10848 40620 10852
rect 40636 10908 40700 10912
rect 40636 10852 40640 10908
rect 40640 10852 40696 10908
rect 40696 10852 40700 10908
rect 40636 10848 40700 10852
rect 79841 10908 79905 10912
rect 79841 10852 79845 10908
rect 79845 10852 79901 10908
rect 79901 10852 79905 10908
rect 79841 10848 79905 10852
rect 79921 10908 79985 10912
rect 79921 10852 79925 10908
rect 79925 10852 79981 10908
rect 79981 10852 79985 10908
rect 79921 10848 79985 10852
rect 80001 10908 80065 10912
rect 80001 10852 80005 10908
rect 80005 10852 80061 10908
rect 80061 10852 80065 10908
rect 80001 10848 80065 10852
rect 80081 10908 80145 10912
rect 80081 10852 80085 10908
rect 80085 10852 80141 10908
rect 80141 10852 80145 10908
rect 80081 10848 80145 10852
rect 119286 10908 119350 10912
rect 119286 10852 119290 10908
rect 119290 10852 119346 10908
rect 119346 10852 119350 10908
rect 119286 10848 119350 10852
rect 119366 10908 119430 10912
rect 119366 10852 119370 10908
rect 119370 10852 119426 10908
rect 119426 10852 119430 10908
rect 119366 10848 119430 10852
rect 119446 10908 119510 10912
rect 119446 10852 119450 10908
rect 119450 10852 119506 10908
rect 119506 10852 119510 10908
rect 119446 10848 119510 10852
rect 119526 10908 119590 10912
rect 119526 10852 119530 10908
rect 119530 10852 119586 10908
rect 119586 10852 119590 10908
rect 119526 10848 119590 10852
rect 158731 10908 158795 10912
rect 158731 10852 158735 10908
rect 158735 10852 158791 10908
rect 158791 10852 158795 10908
rect 158731 10848 158795 10852
rect 158811 10908 158875 10912
rect 158811 10852 158815 10908
rect 158815 10852 158871 10908
rect 158871 10852 158875 10908
rect 158811 10848 158875 10852
rect 158891 10908 158955 10912
rect 158891 10852 158895 10908
rect 158895 10852 158951 10908
rect 158951 10852 158955 10908
rect 158891 10848 158955 10852
rect 158971 10908 159035 10912
rect 158971 10852 158975 10908
rect 158975 10852 159031 10908
rect 159031 10852 159035 10908
rect 158971 10848 159035 10852
rect 20674 10364 20738 10368
rect 20674 10308 20678 10364
rect 20678 10308 20734 10364
rect 20734 10308 20738 10364
rect 20674 10304 20738 10308
rect 20754 10364 20818 10368
rect 20754 10308 20758 10364
rect 20758 10308 20814 10364
rect 20814 10308 20818 10364
rect 20754 10304 20818 10308
rect 20834 10364 20898 10368
rect 20834 10308 20838 10364
rect 20838 10308 20894 10364
rect 20894 10308 20898 10364
rect 20834 10304 20898 10308
rect 20914 10364 20978 10368
rect 20914 10308 20918 10364
rect 20918 10308 20974 10364
rect 20974 10308 20978 10364
rect 20914 10304 20978 10308
rect 60119 10364 60183 10368
rect 60119 10308 60123 10364
rect 60123 10308 60179 10364
rect 60179 10308 60183 10364
rect 60119 10304 60183 10308
rect 60199 10364 60263 10368
rect 60199 10308 60203 10364
rect 60203 10308 60259 10364
rect 60259 10308 60263 10364
rect 60199 10304 60263 10308
rect 60279 10364 60343 10368
rect 60279 10308 60283 10364
rect 60283 10308 60339 10364
rect 60339 10308 60343 10364
rect 60279 10304 60343 10308
rect 60359 10364 60423 10368
rect 60359 10308 60363 10364
rect 60363 10308 60419 10364
rect 60419 10308 60423 10364
rect 60359 10304 60423 10308
rect 99564 10364 99628 10368
rect 99564 10308 99568 10364
rect 99568 10308 99624 10364
rect 99624 10308 99628 10364
rect 99564 10304 99628 10308
rect 99644 10364 99708 10368
rect 99644 10308 99648 10364
rect 99648 10308 99704 10364
rect 99704 10308 99708 10364
rect 99644 10304 99708 10308
rect 99724 10364 99788 10368
rect 99724 10308 99728 10364
rect 99728 10308 99784 10364
rect 99784 10308 99788 10364
rect 99724 10304 99788 10308
rect 99804 10364 99868 10368
rect 99804 10308 99808 10364
rect 99808 10308 99864 10364
rect 99864 10308 99868 10364
rect 99804 10304 99868 10308
rect 139009 10364 139073 10368
rect 139009 10308 139013 10364
rect 139013 10308 139069 10364
rect 139069 10308 139073 10364
rect 139009 10304 139073 10308
rect 139089 10364 139153 10368
rect 139089 10308 139093 10364
rect 139093 10308 139149 10364
rect 139149 10308 139153 10364
rect 139089 10304 139153 10308
rect 139169 10364 139233 10368
rect 139169 10308 139173 10364
rect 139173 10308 139229 10364
rect 139229 10308 139233 10364
rect 139169 10304 139233 10308
rect 139249 10364 139313 10368
rect 139249 10308 139253 10364
rect 139253 10308 139309 10364
rect 139309 10308 139313 10364
rect 139249 10304 139313 10308
rect 150388 10236 150452 10300
rect 40396 9820 40460 9824
rect 40396 9764 40400 9820
rect 40400 9764 40456 9820
rect 40456 9764 40460 9820
rect 40396 9760 40460 9764
rect 40476 9820 40540 9824
rect 40476 9764 40480 9820
rect 40480 9764 40536 9820
rect 40536 9764 40540 9820
rect 40476 9760 40540 9764
rect 40556 9820 40620 9824
rect 40556 9764 40560 9820
rect 40560 9764 40616 9820
rect 40616 9764 40620 9820
rect 40556 9760 40620 9764
rect 40636 9820 40700 9824
rect 40636 9764 40640 9820
rect 40640 9764 40696 9820
rect 40696 9764 40700 9820
rect 40636 9760 40700 9764
rect 79841 9820 79905 9824
rect 79841 9764 79845 9820
rect 79845 9764 79901 9820
rect 79901 9764 79905 9820
rect 79841 9760 79905 9764
rect 79921 9820 79985 9824
rect 79921 9764 79925 9820
rect 79925 9764 79981 9820
rect 79981 9764 79985 9820
rect 79921 9760 79985 9764
rect 80001 9820 80065 9824
rect 80001 9764 80005 9820
rect 80005 9764 80061 9820
rect 80061 9764 80065 9820
rect 80001 9760 80065 9764
rect 80081 9820 80145 9824
rect 80081 9764 80085 9820
rect 80085 9764 80141 9820
rect 80141 9764 80145 9820
rect 80081 9760 80145 9764
rect 119286 9820 119350 9824
rect 119286 9764 119290 9820
rect 119290 9764 119346 9820
rect 119346 9764 119350 9820
rect 119286 9760 119350 9764
rect 119366 9820 119430 9824
rect 119366 9764 119370 9820
rect 119370 9764 119426 9820
rect 119426 9764 119430 9820
rect 119366 9760 119430 9764
rect 119446 9820 119510 9824
rect 119446 9764 119450 9820
rect 119450 9764 119506 9820
rect 119506 9764 119510 9820
rect 119446 9760 119510 9764
rect 119526 9820 119590 9824
rect 119526 9764 119530 9820
rect 119530 9764 119586 9820
rect 119586 9764 119590 9820
rect 119526 9760 119590 9764
rect 158731 9820 158795 9824
rect 158731 9764 158735 9820
rect 158735 9764 158791 9820
rect 158791 9764 158795 9820
rect 158731 9760 158795 9764
rect 158811 9820 158875 9824
rect 158811 9764 158815 9820
rect 158815 9764 158871 9820
rect 158871 9764 158875 9820
rect 158811 9760 158875 9764
rect 158891 9820 158955 9824
rect 158891 9764 158895 9820
rect 158895 9764 158951 9820
rect 158951 9764 158955 9820
rect 158891 9760 158955 9764
rect 158971 9820 159035 9824
rect 158971 9764 158975 9820
rect 158975 9764 159031 9820
rect 159031 9764 159035 9820
rect 158971 9760 159035 9764
rect 124444 9752 124508 9756
rect 124444 9696 124458 9752
rect 124458 9696 124508 9752
rect 124444 9692 124508 9696
rect 152596 9616 152660 9620
rect 152596 9560 152610 9616
rect 152610 9560 152660 9616
rect 152596 9556 152660 9560
rect 20674 9276 20738 9280
rect 20674 9220 20678 9276
rect 20678 9220 20734 9276
rect 20734 9220 20738 9276
rect 20674 9216 20738 9220
rect 20754 9276 20818 9280
rect 20754 9220 20758 9276
rect 20758 9220 20814 9276
rect 20814 9220 20818 9276
rect 20754 9216 20818 9220
rect 20834 9276 20898 9280
rect 20834 9220 20838 9276
rect 20838 9220 20894 9276
rect 20894 9220 20898 9276
rect 20834 9216 20898 9220
rect 20914 9276 20978 9280
rect 20914 9220 20918 9276
rect 20918 9220 20974 9276
rect 20974 9220 20978 9276
rect 20914 9216 20978 9220
rect 60119 9276 60183 9280
rect 60119 9220 60123 9276
rect 60123 9220 60179 9276
rect 60179 9220 60183 9276
rect 60119 9216 60183 9220
rect 60199 9276 60263 9280
rect 60199 9220 60203 9276
rect 60203 9220 60259 9276
rect 60259 9220 60263 9276
rect 60199 9216 60263 9220
rect 60279 9276 60343 9280
rect 60279 9220 60283 9276
rect 60283 9220 60339 9276
rect 60339 9220 60343 9276
rect 60279 9216 60343 9220
rect 60359 9276 60423 9280
rect 60359 9220 60363 9276
rect 60363 9220 60419 9276
rect 60419 9220 60423 9276
rect 60359 9216 60423 9220
rect 99564 9276 99628 9280
rect 99564 9220 99568 9276
rect 99568 9220 99624 9276
rect 99624 9220 99628 9276
rect 99564 9216 99628 9220
rect 99644 9276 99708 9280
rect 99644 9220 99648 9276
rect 99648 9220 99704 9276
rect 99704 9220 99708 9276
rect 99644 9216 99708 9220
rect 99724 9276 99788 9280
rect 99724 9220 99728 9276
rect 99728 9220 99784 9276
rect 99784 9220 99788 9276
rect 99724 9216 99788 9220
rect 99804 9276 99868 9280
rect 99804 9220 99808 9276
rect 99808 9220 99864 9276
rect 99864 9220 99868 9276
rect 99804 9216 99868 9220
rect 139009 9276 139073 9280
rect 139009 9220 139013 9276
rect 139013 9220 139069 9276
rect 139069 9220 139073 9276
rect 139009 9216 139073 9220
rect 139089 9276 139153 9280
rect 139089 9220 139093 9276
rect 139093 9220 139149 9276
rect 139149 9220 139153 9276
rect 139089 9216 139153 9220
rect 139169 9276 139233 9280
rect 139169 9220 139173 9276
rect 139173 9220 139229 9276
rect 139229 9220 139233 9276
rect 139169 9216 139233 9220
rect 139249 9276 139313 9280
rect 139249 9220 139253 9276
rect 139253 9220 139309 9276
rect 139309 9220 139313 9276
rect 139249 9216 139313 9220
rect 139716 8876 139780 8940
rect 148548 8876 148612 8940
rect 154804 8876 154868 8940
rect 127204 8740 127268 8804
rect 150388 8740 150452 8804
rect 40396 8732 40460 8736
rect 40396 8676 40400 8732
rect 40400 8676 40456 8732
rect 40456 8676 40460 8732
rect 40396 8672 40460 8676
rect 40476 8732 40540 8736
rect 40476 8676 40480 8732
rect 40480 8676 40536 8732
rect 40536 8676 40540 8732
rect 40476 8672 40540 8676
rect 40556 8732 40620 8736
rect 40556 8676 40560 8732
rect 40560 8676 40616 8732
rect 40616 8676 40620 8732
rect 40556 8672 40620 8676
rect 40636 8732 40700 8736
rect 40636 8676 40640 8732
rect 40640 8676 40696 8732
rect 40696 8676 40700 8732
rect 40636 8672 40700 8676
rect 79841 8732 79905 8736
rect 79841 8676 79845 8732
rect 79845 8676 79901 8732
rect 79901 8676 79905 8732
rect 79841 8672 79905 8676
rect 79921 8732 79985 8736
rect 79921 8676 79925 8732
rect 79925 8676 79981 8732
rect 79981 8676 79985 8732
rect 79921 8672 79985 8676
rect 80001 8732 80065 8736
rect 80001 8676 80005 8732
rect 80005 8676 80061 8732
rect 80061 8676 80065 8732
rect 80001 8672 80065 8676
rect 80081 8732 80145 8736
rect 80081 8676 80085 8732
rect 80085 8676 80141 8732
rect 80141 8676 80145 8732
rect 80081 8672 80145 8676
rect 119286 8732 119350 8736
rect 119286 8676 119290 8732
rect 119290 8676 119346 8732
rect 119346 8676 119350 8732
rect 119286 8672 119350 8676
rect 119366 8732 119430 8736
rect 119366 8676 119370 8732
rect 119370 8676 119426 8732
rect 119426 8676 119430 8732
rect 119366 8672 119430 8676
rect 119446 8732 119510 8736
rect 119446 8676 119450 8732
rect 119450 8676 119506 8732
rect 119506 8676 119510 8732
rect 119446 8672 119510 8676
rect 119526 8732 119590 8736
rect 119526 8676 119530 8732
rect 119530 8676 119586 8732
rect 119586 8676 119590 8732
rect 119526 8672 119590 8676
rect 158731 8732 158795 8736
rect 158731 8676 158735 8732
rect 158735 8676 158791 8732
rect 158791 8676 158795 8732
rect 158731 8672 158795 8676
rect 158811 8732 158875 8736
rect 158811 8676 158815 8732
rect 158815 8676 158871 8732
rect 158871 8676 158875 8732
rect 158811 8672 158875 8676
rect 158891 8732 158955 8736
rect 158891 8676 158895 8732
rect 158895 8676 158951 8732
rect 158951 8676 158955 8732
rect 158891 8672 158955 8676
rect 158971 8732 159035 8736
rect 158971 8676 158975 8732
rect 158975 8676 159031 8732
rect 159031 8676 159035 8732
rect 158971 8672 159035 8676
rect 147076 8604 147140 8668
rect 149652 8664 149716 8668
rect 149652 8608 149666 8664
rect 149666 8608 149716 8664
rect 149652 8604 149716 8608
rect 150204 8664 150268 8668
rect 150204 8608 150218 8664
rect 150218 8608 150268 8664
rect 150204 8604 150268 8608
rect 124260 8332 124324 8396
rect 153148 8332 153212 8396
rect 20674 8188 20738 8192
rect 20674 8132 20678 8188
rect 20678 8132 20734 8188
rect 20734 8132 20738 8188
rect 20674 8128 20738 8132
rect 20754 8188 20818 8192
rect 20754 8132 20758 8188
rect 20758 8132 20814 8188
rect 20814 8132 20818 8188
rect 20754 8128 20818 8132
rect 20834 8188 20898 8192
rect 20834 8132 20838 8188
rect 20838 8132 20894 8188
rect 20894 8132 20898 8188
rect 20834 8128 20898 8132
rect 20914 8188 20978 8192
rect 20914 8132 20918 8188
rect 20918 8132 20974 8188
rect 20974 8132 20978 8188
rect 20914 8128 20978 8132
rect 60119 8188 60183 8192
rect 60119 8132 60123 8188
rect 60123 8132 60179 8188
rect 60179 8132 60183 8188
rect 60119 8128 60183 8132
rect 60199 8188 60263 8192
rect 60199 8132 60203 8188
rect 60203 8132 60259 8188
rect 60259 8132 60263 8188
rect 60199 8128 60263 8132
rect 60279 8188 60343 8192
rect 60279 8132 60283 8188
rect 60283 8132 60339 8188
rect 60339 8132 60343 8188
rect 60279 8128 60343 8132
rect 60359 8188 60423 8192
rect 60359 8132 60363 8188
rect 60363 8132 60419 8188
rect 60419 8132 60423 8188
rect 60359 8128 60423 8132
rect 99564 8188 99628 8192
rect 99564 8132 99568 8188
rect 99568 8132 99624 8188
rect 99624 8132 99628 8188
rect 99564 8128 99628 8132
rect 99644 8188 99708 8192
rect 99644 8132 99648 8188
rect 99648 8132 99704 8188
rect 99704 8132 99708 8188
rect 99644 8128 99708 8132
rect 99724 8188 99788 8192
rect 99724 8132 99728 8188
rect 99728 8132 99784 8188
rect 99784 8132 99788 8188
rect 99724 8128 99788 8132
rect 99804 8188 99868 8192
rect 99804 8132 99808 8188
rect 99808 8132 99864 8188
rect 99864 8132 99868 8188
rect 99804 8128 99868 8132
rect 145052 8196 145116 8260
rect 139009 8188 139073 8192
rect 139009 8132 139013 8188
rect 139013 8132 139069 8188
rect 139069 8132 139073 8188
rect 139009 8128 139073 8132
rect 139089 8188 139153 8192
rect 139089 8132 139093 8188
rect 139093 8132 139149 8188
rect 139149 8132 139153 8188
rect 139089 8128 139153 8132
rect 139169 8188 139233 8192
rect 139169 8132 139173 8188
rect 139173 8132 139229 8188
rect 139229 8132 139233 8188
rect 139169 8128 139233 8132
rect 139249 8188 139313 8192
rect 139249 8132 139253 8188
rect 139253 8132 139309 8188
rect 139309 8132 139313 8188
rect 139249 8128 139313 8132
rect 146892 8060 146956 8124
rect 147260 8120 147324 8124
rect 147260 8064 147274 8120
rect 147274 8064 147324 8120
rect 147260 8060 147324 8064
rect 148916 8196 148980 8260
rect 150388 8196 150452 8260
rect 151676 8196 151740 8260
rect 154252 7788 154316 7852
rect 40396 7644 40460 7648
rect 40396 7588 40400 7644
rect 40400 7588 40456 7644
rect 40456 7588 40460 7644
rect 40396 7584 40460 7588
rect 40476 7644 40540 7648
rect 40476 7588 40480 7644
rect 40480 7588 40536 7644
rect 40536 7588 40540 7644
rect 40476 7584 40540 7588
rect 40556 7644 40620 7648
rect 40556 7588 40560 7644
rect 40560 7588 40616 7644
rect 40616 7588 40620 7644
rect 40556 7584 40620 7588
rect 40636 7644 40700 7648
rect 40636 7588 40640 7644
rect 40640 7588 40696 7644
rect 40696 7588 40700 7644
rect 40636 7584 40700 7588
rect 79841 7644 79905 7648
rect 79841 7588 79845 7644
rect 79845 7588 79901 7644
rect 79901 7588 79905 7644
rect 79841 7584 79905 7588
rect 79921 7644 79985 7648
rect 79921 7588 79925 7644
rect 79925 7588 79981 7644
rect 79981 7588 79985 7644
rect 79921 7584 79985 7588
rect 80001 7644 80065 7648
rect 80001 7588 80005 7644
rect 80005 7588 80061 7644
rect 80061 7588 80065 7644
rect 80001 7584 80065 7588
rect 80081 7644 80145 7648
rect 80081 7588 80085 7644
rect 80085 7588 80141 7644
rect 80141 7588 80145 7644
rect 80081 7584 80145 7588
rect 119286 7644 119350 7648
rect 119286 7588 119290 7644
rect 119290 7588 119346 7644
rect 119346 7588 119350 7644
rect 119286 7584 119350 7588
rect 119366 7644 119430 7648
rect 119366 7588 119370 7644
rect 119370 7588 119426 7644
rect 119426 7588 119430 7644
rect 119366 7584 119430 7588
rect 119446 7644 119510 7648
rect 119446 7588 119450 7644
rect 119450 7588 119506 7644
rect 119506 7588 119510 7644
rect 119446 7584 119510 7588
rect 119526 7644 119590 7648
rect 119526 7588 119530 7644
rect 119530 7588 119586 7644
rect 119586 7588 119590 7644
rect 119526 7584 119590 7588
rect 158731 7644 158795 7648
rect 158731 7588 158735 7644
rect 158735 7588 158791 7644
rect 158791 7588 158795 7644
rect 158731 7584 158795 7588
rect 158811 7644 158875 7648
rect 158811 7588 158815 7644
rect 158815 7588 158871 7644
rect 158871 7588 158875 7644
rect 158811 7584 158875 7588
rect 158891 7644 158955 7648
rect 158891 7588 158895 7644
rect 158895 7588 158951 7644
rect 158951 7588 158955 7644
rect 158891 7584 158955 7588
rect 158971 7644 159035 7648
rect 158971 7588 158975 7644
rect 158975 7588 159031 7644
rect 159031 7588 159035 7644
rect 158971 7584 159035 7588
rect 150388 7380 150452 7444
rect 150756 7576 150820 7580
rect 150756 7520 150806 7576
rect 150806 7520 150820 7576
rect 150756 7516 150820 7520
rect 20674 7100 20738 7104
rect 20674 7044 20678 7100
rect 20678 7044 20734 7100
rect 20734 7044 20738 7100
rect 20674 7040 20738 7044
rect 20754 7100 20818 7104
rect 20754 7044 20758 7100
rect 20758 7044 20814 7100
rect 20814 7044 20818 7100
rect 20754 7040 20818 7044
rect 20834 7100 20898 7104
rect 20834 7044 20838 7100
rect 20838 7044 20894 7100
rect 20894 7044 20898 7100
rect 20834 7040 20898 7044
rect 20914 7100 20978 7104
rect 20914 7044 20918 7100
rect 20918 7044 20974 7100
rect 20974 7044 20978 7100
rect 20914 7040 20978 7044
rect 60119 7100 60183 7104
rect 60119 7044 60123 7100
rect 60123 7044 60179 7100
rect 60179 7044 60183 7100
rect 60119 7040 60183 7044
rect 60199 7100 60263 7104
rect 60199 7044 60203 7100
rect 60203 7044 60259 7100
rect 60259 7044 60263 7100
rect 60199 7040 60263 7044
rect 60279 7100 60343 7104
rect 60279 7044 60283 7100
rect 60283 7044 60339 7100
rect 60339 7044 60343 7100
rect 60279 7040 60343 7044
rect 60359 7100 60423 7104
rect 60359 7044 60363 7100
rect 60363 7044 60419 7100
rect 60419 7044 60423 7100
rect 60359 7040 60423 7044
rect 99564 7100 99628 7104
rect 99564 7044 99568 7100
rect 99568 7044 99624 7100
rect 99624 7044 99628 7100
rect 99564 7040 99628 7044
rect 99644 7100 99708 7104
rect 99644 7044 99648 7100
rect 99648 7044 99704 7100
rect 99704 7044 99708 7100
rect 99644 7040 99708 7044
rect 99724 7100 99788 7104
rect 99724 7044 99728 7100
rect 99728 7044 99784 7100
rect 99784 7044 99788 7100
rect 99724 7040 99788 7044
rect 99804 7100 99868 7104
rect 99804 7044 99808 7100
rect 99808 7044 99864 7100
rect 99864 7044 99868 7100
rect 99804 7040 99868 7044
rect 131068 7108 131132 7172
rect 146892 7108 146956 7172
rect 147444 7108 147508 7172
rect 147812 7108 147876 7172
rect 139009 7100 139073 7104
rect 139009 7044 139013 7100
rect 139013 7044 139069 7100
rect 139069 7044 139073 7100
rect 139009 7040 139073 7044
rect 139089 7100 139153 7104
rect 139089 7044 139093 7100
rect 139093 7044 139149 7100
rect 139149 7044 139153 7100
rect 139089 7040 139153 7044
rect 139169 7100 139233 7104
rect 139169 7044 139173 7100
rect 139173 7044 139229 7100
rect 139229 7044 139233 7100
rect 139169 7040 139233 7044
rect 139249 7100 139313 7104
rect 139249 7044 139253 7100
rect 139253 7044 139309 7100
rect 139309 7044 139313 7100
rect 139249 7040 139313 7044
rect 145052 7032 145116 7036
rect 145052 6976 145066 7032
rect 145066 6976 145116 7032
rect 145052 6972 145116 6976
rect 153332 6972 153396 7036
rect 133460 6896 133524 6900
rect 133460 6840 133474 6896
rect 133474 6840 133524 6896
rect 133460 6836 133524 6840
rect 147812 6836 147876 6900
rect 127204 6564 127268 6628
rect 40396 6556 40460 6560
rect 40396 6500 40400 6556
rect 40400 6500 40456 6556
rect 40456 6500 40460 6556
rect 40396 6496 40460 6500
rect 40476 6556 40540 6560
rect 40476 6500 40480 6556
rect 40480 6500 40536 6556
rect 40536 6500 40540 6556
rect 40476 6496 40540 6500
rect 40556 6556 40620 6560
rect 40556 6500 40560 6556
rect 40560 6500 40616 6556
rect 40616 6500 40620 6556
rect 40556 6496 40620 6500
rect 40636 6556 40700 6560
rect 40636 6500 40640 6556
rect 40640 6500 40696 6556
rect 40696 6500 40700 6556
rect 40636 6496 40700 6500
rect 79841 6556 79905 6560
rect 79841 6500 79845 6556
rect 79845 6500 79901 6556
rect 79901 6500 79905 6556
rect 79841 6496 79905 6500
rect 79921 6556 79985 6560
rect 79921 6500 79925 6556
rect 79925 6500 79981 6556
rect 79981 6500 79985 6556
rect 79921 6496 79985 6500
rect 80001 6556 80065 6560
rect 80001 6500 80005 6556
rect 80005 6500 80061 6556
rect 80061 6500 80065 6556
rect 80001 6496 80065 6500
rect 80081 6556 80145 6560
rect 80081 6500 80085 6556
rect 80085 6500 80141 6556
rect 80141 6500 80145 6556
rect 80081 6496 80145 6500
rect 119286 6556 119350 6560
rect 119286 6500 119290 6556
rect 119290 6500 119346 6556
rect 119346 6500 119350 6556
rect 119286 6496 119350 6500
rect 119366 6556 119430 6560
rect 119366 6500 119370 6556
rect 119370 6500 119426 6556
rect 119426 6500 119430 6556
rect 119366 6496 119430 6500
rect 119446 6556 119510 6560
rect 119446 6500 119450 6556
rect 119450 6500 119506 6556
rect 119506 6500 119510 6556
rect 119446 6496 119510 6500
rect 119526 6556 119590 6560
rect 119526 6500 119530 6556
rect 119530 6500 119586 6556
rect 119586 6500 119590 6556
rect 119526 6496 119590 6500
rect 158731 6556 158795 6560
rect 158731 6500 158735 6556
rect 158735 6500 158791 6556
rect 158791 6500 158795 6556
rect 158731 6496 158795 6500
rect 158811 6556 158875 6560
rect 158811 6500 158815 6556
rect 158815 6500 158871 6556
rect 158871 6500 158875 6556
rect 158811 6496 158875 6500
rect 158891 6556 158955 6560
rect 158891 6500 158895 6556
rect 158895 6500 158951 6556
rect 158951 6500 158955 6556
rect 158891 6496 158955 6500
rect 158971 6556 159035 6560
rect 158971 6500 158975 6556
rect 158975 6500 159031 6556
rect 159031 6500 159035 6556
rect 158971 6496 159035 6500
rect 146340 6428 146404 6492
rect 139716 6292 139780 6356
rect 149284 6156 149348 6220
rect 20674 6012 20738 6016
rect 20674 5956 20678 6012
rect 20678 5956 20734 6012
rect 20734 5956 20738 6012
rect 20674 5952 20738 5956
rect 20754 6012 20818 6016
rect 20754 5956 20758 6012
rect 20758 5956 20814 6012
rect 20814 5956 20818 6012
rect 20754 5952 20818 5956
rect 20834 6012 20898 6016
rect 20834 5956 20838 6012
rect 20838 5956 20894 6012
rect 20894 5956 20898 6012
rect 20834 5952 20898 5956
rect 20914 6012 20978 6016
rect 20914 5956 20918 6012
rect 20918 5956 20974 6012
rect 20974 5956 20978 6012
rect 20914 5952 20978 5956
rect 60119 6012 60183 6016
rect 60119 5956 60123 6012
rect 60123 5956 60179 6012
rect 60179 5956 60183 6012
rect 60119 5952 60183 5956
rect 60199 6012 60263 6016
rect 60199 5956 60203 6012
rect 60203 5956 60259 6012
rect 60259 5956 60263 6012
rect 60199 5952 60263 5956
rect 60279 6012 60343 6016
rect 60279 5956 60283 6012
rect 60283 5956 60339 6012
rect 60339 5956 60343 6012
rect 60279 5952 60343 5956
rect 60359 6012 60423 6016
rect 60359 5956 60363 6012
rect 60363 5956 60419 6012
rect 60419 5956 60423 6012
rect 60359 5952 60423 5956
rect 99564 6012 99628 6016
rect 99564 5956 99568 6012
rect 99568 5956 99624 6012
rect 99624 5956 99628 6012
rect 99564 5952 99628 5956
rect 99644 6012 99708 6016
rect 99644 5956 99648 6012
rect 99648 5956 99704 6012
rect 99704 5956 99708 6012
rect 99644 5952 99708 5956
rect 99724 6012 99788 6016
rect 99724 5956 99728 6012
rect 99728 5956 99784 6012
rect 99784 5956 99788 6012
rect 99724 5952 99788 5956
rect 99804 6012 99868 6016
rect 99804 5956 99808 6012
rect 99808 5956 99864 6012
rect 99864 5956 99868 6012
rect 99804 5952 99868 5956
rect 124260 5884 124324 5948
rect 139009 6012 139073 6016
rect 139009 5956 139013 6012
rect 139013 5956 139069 6012
rect 139069 5956 139073 6012
rect 139009 5952 139073 5956
rect 139089 6012 139153 6016
rect 139089 5956 139093 6012
rect 139093 5956 139149 6012
rect 139149 5956 139153 6012
rect 139089 5952 139153 5956
rect 139169 6012 139233 6016
rect 139169 5956 139173 6012
rect 139173 5956 139229 6012
rect 139229 5956 139233 6012
rect 139169 5952 139233 5956
rect 139249 6012 139313 6016
rect 139249 5956 139253 6012
rect 139253 5956 139309 6012
rect 139309 5956 139313 6012
rect 139249 5952 139313 5956
rect 150204 5612 150268 5676
rect 151860 5612 151924 5676
rect 155908 5672 155972 5676
rect 155908 5616 155958 5672
rect 155958 5616 155972 5672
rect 155908 5612 155972 5616
rect 147260 5476 147324 5540
rect 40396 5468 40460 5472
rect 40396 5412 40400 5468
rect 40400 5412 40456 5468
rect 40456 5412 40460 5468
rect 40396 5408 40460 5412
rect 40476 5468 40540 5472
rect 40476 5412 40480 5468
rect 40480 5412 40536 5468
rect 40536 5412 40540 5468
rect 40476 5408 40540 5412
rect 40556 5468 40620 5472
rect 40556 5412 40560 5468
rect 40560 5412 40616 5468
rect 40616 5412 40620 5468
rect 40556 5408 40620 5412
rect 40636 5468 40700 5472
rect 40636 5412 40640 5468
rect 40640 5412 40696 5468
rect 40696 5412 40700 5468
rect 40636 5408 40700 5412
rect 79841 5468 79905 5472
rect 79841 5412 79845 5468
rect 79845 5412 79901 5468
rect 79901 5412 79905 5468
rect 79841 5408 79905 5412
rect 79921 5468 79985 5472
rect 79921 5412 79925 5468
rect 79925 5412 79981 5468
rect 79981 5412 79985 5468
rect 79921 5408 79985 5412
rect 80001 5468 80065 5472
rect 80001 5412 80005 5468
rect 80005 5412 80061 5468
rect 80061 5412 80065 5468
rect 80001 5408 80065 5412
rect 80081 5468 80145 5472
rect 80081 5412 80085 5468
rect 80085 5412 80141 5468
rect 80141 5412 80145 5468
rect 80081 5408 80145 5412
rect 119286 5468 119350 5472
rect 119286 5412 119290 5468
rect 119290 5412 119346 5468
rect 119346 5412 119350 5468
rect 119286 5408 119350 5412
rect 119366 5468 119430 5472
rect 119366 5412 119370 5468
rect 119370 5412 119426 5468
rect 119426 5412 119430 5468
rect 119366 5408 119430 5412
rect 119446 5468 119510 5472
rect 119446 5412 119450 5468
rect 119450 5412 119506 5468
rect 119506 5412 119510 5468
rect 119446 5408 119510 5412
rect 119526 5468 119590 5472
rect 119526 5412 119530 5468
rect 119530 5412 119586 5468
rect 119586 5412 119590 5468
rect 119526 5408 119590 5412
rect 158731 5468 158795 5472
rect 158731 5412 158735 5468
rect 158735 5412 158791 5468
rect 158791 5412 158795 5468
rect 158731 5408 158795 5412
rect 158811 5468 158875 5472
rect 158811 5412 158815 5468
rect 158815 5412 158871 5468
rect 158871 5412 158875 5468
rect 158811 5408 158875 5412
rect 158891 5468 158955 5472
rect 158891 5412 158895 5468
rect 158895 5412 158951 5468
rect 158951 5412 158955 5468
rect 158891 5408 158955 5412
rect 158971 5468 159035 5472
rect 158971 5412 158975 5468
rect 158975 5412 159031 5468
rect 159031 5412 159035 5468
rect 158971 5408 159035 5412
rect 147996 5340 148060 5404
rect 156828 5400 156892 5404
rect 156828 5344 156842 5400
rect 156842 5344 156892 5400
rect 156828 5340 156892 5344
rect 148916 5204 148980 5268
rect 147076 5068 147140 5132
rect 154252 5128 154316 5132
rect 154252 5072 154302 5128
rect 154302 5072 154316 5128
rect 154252 5068 154316 5072
rect 20674 4924 20738 4928
rect 20674 4868 20678 4924
rect 20678 4868 20734 4924
rect 20734 4868 20738 4924
rect 20674 4864 20738 4868
rect 20754 4924 20818 4928
rect 20754 4868 20758 4924
rect 20758 4868 20814 4924
rect 20814 4868 20818 4924
rect 20754 4864 20818 4868
rect 20834 4924 20898 4928
rect 20834 4868 20838 4924
rect 20838 4868 20894 4924
rect 20894 4868 20898 4924
rect 20834 4864 20898 4868
rect 20914 4924 20978 4928
rect 20914 4868 20918 4924
rect 20918 4868 20974 4924
rect 20974 4868 20978 4924
rect 20914 4864 20978 4868
rect 60119 4924 60183 4928
rect 60119 4868 60123 4924
rect 60123 4868 60179 4924
rect 60179 4868 60183 4924
rect 60119 4864 60183 4868
rect 60199 4924 60263 4928
rect 60199 4868 60203 4924
rect 60203 4868 60259 4924
rect 60259 4868 60263 4924
rect 60199 4864 60263 4868
rect 60279 4924 60343 4928
rect 60279 4868 60283 4924
rect 60283 4868 60339 4924
rect 60339 4868 60343 4924
rect 60279 4864 60343 4868
rect 60359 4924 60423 4928
rect 60359 4868 60363 4924
rect 60363 4868 60419 4924
rect 60419 4868 60423 4924
rect 60359 4864 60423 4868
rect 99564 4924 99628 4928
rect 99564 4868 99568 4924
rect 99568 4868 99624 4924
rect 99624 4868 99628 4924
rect 99564 4864 99628 4868
rect 99644 4924 99708 4928
rect 99644 4868 99648 4924
rect 99648 4868 99704 4924
rect 99704 4868 99708 4924
rect 99644 4864 99708 4868
rect 99724 4924 99788 4928
rect 99724 4868 99728 4924
rect 99728 4868 99784 4924
rect 99784 4868 99788 4924
rect 99724 4864 99788 4868
rect 99804 4924 99868 4928
rect 99804 4868 99808 4924
rect 99808 4868 99864 4924
rect 99864 4868 99868 4924
rect 99804 4864 99868 4868
rect 139009 4924 139073 4928
rect 139009 4868 139013 4924
rect 139013 4868 139069 4924
rect 139069 4868 139073 4924
rect 139009 4864 139073 4868
rect 139089 4924 139153 4928
rect 139089 4868 139093 4924
rect 139093 4868 139149 4924
rect 139149 4868 139153 4924
rect 139089 4864 139153 4868
rect 139169 4924 139233 4928
rect 139169 4868 139173 4924
rect 139173 4868 139229 4924
rect 139229 4868 139233 4924
rect 139169 4864 139233 4868
rect 139249 4924 139313 4928
rect 139249 4868 139253 4924
rect 139253 4868 139309 4924
rect 139309 4868 139313 4924
rect 139249 4864 139313 4868
rect 40396 4380 40460 4384
rect 40396 4324 40400 4380
rect 40400 4324 40456 4380
rect 40456 4324 40460 4380
rect 40396 4320 40460 4324
rect 40476 4380 40540 4384
rect 40476 4324 40480 4380
rect 40480 4324 40536 4380
rect 40536 4324 40540 4380
rect 40476 4320 40540 4324
rect 40556 4380 40620 4384
rect 40556 4324 40560 4380
rect 40560 4324 40616 4380
rect 40616 4324 40620 4380
rect 40556 4320 40620 4324
rect 40636 4380 40700 4384
rect 40636 4324 40640 4380
rect 40640 4324 40696 4380
rect 40696 4324 40700 4380
rect 40636 4320 40700 4324
rect 79841 4380 79905 4384
rect 79841 4324 79845 4380
rect 79845 4324 79901 4380
rect 79901 4324 79905 4380
rect 79841 4320 79905 4324
rect 79921 4380 79985 4384
rect 79921 4324 79925 4380
rect 79925 4324 79981 4380
rect 79981 4324 79985 4380
rect 79921 4320 79985 4324
rect 80001 4380 80065 4384
rect 80001 4324 80005 4380
rect 80005 4324 80061 4380
rect 80061 4324 80065 4380
rect 80001 4320 80065 4324
rect 80081 4380 80145 4384
rect 80081 4324 80085 4380
rect 80085 4324 80141 4380
rect 80141 4324 80145 4380
rect 80081 4320 80145 4324
rect 119286 4380 119350 4384
rect 119286 4324 119290 4380
rect 119290 4324 119346 4380
rect 119346 4324 119350 4380
rect 119286 4320 119350 4324
rect 119366 4380 119430 4384
rect 119366 4324 119370 4380
rect 119370 4324 119426 4380
rect 119426 4324 119430 4380
rect 119366 4320 119430 4324
rect 119446 4380 119510 4384
rect 119446 4324 119450 4380
rect 119450 4324 119506 4380
rect 119506 4324 119510 4380
rect 119446 4320 119510 4324
rect 119526 4380 119590 4384
rect 119526 4324 119530 4380
rect 119530 4324 119586 4380
rect 119586 4324 119590 4380
rect 119526 4320 119590 4324
rect 158731 4380 158795 4384
rect 158731 4324 158735 4380
rect 158735 4324 158791 4380
rect 158791 4324 158795 4380
rect 158731 4320 158795 4324
rect 158811 4380 158875 4384
rect 158811 4324 158815 4380
rect 158815 4324 158871 4380
rect 158871 4324 158875 4380
rect 158811 4320 158875 4324
rect 158891 4380 158955 4384
rect 158891 4324 158895 4380
rect 158895 4324 158951 4380
rect 158951 4324 158955 4380
rect 158891 4320 158955 4324
rect 158971 4380 159035 4384
rect 158971 4324 158975 4380
rect 158975 4324 159031 4380
rect 159031 4324 159035 4380
rect 158971 4320 159035 4324
rect 153148 4252 153212 4316
rect 152596 4116 152660 4180
rect 155172 4040 155236 4044
rect 155172 3984 155186 4040
rect 155186 3984 155236 4040
rect 155172 3980 155236 3984
rect 155724 4040 155788 4044
rect 155724 3984 155774 4040
rect 155774 3984 155788 4040
rect 155724 3980 155788 3984
rect 20674 3836 20738 3840
rect 20674 3780 20678 3836
rect 20678 3780 20734 3836
rect 20734 3780 20738 3836
rect 20674 3776 20738 3780
rect 20754 3836 20818 3840
rect 20754 3780 20758 3836
rect 20758 3780 20814 3836
rect 20814 3780 20818 3836
rect 20754 3776 20818 3780
rect 20834 3836 20898 3840
rect 20834 3780 20838 3836
rect 20838 3780 20894 3836
rect 20894 3780 20898 3836
rect 20834 3776 20898 3780
rect 20914 3836 20978 3840
rect 20914 3780 20918 3836
rect 20918 3780 20974 3836
rect 20974 3780 20978 3836
rect 20914 3776 20978 3780
rect 60119 3836 60183 3840
rect 60119 3780 60123 3836
rect 60123 3780 60179 3836
rect 60179 3780 60183 3836
rect 60119 3776 60183 3780
rect 60199 3836 60263 3840
rect 60199 3780 60203 3836
rect 60203 3780 60259 3836
rect 60259 3780 60263 3836
rect 60199 3776 60263 3780
rect 60279 3836 60343 3840
rect 60279 3780 60283 3836
rect 60283 3780 60339 3836
rect 60339 3780 60343 3836
rect 60279 3776 60343 3780
rect 60359 3836 60423 3840
rect 60359 3780 60363 3836
rect 60363 3780 60419 3836
rect 60419 3780 60423 3836
rect 60359 3776 60423 3780
rect 99564 3836 99628 3840
rect 99564 3780 99568 3836
rect 99568 3780 99624 3836
rect 99624 3780 99628 3836
rect 99564 3776 99628 3780
rect 99644 3836 99708 3840
rect 99644 3780 99648 3836
rect 99648 3780 99704 3836
rect 99704 3780 99708 3836
rect 99644 3776 99708 3780
rect 99724 3836 99788 3840
rect 99724 3780 99728 3836
rect 99728 3780 99784 3836
rect 99784 3780 99788 3836
rect 99724 3776 99788 3780
rect 99804 3836 99868 3840
rect 99804 3780 99808 3836
rect 99808 3780 99864 3836
rect 99864 3780 99868 3836
rect 99804 3776 99868 3780
rect 139009 3836 139073 3840
rect 139009 3780 139013 3836
rect 139013 3780 139069 3836
rect 139069 3780 139073 3836
rect 139009 3776 139073 3780
rect 139089 3836 139153 3840
rect 139089 3780 139093 3836
rect 139093 3780 139149 3836
rect 139149 3780 139153 3836
rect 139089 3776 139153 3780
rect 139169 3836 139233 3840
rect 139169 3780 139173 3836
rect 139173 3780 139229 3836
rect 139229 3780 139233 3836
rect 139169 3776 139233 3780
rect 139249 3836 139313 3840
rect 139249 3780 139253 3836
rect 139253 3780 139309 3836
rect 139309 3780 139313 3836
rect 139249 3776 139313 3780
rect 151860 3708 151924 3772
rect 152780 3768 152844 3772
rect 152780 3712 152830 3768
rect 152830 3712 152844 3768
rect 152780 3708 152844 3712
rect 154804 3708 154868 3772
rect 151676 3436 151740 3500
rect 40396 3292 40460 3296
rect 40396 3236 40400 3292
rect 40400 3236 40456 3292
rect 40456 3236 40460 3292
rect 40396 3232 40460 3236
rect 40476 3292 40540 3296
rect 40476 3236 40480 3292
rect 40480 3236 40536 3292
rect 40536 3236 40540 3292
rect 40476 3232 40540 3236
rect 40556 3292 40620 3296
rect 40556 3236 40560 3292
rect 40560 3236 40616 3292
rect 40616 3236 40620 3292
rect 40556 3232 40620 3236
rect 40636 3292 40700 3296
rect 40636 3236 40640 3292
rect 40640 3236 40696 3292
rect 40696 3236 40700 3292
rect 40636 3232 40700 3236
rect 79841 3292 79905 3296
rect 79841 3236 79845 3292
rect 79845 3236 79901 3292
rect 79901 3236 79905 3292
rect 79841 3232 79905 3236
rect 79921 3292 79985 3296
rect 79921 3236 79925 3292
rect 79925 3236 79981 3292
rect 79981 3236 79985 3292
rect 79921 3232 79985 3236
rect 80001 3292 80065 3296
rect 80001 3236 80005 3292
rect 80005 3236 80061 3292
rect 80061 3236 80065 3292
rect 80001 3232 80065 3236
rect 80081 3292 80145 3296
rect 80081 3236 80085 3292
rect 80085 3236 80141 3292
rect 80141 3236 80145 3292
rect 80081 3232 80145 3236
rect 119286 3292 119350 3296
rect 119286 3236 119290 3292
rect 119290 3236 119346 3292
rect 119346 3236 119350 3292
rect 119286 3232 119350 3236
rect 119366 3292 119430 3296
rect 119366 3236 119370 3292
rect 119370 3236 119426 3292
rect 119426 3236 119430 3292
rect 119366 3232 119430 3236
rect 119446 3292 119510 3296
rect 119446 3236 119450 3292
rect 119450 3236 119506 3292
rect 119506 3236 119510 3292
rect 119446 3232 119510 3236
rect 119526 3292 119590 3296
rect 119526 3236 119530 3292
rect 119530 3236 119586 3292
rect 119586 3236 119590 3292
rect 119526 3232 119590 3236
rect 158731 3292 158795 3296
rect 158731 3236 158735 3292
rect 158735 3236 158791 3292
rect 158791 3236 158795 3292
rect 158731 3232 158795 3236
rect 158811 3292 158875 3296
rect 158811 3236 158815 3292
rect 158815 3236 158871 3292
rect 158871 3236 158875 3292
rect 158811 3232 158875 3236
rect 158891 3292 158955 3296
rect 158891 3236 158895 3292
rect 158895 3236 158951 3292
rect 158951 3236 158955 3292
rect 158891 3232 158955 3236
rect 158971 3292 159035 3296
rect 158971 3236 158975 3292
rect 158975 3236 159031 3292
rect 159031 3236 159035 3292
rect 158971 3232 159035 3236
rect 20674 2748 20738 2752
rect 20674 2692 20678 2748
rect 20678 2692 20734 2748
rect 20734 2692 20738 2748
rect 20674 2688 20738 2692
rect 20754 2748 20818 2752
rect 20754 2692 20758 2748
rect 20758 2692 20814 2748
rect 20814 2692 20818 2748
rect 20754 2688 20818 2692
rect 20834 2748 20898 2752
rect 20834 2692 20838 2748
rect 20838 2692 20894 2748
rect 20894 2692 20898 2748
rect 20834 2688 20898 2692
rect 20914 2748 20978 2752
rect 20914 2692 20918 2748
rect 20918 2692 20974 2748
rect 20974 2692 20978 2748
rect 20914 2688 20978 2692
rect 60119 2748 60183 2752
rect 60119 2692 60123 2748
rect 60123 2692 60179 2748
rect 60179 2692 60183 2748
rect 60119 2688 60183 2692
rect 60199 2748 60263 2752
rect 60199 2692 60203 2748
rect 60203 2692 60259 2748
rect 60259 2692 60263 2748
rect 60199 2688 60263 2692
rect 60279 2748 60343 2752
rect 60279 2692 60283 2748
rect 60283 2692 60339 2748
rect 60339 2692 60343 2748
rect 60279 2688 60343 2692
rect 60359 2748 60423 2752
rect 60359 2692 60363 2748
rect 60363 2692 60419 2748
rect 60419 2692 60423 2748
rect 60359 2688 60423 2692
rect 99564 2748 99628 2752
rect 99564 2692 99568 2748
rect 99568 2692 99624 2748
rect 99624 2692 99628 2748
rect 99564 2688 99628 2692
rect 99644 2748 99708 2752
rect 99644 2692 99648 2748
rect 99648 2692 99704 2748
rect 99704 2692 99708 2748
rect 99644 2688 99708 2692
rect 99724 2748 99788 2752
rect 99724 2692 99728 2748
rect 99728 2692 99784 2748
rect 99784 2692 99788 2748
rect 99724 2688 99788 2692
rect 99804 2748 99868 2752
rect 99804 2692 99808 2748
rect 99808 2692 99864 2748
rect 99864 2692 99868 2748
rect 99804 2688 99868 2692
rect 139009 2748 139073 2752
rect 139009 2692 139013 2748
rect 139013 2692 139069 2748
rect 139069 2692 139073 2748
rect 139009 2688 139073 2692
rect 139089 2748 139153 2752
rect 139089 2692 139093 2748
rect 139093 2692 139149 2748
rect 139149 2692 139153 2748
rect 139089 2688 139153 2692
rect 139169 2748 139233 2752
rect 139169 2692 139173 2748
rect 139173 2692 139229 2748
rect 139229 2692 139233 2748
rect 139169 2688 139233 2692
rect 139249 2748 139313 2752
rect 139249 2692 139253 2748
rect 139253 2692 139309 2748
rect 139309 2692 139313 2748
rect 139249 2688 139313 2692
rect 40396 2204 40460 2208
rect 40396 2148 40400 2204
rect 40400 2148 40456 2204
rect 40456 2148 40460 2204
rect 40396 2144 40460 2148
rect 40476 2204 40540 2208
rect 40476 2148 40480 2204
rect 40480 2148 40536 2204
rect 40536 2148 40540 2204
rect 40476 2144 40540 2148
rect 40556 2204 40620 2208
rect 40556 2148 40560 2204
rect 40560 2148 40616 2204
rect 40616 2148 40620 2204
rect 40556 2144 40620 2148
rect 40636 2204 40700 2208
rect 40636 2148 40640 2204
rect 40640 2148 40696 2204
rect 40696 2148 40700 2204
rect 40636 2144 40700 2148
rect 79841 2204 79905 2208
rect 79841 2148 79845 2204
rect 79845 2148 79901 2204
rect 79901 2148 79905 2204
rect 79841 2144 79905 2148
rect 79921 2204 79985 2208
rect 79921 2148 79925 2204
rect 79925 2148 79981 2204
rect 79981 2148 79985 2204
rect 79921 2144 79985 2148
rect 80001 2204 80065 2208
rect 80001 2148 80005 2204
rect 80005 2148 80061 2204
rect 80061 2148 80065 2204
rect 80001 2144 80065 2148
rect 80081 2204 80145 2208
rect 80081 2148 80085 2204
rect 80085 2148 80141 2204
rect 80141 2148 80145 2204
rect 80081 2144 80145 2148
rect 119286 2204 119350 2208
rect 119286 2148 119290 2204
rect 119290 2148 119346 2204
rect 119346 2148 119350 2204
rect 119286 2144 119350 2148
rect 119366 2204 119430 2208
rect 119366 2148 119370 2204
rect 119370 2148 119426 2204
rect 119426 2148 119430 2204
rect 119366 2144 119430 2148
rect 119446 2204 119510 2208
rect 119446 2148 119450 2204
rect 119450 2148 119506 2204
rect 119506 2148 119510 2204
rect 119446 2144 119510 2148
rect 119526 2204 119590 2208
rect 119526 2148 119530 2204
rect 119530 2148 119586 2204
rect 119586 2148 119590 2204
rect 119526 2144 119590 2148
rect 158731 2204 158795 2208
rect 158731 2148 158735 2204
rect 158735 2148 158791 2204
rect 158791 2148 158795 2204
rect 158731 2144 158795 2148
rect 158811 2204 158875 2208
rect 158811 2148 158815 2204
rect 158815 2148 158871 2204
rect 158871 2148 158875 2204
rect 158811 2144 158875 2148
rect 158891 2204 158955 2208
rect 158891 2148 158895 2204
rect 158895 2148 158951 2204
rect 158951 2148 158955 2204
rect 158891 2144 158955 2148
rect 158971 2204 159035 2208
rect 158971 2148 158975 2204
rect 158975 2148 159031 2204
rect 159031 2148 159035 2204
rect 158971 2144 159035 2148
rect 131068 2076 131132 2140
rect 153332 1804 153396 1868
rect 155908 1260 155972 1324
rect 124444 1124 124508 1188
<< metal4 >>
rect 150755 14516 150821 14517
rect 150755 14452 150756 14516
rect 150820 14452 150821 14516
rect 150755 14451 150821 14452
rect 20666 13632 20986 13648
rect 20666 13568 20674 13632
rect 20738 13568 20754 13632
rect 20818 13568 20834 13632
rect 20898 13568 20914 13632
rect 20978 13568 20986 13632
rect 20666 12544 20986 13568
rect 20666 12480 20674 12544
rect 20738 12480 20754 12544
rect 20818 12480 20834 12544
rect 20898 12480 20914 12544
rect 20978 12480 20986 12544
rect 20666 11456 20986 12480
rect 20666 11392 20674 11456
rect 20738 11392 20754 11456
rect 20818 11392 20834 11456
rect 20898 11392 20914 11456
rect 20978 11392 20986 11456
rect 20666 10368 20986 11392
rect 20666 10304 20674 10368
rect 20738 10304 20754 10368
rect 20818 10304 20834 10368
rect 20898 10304 20914 10368
rect 20978 10304 20986 10368
rect 20666 9280 20986 10304
rect 20666 9216 20674 9280
rect 20738 9216 20754 9280
rect 20818 9216 20834 9280
rect 20898 9216 20914 9280
rect 20978 9216 20986 9280
rect 20666 8192 20986 9216
rect 20666 8128 20674 8192
rect 20738 8128 20754 8192
rect 20818 8128 20834 8192
rect 20898 8128 20914 8192
rect 20978 8128 20986 8192
rect 20666 7104 20986 8128
rect 20666 7040 20674 7104
rect 20738 7040 20754 7104
rect 20818 7040 20834 7104
rect 20898 7040 20914 7104
rect 20978 7040 20986 7104
rect 20666 6016 20986 7040
rect 20666 5952 20674 6016
rect 20738 5952 20754 6016
rect 20818 5952 20834 6016
rect 20898 5952 20914 6016
rect 20978 5952 20986 6016
rect 20666 4928 20986 5952
rect 20666 4864 20674 4928
rect 20738 4864 20754 4928
rect 20818 4864 20834 4928
rect 20898 4864 20914 4928
rect 20978 4864 20986 4928
rect 20666 3840 20986 4864
rect 20666 3776 20674 3840
rect 20738 3776 20754 3840
rect 20818 3776 20834 3840
rect 20898 3776 20914 3840
rect 20978 3776 20986 3840
rect 20666 2752 20986 3776
rect 20666 2688 20674 2752
rect 20738 2688 20754 2752
rect 20818 2688 20834 2752
rect 20898 2688 20914 2752
rect 20978 2688 20986 2752
rect 20666 2128 20986 2688
rect 40388 13088 40708 13648
rect 40388 13024 40396 13088
rect 40460 13024 40476 13088
rect 40540 13024 40556 13088
rect 40620 13024 40636 13088
rect 40700 13024 40708 13088
rect 40388 12000 40708 13024
rect 40388 11936 40396 12000
rect 40460 11936 40476 12000
rect 40540 11936 40556 12000
rect 40620 11936 40636 12000
rect 40700 11936 40708 12000
rect 40388 10912 40708 11936
rect 40388 10848 40396 10912
rect 40460 10848 40476 10912
rect 40540 10848 40556 10912
rect 40620 10848 40636 10912
rect 40700 10848 40708 10912
rect 40388 9824 40708 10848
rect 40388 9760 40396 9824
rect 40460 9760 40476 9824
rect 40540 9760 40556 9824
rect 40620 9760 40636 9824
rect 40700 9760 40708 9824
rect 40388 8736 40708 9760
rect 40388 8672 40396 8736
rect 40460 8672 40476 8736
rect 40540 8672 40556 8736
rect 40620 8672 40636 8736
rect 40700 8672 40708 8736
rect 40388 7648 40708 8672
rect 40388 7584 40396 7648
rect 40460 7584 40476 7648
rect 40540 7584 40556 7648
rect 40620 7584 40636 7648
rect 40700 7584 40708 7648
rect 40388 6560 40708 7584
rect 40388 6496 40396 6560
rect 40460 6496 40476 6560
rect 40540 6496 40556 6560
rect 40620 6496 40636 6560
rect 40700 6496 40708 6560
rect 40388 5472 40708 6496
rect 40388 5408 40396 5472
rect 40460 5408 40476 5472
rect 40540 5408 40556 5472
rect 40620 5408 40636 5472
rect 40700 5408 40708 5472
rect 40388 4384 40708 5408
rect 40388 4320 40396 4384
rect 40460 4320 40476 4384
rect 40540 4320 40556 4384
rect 40620 4320 40636 4384
rect 40700 4320 40708 4384
rect 40388 3296 40708 4320
rect 40388 3232 40396 3296
rect 40460 3232 40476 3296
rect 40540 3232 40556 3296
rect 40620 3232 40636 3296
rect 40700 3232 40708 3296
rect 40388 2208 40708 3232
rect 40388 2144 40396 2208
rect 40460 2144 40476 2208
rect 40540 2144 40556 2208
rect 40620 2144 40636 2208
rect 40700 2144 40708 2208
rect 40388 2128 40708 2144
rect 60111 13632 60431 13648
rect 60111 13568 60119 13632
rect 60183 13568 60199 13632
rect 60263 13568 60279 13632
rect 60343 13568 60359 13632
rect 60423 13568 60431 13632
rect 60111 12544 60431 13568
rect 60111 12480 60119 12544
rect 60183 12480 60199 12544
rect 60263 12480 60279 12544
rect 60343 12480 60359 12544
rect 60423 12480 60431 12544
rect 60111 11456 60431 12480
rect 60111 11392 60119 11456
rect 60183 11392 60199 11456
rect 60263 11392 60279 11456
rect 60343 11392 60359 11456
rect 60423 11392 60431 11456
rect 60111 10368 60431 11392
rect 60111 10304 60119 10368
rect 60183 10304 60199 10368
rect 60263 10304 60279 10368
rect 60343 10304 60359 10368
rect 60423 10304 60431 10368
rect 60111 9280 60431 10304
rect 60111 9216 60119 9280
rect 60183 9216 60199 9280
rect 60263 9216 60279 9280
rect 60343 9216 60359 9280
rect 60423 9216 60431 9280
rect 60111 8192 60431 9216
rect 60111 8128 60119 8192
rect 60183 8128 60199 8192
rect 60263 8128 60279 8192
rect 60343 8128 60359 8192
rect 60423 8128 60431 8192
rect 60111 7104 60431 8128
rect 60111 7040 60119 7104
rect 60183 7040 60199 7104
rect 60263 7040 60279 7104
rect 60343 7040 60359 7104
rect 60423 7040 60431 7104
rect 60111 6016 60431 7040
rect 60111 5952 60119 6016
rect 60183 5952 60199 6016
rect 60263 5952 60279 6016
rect 60343 5952 60359 6016
rect 60423 5952 60431 6016
rect 60111 4928 60431 5952
rect 60111 4864 60119 4928
rect 60183 4864 60199 4928
rect 60263 4864 60279 4928
rect 60343 4864 60359 4928
rect 60423 4864 60431 4928
rect 60111 3840 60431 4864
rect 60111 3776 60119 3840
rect 60183 3776 60199 3840
rect 60263 3776 60279 3840
rect 60343 3776 60359 3840
rect 60423 3776 60431 3840
rect 60111 2752 60431 3776
rect 60111 2688 60119 2752
rect 60183 2688 60199 2752
rect 60263 2688 60279 2752
rect 60343 2688 60359 2752
rect 60423 2688 60431 2752
rect 60111 2128 60431 2688
rect 79833 13088 80153 13648
rect 79833 13024 79841 13088
rect 79905 13024 79921 13088
rect 79985 13024 80001 13088
rect 80065 13024 80081 13088
rect 80145 13024 80153 13088
rect 79833 12000 80153 13024
rect 79833 11936 79841 12000
rect 79905 11936 79921 12000
rect 79985 11936 80001 12000
rect 80065 11936 80081 12000
rect 80145 11936 80153 12000
rect 79833 10912 80153 11936
rect 79833 10848 79841 10912
rect 79905 10848 79921 10912
rect 79985 10848 80001 10912
rect 80065 10848 80081 10912
rect 80145 10848 80153 10912
rect 79833 9824 80153 10848
rect 79833 9760 79841 9824
rect 79905 9760 79921 9824
rect 79985 9760 80001 9824
rect 80065 9760 80081 9824
rect 80145 9760 80153 9824
rect 79833 8736 80153 9760
rect 79833 8672 79841 8736
rect 79905 8672 79921 8736
rect 79985 8672 80001 8736
rect 80065 8672 80081 8736
rect 80145 8672 80153 8736
rect 79833 7648 80153 8672
rect 79833 7584 79841 7648
rect 79905 7584 79921 7648
rect 79985 7584 80001 7648
rect 80065 7584 80081 7648
rect 80145 7584 80153 7648
rect 79833 6560 80153 7584
rect 79833 6496 79841 6560
rect 79905 6496 79921 6560
rect 79985 6496 80001 6560
rect 80065 6496 80081 6560
rect 80145 6496 80153 6560
rect 79833 5472 80153 6496
rect 79833 5408 79841 5472
rect 79905 5408 79921 5472
rect 79985 5408 80001 5472
rect 80065 5408 80081 5472
rect 80145 5408 80153 5472
rect 79833 4384 80153 5408
rect 79833 4320 79841 4384
rect 79905 4320 79921 4384
rect 79985 4320 80001 4384
rect 80065 4320 80081 4384
rect 80145 4320 80153 4384
rect 79833 3296 80153 4320
rect 79833 3232 79841 3296
rect 79905 3232 79921 3296
rect 79985 3232 80001 3296
rect 80065 3232 80081 3296
rect 80145 3232 80153 3296
rect 79833 2208 80153 3232
rect 79833 2144 79841 2208
rect 79905 2144 79921 2208
rect 79985 2144 80001 2208
rect 80065 2144 80081 2208
rect 80145 2144 80153 2208
rect 79833 2128 80153 2144
rect 99556 13632 99876 13648
rect 99556 13568 99564 13632
rect 99628 13568 99644 13632
rect 99708 13568 99724 13632
rect 99788 13568 99804 13632
rect 99868 13568 99876 13632
rect 99556 12544 99876 13568
rect 99556 12480 99564 12544
rect 99628 12480 99644 12544
rect 99708 12480 99724 12544
rect 99788 12480 99804 12544
rect 99868 12480 99876 12544
rect 99556 11456 99876 12480
rect 99556 11392 99564 11456
rect 99628 11392 99644 11456
rect 99708 11392 99724 11456
rect 99788 11392 99804 11456
rect 99868 11392 99876 11456
rect 99556 10368 99876 11392
rect 99556 10304 99564 10368
rect 99628 10304 99644 10368
rect 99708 10304 99724 10368
rect 99788 10304 99804 10368
rect 99868 10304 99876 10368
rect 99556 9280 99876 10304
rect 99556 9216 99564 9280
rect 99628 9216 99644 9280
rect 99708 9216 99724 9280
rect 99788 9216 99804 9280
rect 99868 9216 99876 9280
rect 99556 8192 99876 9216
rect 99556 8128 99564 8192
rect 99628 8128 99644 8192
rect 99708 8128 99724 8192
rect 99788 8128 99804 8192
rect 99868 8128 99876 8192
rect 99556 7104 99876 8128
rect 99556 7040 99564 7104
rect 99628 7040 99644 7104
rect 99708 7040 99724 7104
rect 99788 7040 99804 7104
rect 99868 7040 99876 7104
rect 99556 6016 99876 7040
rect 99556 5952 99564 6016
rect 99628 5952 99644 6016
rect 99708 5952 99724 6016
rect 99788 5952 99804 6016
rect 99868 5952 99876 6016
rect 99556 4928 99876 5952
rect 99556 4864 99564 4928
rect 99628 4864 99644 4928
rect 99708 4864 99724 4928
rect 99788 4864 99804 4928
rect 99868 4864 99876 4928
rect 99556 3840 99876 4864
rect 99556 3776 99564 3840
rect 99628 3776 99644 3840
rect 99708 3776 99724 3840
rect 99788 3776 99804 3840
rect 99868 3776 99876 3840
rect 99556 2752 99876 3776
rect 99556 2688 99564 2752
rect 99628 2688 99644 2752
rect 99708 2688 99724 2752
rect 99788 2688 99804 2752
rect 99868 2688 99876 2752
rect 99556 2128 99876 2688
rect 119278 13088 119598 13648
rect 119278 13024 119286 13088
rect 119350 13024 119366 13088
rect 119430 13024 119446 13088
rect 119510 13024 119526 13088
rect 119590 13024 119598 13088
rect 119278 12000 119598 13024
rect 139001 13632 139321 13648
rect 139001 13568 139009 13632
rect 139073 13568 139089 13632
rect 139153 13568 139169 13632
rect 139233 13568 139249 13632
rect 139313 13568 139321 13632
rect 139001 12544 139321 13568
rect 149651 13020 149717 13021
rect 149651 12956 149652 13020
rect 149716 12956 149717 13020
rect 149651 12955 149717 12956
rect 139001 12480 139009 12544
rect 139073 12480 139089 12544
rect 139153 12480 139169 12544
rect 139233 12480 139249 12544
rect 139313 12480 139321 12544
rect 127203 12068 127269 12069
rect 127203 12004 127204 12068
rect 127268 12004 127269 12068
rect 127203 12003 127269 12004
rect 119278 11936 119286 12000
rect 119350 11936 119366 12000
rect 119430 11936 119446 12000
rect 119510 11936 119526 12000
rect 119590 11936 119598 12000
rect 119278 10912 119598 11936
rect 119278 10848 119286 10912
rect 119350 10848 119366 10912
rect 119430 10848 119446 10912
rect 119510 10848 119526 10912
rect 119590 10848 119598 10912
rect 119278 9824 119598 10848
rect 119278 9760 119286 9824
rect 119350 9760 119366 9824
rect 119430 9760 119446 9824
rect 119510 9760 119526 9824
rect 119590 9760 119598 9824
rect 119278 8736 119598 9760
rect 124443 9756 124509 9757
rect 124443 9692 124444 9756
rect 124508 9692 124509 9756
rect 124443 9691 124509 9692
rect 119278 8672 119286 8736
rect 119350 8672 119366 8736
rect 119430 8672 119446 8736
rect 119510 8672 119526 8736
rect 119590 8672 119598 8736
rect 119278 7648 119598 8672
rect 124259 8396 124325 8397
rect 124259 8332 124260 8396
rect 124324 8332 124325 8396
rect 124259 8331 124325 8332
rect 119278 7584 119286 7648
rect 119350 7584 119366 7648
rect 119430 7584 119446 7648
rect 119510 7584 119526 7648
rect 119590 7584 119598 7648
rect 119278 6560 119598 7584
rect 119278 6496 119286 6560
rect 119350 6496 119366 6560
rect 119430 6496 119446 6560
rect 119510 6496 119526 6560
rect 119590 6496 119598 6560
rect 119278 5472 119598 6496
rect 124262 5949 124322 8331
rect 124259 5948 124325 5949
rect 124259 5884 124260 5948
rect 124324 5884 124325 5948
rect 124259 5883 124325 5884
rect 119278 5408 119286 5472
rect 119350 5408 119366 5472
rect 119430 5408 119446 5472
rect 119510 5408 119526 5472
rect 119590 5408 119598 5472
rect 119278 4384 119598 5408
rect 119278 4320 119286 4384
rect 119350 4320 119366 4384
rect 119430 4320 119446 4384
rect 119510 4320 119526 4384
rect 119590 4320 119598 4384
rect 119278 3296 119598 4320
rect 119278 3232 119286 3296
rect 119350 3232 119366 3296
rect 119430 3232 119446 3296
rect 119510 3232 119526 3296
rect 119590 3232 119598 3296
rect 119278 2208 119598 3232
rect 119278 2144 119286 2208
rect 119350 2144 119366 2208
rect 119430 2144 119446 2208
rect 119510 2144 119526 2208
rect 119590 2144 119598 2208
rect 119278 2128 119598 2144
rect 124446 1189 124506 9691
rect 127206 8805 127266 12003
rect 131067 11932 131133 11933
rect 131067 11868 131068 11932
rect 131132 11868 131133 11932
rect 131067 11867 131133 11868
rect 127203 8804 127269 8805
rect 127203 8740 127204 8804
rect 127268 8740 127269 8804
rect 127203 8739 127269 8740
rect 127206 6629 127266 8739
rect 131070 7173 131130 11867
rect 133459 11796 133525 11797
rect 133459 11732 133460 11796
rect 133524 11732 133525 11796
rect 133459 11731 133525 11732
rect 131067 7172 131133 7173
rect 131067 7108 131068 7172
rect 131132 7108 131133 7172
rect 131067 7107 131133 7108
rect 127203 6628 127269 6629
rect 127203 6564 127204 6628
rect 127268 6564 127269 6628
rect 127203 6563 127269 6564
rect 131070 2141 131130 7107
rect 133462 6901 133522 11731
rect 139001 11456 139321 12480
rect 147995 11932 148061 11933
rect 147995 11868 147996 11932
rect 148060 11868 148061 11932
rect 147995 11867 148061 11868
rect 139001 11392 139009 11456
rect 139073 11392 139089 11456
rect 139153 11392 139169 11456
rect 139233 11392 139249 11456
rect 139313 11392 139321 11456
rect 139001 10368 139321 11392
rect 147443 11116 147509 11117
rect 147443 11052 147444 11116
rect 147508 11052 147509 11116
rect 147443 11051 147509 11052
rect 146339 10980 146405 10981
rect 146339 10916 146340 10980
rect 146404 10916 146405 10980
rect 146339 10915 146405 10916
rect 139001 10304 139009 10368
rect 139073 10304 139089 10368
rect 139153 10304 139169 10368
rect 139233 10304 139249 10368
rect 139313 10304 139321 10368
rect 139001 9280 139321 10304
rect 139001 9216 139009 9280
rect 139073 9216 139089 9280
rect 139153 9216 139169 9280
rect 139233 9216 139249 9280
rect 139313 9216 139321 9280
rect 139001 8192 139321 9216
rect 139715 8940 139781 8941
rect 139715 8876 139716 8940
rect 139780 8876 139781 8940
rect 139715 8875 139781 8876
rect 139001 8128 139009 8192
rect 139073 8128 139089 8192
rect 139153 8128 139169 8192
rect 139233 8128 139249 8192
rect 139313 8128 139321 8192
rect 139001 7104 139321 8128
rect 139001 7040 139009 7104
rect 139073 7040 139089 7104
rect 139153 7040 139169 7104
rect 139233 7040 139249 7104
rect 139313 7040 139321 7104
rect 133459 6900 133525 6901
rect 133459 6836 133460 6900
rect 133524 6836 133525 6900
rect 133459 6835 133525 6836
rect 139001 6016 139321 7040
rect 139718 6357 139778 8875
rect 145051 8260 145117 8261
rect 145051 8196 145052 8260
rect 145116 8196 145117 8260
rect 145051 8195 145117 8196
rect 145054 7037 145114 8195
rect 145051 7036 145117 7037
rect 145051 6972 145052 7036
rect 145116 6972 145117 7036
rect 145051 6971 145117 6972
rect 146342 6493 146402 10915
rect 147075 8668 147141 8669
rect 147075 8604 147076 8668
rect 147140 8604 147141 8668
rect 147075 8603 147141 8604
rect 146891 8124 146957 8125
rect 146891 8060 146892 8124
rect 146956 8060 146957 8124
rect 146891 8059 146957 8060
rect 146894 7173 146954 8059
rect 146891 7172 146957 7173
rect 146891 7108 146892 7172
rect 146956 7108 146957 7172
rect 146891 7107 146957 7108
rect 146339 6492 146405 6493
rect 146339 6428 146340 6492
rect 146404 6428 146405 6492
rect 146339 6427 146405 6428
rect 139715 6356 139781 6357
rect 139715 6292 139716 6356
rect 139780 6292 139781 6356
rect 139715 6291 139781 6292
rect 139001 5952 139009 6016
rect 139073 5952 139089 6016
rect 139153 5952 139169 6016
rect 139233 5952 139249 6016
rect 139313 5952 139321 6016
rect 139001 4928 139321 5952
rect 147078 5133 147138 8603
rect 147259 8124 147325 8125
rect 147259 8060 147260 8124
rect 147324 8060 147325 8124
rect 147259 8059 147325 8060
rect 147262 5541 147322 8059
rect 147446 7173 147506 11051
rect 147443 7172 147509 7173
rect 147443 7108 147444 7172
rect 147508 7108 147509 7172
rect 147443 7107 147509 7108
rect 147811 7172 147877 7173
rect 147811 7108 147812 7172
rect 147876 7108 147877 7172
rect 147811 7107 147877 7108
rect 147814 6901 147874 7107
rect 147811 6900 147877 6901
rect 147811 6836 147812 6900
rect 147876 6836 147877 6900
rect 147811 6835 147877 6836
rect 147259 5540 147325 5541
rect 147259 5476 147260 5540
rect 147324 5476 147325 5540
rect 147259 5475 147325 5476
rect 147998 5405 148058 11867
rect 148547 8940 148613 8941
rect 148547 8876 148548 8940
rect 148612 8938 148613 8940
rect 148612 8878 149346 8938
rect 148612 8876 148613 8878
rect 148547 8875 148613 8876
rect 148915 8260 148981 8261
rect 148915 8196 148916 8260
rect 148980 8196 148981 8260
rect 148915 8195 148981 8196
rect 147995 5404 148061 5405
rect 147995 5340 147996 5404
rect 148060 5340 148061 5404
rect 147995 5339 148061 5340
rect 148918 5269 148978 8195
rect 149286 6221 149346 8878
rect 149654 8669 149714 12955
rect 150387 10300 150453 10301
rect 150387 10236 150388 10300
rect 150452 10236 150453 10300
rect 150387 10235 150453 10236
rect 150390 8805 150450 10235
rect 150387 8804 150453 8805
rect 150387 8740 150388 8804
rect 150452 8740 150453 8804
rect 150387 8739 150453 8740
rect 149651 8668 149717 8669
rect 149651 8604 149652 8668
rect 149716 8604 149717 8668
rect 149651 8603 149717 8604
rect 150203 8668 150269 8669
rect 150203 8604 150204 8668
rect 150268 8604 150269 8668
rect 150203 8603 150269 8604
rect 149283 6220 149349 6221
rect 149283 6156 149284 6220
rect 149348 6156 149349 6220
rect 149283 6155 149349 6156
rect 150206 5677 150266 8603
rect 150387 8260 150453 8261
rect 150387 8196 150388 8260
rect 150452 8196 150453 8260
rect 150387 8195 150453 8196
rect 150390 7445 150450 8195
rect 150758 7581 150818 14451
rect 156827 14244 156893 14245
rect 156827 14180 156828 14244
rect 156892 14180 156893 14244
rect 156827 14179 156893 14180
rect 155723 14108 155789 14109
rect 155723 14044 155724 14108
rect 155788 14044 155789 14108
rect 155723 14043 155789 14044
rect 155171 13972 155237 13973
rect 155171 13908 155172 13972
rect 155236 13908 155237 13972
rect 155171 13907 155237 13908
rect 152779 11116 152845 11117
rect 152779 11052 152780 11116
rect 152844 11052 152845 11116
rect 152779 11051 152845 11052
rect 152595 9620 152661 9621
rect 152595 9556 152596 9620
rect 152660 9556 152661 9620
rect 152595 9555 152661 9556
rect 151675 8260 151741 8261
rect 151675 8196 151676 8260
rect 151740 8196 151741 8260
rect 151675 8195 151741 8196
rect 150755 7580 150821 7581
rect 150755 7516 150756 7580
rect 150820 7516 150821 7580
rect 150755 7515 150821 7516
rect 150387 7444 150453 7445
rect 150387 7380 150388 7444
rect 150452 7380 150453 7444
rect 150387 7379 150453 7380
rect 150203 5676 150269 5677
rect 150203 5612 150204 5676
rect 150268 5612 150269 5676
rect 150203 5611 150269 5612
rect 148915 5268 148981 5269
rect 148915 5204 148916 5268
rect 148980 5204 148981 5268
rect 148915 5203 148981 5204
rect 147075 5132 147141 5133
rect 147075 5068 147076 5132
rect 147140 5068 147141 5132
rect 147075 5067 147141 5068
rect 139001 4864 139009 4928
rect 139073 4864 139089 4928
rect 139153 4864 139169 4928
rect 139233 4864 139249 4928
rect 139313 4864 139321 4928
rect 139001 3840 139321 4864
rect 139001 3776 139009 3840
rect 139073 3776 139089 3840
rect 139153 3776 139169 3840
rect 139233 3776 139249 3840
rect 139313 3776 139321 3840
rect 139001 2752 139321 3776
rect 151678 3501 151738 8195
rect 151859 5676 151925 5677
rect 151859 5612 151860 5676
rect 151924 5612 151925 5676
rect 151859 5611 151925 5612
rect 151862 3773 151922 5611
rect 152598 4181 152658 9555
rect 152595 4180 152661 4181
rect 152595 4116 152596 4180
rect 152660 4116 152661 4180
rect 152595 4115 152661 4116
rect 152782 3773 152842 11051
rect 154803 8940 154869 8941
rect 154803 8876 154804 8940
rect 154868 8876 154869 8940
rect 154803 8875 154869 8876
rect 153147 8396 153213 8397
rect 153147 8332 153148 8396
rect 153212 8332 153213 8396
rect 153147 8331 153213 8332
rect 153150 4317 153210 8331
rect 154251 7852 154317 7853
rect 154251 7788 154252 7852
rect 154316 7788 154317 7852
rect 154251 7787 154317 7788
rect 153331 7036 153397 7037
rect 153331 6972 153332 7036
rect 153396 6972 153397 7036
rect 153331 6971 153397 6972
rect 153147 4316 153213 4317
rect 153147 4252 153148 4316
rect 153212 4252 153213 4316
rect 153147 4251 153213 4252
rect 151859 3772 151925 3773
rect 151859 3708 151860 3772
rect 151924 3708 151925 3772
rect 151859 3707 151925 3708
rect 152779 3772 152845 3773
rect 152779 3708 152780 3772
rect 152844 3708 152845 3772
rect 152779 3707 152845 3708
rect 151675 3500 151741 3501
rect 151675 3436 151676 3500
rect 151740 3436 151741 3500
rect 151675 3435 151741 3436
rect 139001 2688 139009 2752
rect 139073 2688 139089 2752
rect 139153 2688 139169 2752
rect 139233 2688 139249 2752
rect 139313 2688 139321 2752
rect 131067 2140 131133 2141
rect 131067 2076 131068 2140
rect 131132 2076 131133 2140
rect 139001 2128 139321 2688
rect 131067 2075 131133 2076
rect 153334 1869 153394 6971
rect 154254 5133 154314 7787
rect 154251 5132 154317 5133
rect 154251 5068 154252 5132
rect 154316 5068 154317 5132
rect 154251 5067 154317 5068
rect 154806 3773 154866 8875
rect 155174 4045 155234 13907
rect 155726 4045 155786 14043
rect 155907 5676 155973 5677
rect 155907 5612 155908 5676
rect 155972 5612 155973 5676
rect 155907 5611 155973 5612
rect 155171 4044 155237 4045
rect 155171 3980 155172 4044
rect 155236 3980 155237 4044
rect 155171 3979 155237 3980
rect 155723 4044 155789 4045
rect 155723 3980 155724 4044
rect 155788 3980 155789 4044
rect 155723 3979 155789 3980
rect 154803 3772 154869 3773
rect 154803 3708 154804 3772
rect 154868 3708 154869 3772
rect 154803 3707 154869 3708
rect 153331 1868 153397 1869
rect 153331 1804 153332 1868
rect 153396 1804 153397 1868
rect 153331 1803 153397 1804
rect 155910 1325 155970 5611
rect 156830 5405 156890 14179
rect 158723 13088 159043 13648
rect 158723 13024 158731 13088
rect 158795 13024 158811 13088
rect 158875 13024 158891 13088
rect 158955 13024 158971 13088
rect 159035 13024 159043 13088
rect 158723 12000 159043 13024
rect 158723 11936 158731 12000
rect 158795 11936 158811 12000
rect 158875 11936 158891 12000
rect 158955 11936 158971 12000
rect 159035 11936 159043 12000
rect 158723 10912 159043 11936
rect 158723 10848 158731 10912
rect 158795 10848 158811 10912
rect 158875 10848 158891 10912
rect 158955 10848 158971 10912
rect 159035 10848 159043 10912
rect 158723 9824 159043 10848
rect 158723 9760 158731 9824
rect 158795 9760 158811 9824
rect 158875 9760 158891 9824
rect 158955 9760 158971 9824
rect 159035 9760 159043 9824
rect 158723 8736 159043 9760
rect 158723 8672 158731 8736
rect 158795 8672 158811 8736
rect 158875 8672 158891 8736
rect 158955 8672 158971 8736
rect 159035 8672 159043 8736
rect 158723 7648 159043 8672
rect 158723 7584 158731 7648
rect 158795 7584 158811 7648
rect 158875 7584 158891 7648
rect 158955 7584 158971 7648
rect 159035 7584 159043 7648
rect 158723 6560 159043 7584
rect 158723 6496 158731 6560
rect 158795 6496 158811 6560
rect 158875 6496 158891 6560
rect 158955 6496 158971 6560
rect 159035 6496 159043 6560
rect 158723 5472 159043 6496
rect 158723 5408 158731 5472
rect 158795 5408 158811 5472
rect 158875 5408 158891 5472
rect 158955 5408 158971 5472
rect 159035 5408 159043 5472
rect 156827 5404 156893 5405
rect 156827 5340 156828 5404
rect 156892 5340 156893 5404
rect 156827 5339 156893 5340
rect 158723 4384 159043 5408
rect 158723 4320 158731 4384
rect 158795 4320 158811 4384
rect 158875 4320 158891 4384
rect 158955 4320 158971 4384
rect 159035 4320 159043 4384
rect 158723 3296 159043 4320
rect 158723 3232 158731 3296
rect 158795 3232 158811 3296
rect 158875 3232 158891 3296
rect 158955 3232 158971 3296
rect 159035 3232 159043 3296
rect 158723 2208 159043 3232
rect 158723 2144 158731 2208
rect 158795 2144 158811 2208
rect 158875 2144 158891 2208
rect 158955 2144 158971 2208
rect 159035 2144 159043 2208
rect 158723 2128 159043 2144
rect 155907 1324 155973 1325
rect 155907 1260 155908 1324
rect 155972 1260 155973 1324
rect 155907 1259 155973 1260
rect 124443 1188 124509 1189
rect 124443 1124 124444 1188
rect 124508 1124 124509 1188
rect 124443 1123 124509 1124
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__B
timestamp 1670771148
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1670771148
transform 1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1670771148
transform 1 0 12788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1670771148
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__B
timestamp 1670771148
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1670771148
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1670771148
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1670771148
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1670771148
transform 1 0 24748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1670771148
transform 1 0 23736 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1670771148
transform 1 0 21804 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1670771148
transform 1 0 25208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1670771148
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A
timestamp 1670771148
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__B
timestamp 1670771148
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1670771148
transform 1 0 8372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A
timestamp 1670771148
transform 1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__B
timestamp 1670771148
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1670771148
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1670771148
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1670771148
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__B
timestamp 1670771148
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1670771148
transform 1 0 5796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__B
timestamp 1670771148
transform 1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A
timestamp 1670771148
transform -1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B
timestamp 1670771148
transform -1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1670771148
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B
timestamp 1670771148
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A
timestamp 1670771148
transform 1 0 7636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B
timestamp 1670771148
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1670771148
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1670771148
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1670771148
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1670771148
transform -1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1670771148
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1670771148
transform -1 0 11040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1670771148
transform 1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1670771148
transform -1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__B
timestamp 1670771148
transform -1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1670771148
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1670771148
transform -1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A
timestamp 1670771148
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1670771148
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1670771148
transform 1 0 10672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A
timestamp 1670771148
transform -1 0 18768 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1670771148
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1670771148
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1670771148
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1670771148
transform -1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__B
timestamp 1670771148
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1670771148
transform 1 0 32384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1670771148
transform -1 0 54648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1670771148
transform 1 0 49680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 1670771148
transform 1 0 46368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1670771148
transform 1 0 49128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A
timestamp 1670771148
transform 1 0 45264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 1670771148
transform 1 0 37628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1670771148
transform 1 0 36432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1670771148
transform 1 0 37812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A
timestamp 1670771148
transform 1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B
timestamp 1670771148
transform 1 0 46184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A
timestamp 1670771148
transform 1 0 40848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A
timestamp 1670771148
transform 1 0 37628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1670771148
transform 1 0 100832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A
timestamp 1670771148
transform -1 0 64400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1670771148
transform 1 0 30084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1670771148
transform 1 0 34224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1670771148
transform 1 0 34132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__B
timestamp 1670771148
transform -1 0 35052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1670771148
transform 1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1670771148
transform 1 0 32384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__B
timestamp 1670771148
transform -1 0 32936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1670771148
transform 1 0 30360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1670771148
transform -1 0 33304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1670771148
transform -1 0 33856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1670771148
transform 1 0 31096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1670771148
transform -1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1670771148
transform 1 0 27232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1670771148
transform 1 0 34132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1670771148
transform -1 0 33672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 1670771148
transform 1 0 79396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1670771148
transform 1 0 38824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 1670771148
transform 1 0 38180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1670771148
transform 1 0 44344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1670771148
transform 1 0 48024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A
timestamp 1670771148
transform 1 0 45724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A
timestamp 1670771148
transform 1 0 37536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 1670771148
transform -1 0 37168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1670771148
transform -1 0 41216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1670771148
transform 1 0 47104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1670771148
transform -1 0 52440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B
timestamp 1670771148
transform 1 0 50876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1670771148
transform 1 0 45816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1670771148
transform -1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1670771148
transform 1 0 66608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1670771148
transform 1 0 46276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1670771148
transform 1 0 55476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B
timestamp 1670771148
transform 1 0 58696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1670771148
transform 1 0 41860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1670771148
transform -1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1670771148
transform 1 0 50416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1670771148
transform 1 0 47748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1670771148
transform -1 0 65780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1670771148
transform 1 0 65964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1670771148
transform 1 0 59708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1670771148
transform 1 0 52072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1670771148
transform 1 0 52624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1670771148
transform 1 0 52256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1670771148
transform -1 0 63388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1670771148
transform -1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1670771148
transform 1 0 59524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1670771148
transform 1 0 51428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1670771148
transform 1 0 59708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1670771148
transform 1 0 61272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1670771148
transform -1 0 58328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1670771148
transform 1 0 63296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1670771148
transform 1 0 65136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1670771148
transform 1 0 55476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1670771148
transform 1 0 54740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1670771148
transform 1 0 57592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1670771148
transform 1 0 65136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1670771148
transform -1 0 49864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A
timestamp 1670771148
transform 1 0 65136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B
timestamp 1670771148
transform 1 0 64492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1670771148
transform 1 0 66884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1670771148
transform 1 0 56856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1670771148
transform 1 0 59248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1670771148
transform 1 0 62468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1670771148
transform 1 0 69552 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1670771148
transform 1 0 71760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1670771148
transform 1 0 72864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1670771148
transform 1 0 67712 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1670771148
transform 1 0 72312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1670771148
transform 1 0 73968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B
timestamp 1670771148
transform 1 0 72588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1670771148
transform 1 0 73508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B
timestamp 1670771148
transform 1 0 73508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1670771148
transform 1 0 77648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1670771148
transform 1 0 81788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1670771148
transform 1 0 87216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1670771148
transform 1 0 81420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A
timestamp 1670771148
transform 1 0 76912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1670771148
transform 1 0 74244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1670771148
transform 1 0 83076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1670771148
transform 1 0 83720 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1670771148
transform 1 0 93012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1670771148
transform 1 0 86388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1670771148
transform 1 0 107180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1670771148
transform 1 0 106996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1670771148
transform 1 0 98532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B
timestamp 1670771148
transform 1 0 97796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1670771148
transform 1 0 82064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 1670771148
transform -1 0 82800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1670771148
transform 1 0 107732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1670771148
transform -1 0 106536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A
timestamp 1670771148
transform -1 0 111412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B
timestamp 1670771148
transform -1 0 110860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1670771148
transform 1 0 99820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B
timestamp 1670771148
transform -1 0 100556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1670771148
transform 1 0 90804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1670771148
transform 1 0 91540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1670771148
transform -1 0 91908 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1670771148
transform 1 0 93932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1670771148
transform 1 0 112148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1670771148
transform -1 0 123188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1670771148
transform -1 0 122636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1670771148
transform 1 0 119600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 1670771148
transform -1 0 120612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1670771148
transform 1 0 115920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B
timestamp 1670771148
transform 1 0 115276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1670771148
transform 1 0 118772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B
timestamp 1670771148
transform 1 0 118220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1670771148
transform 1 0 120888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B
timestamp 1670771148
transform 1 0 120520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1670771148
transform 1 0 108560 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1670771148
transform -1 0 107732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1670771148
transform 1 0 116840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B
timestamp 1670771148
transform 1 0 117392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1670771148
transform -1 0 115736 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B
timestamp 1670771148
transform -1 0 114264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1670771148
transform 1 0 116196 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1670771148
transform -1 0 117484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1670771148
transform 1 0 113068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1670771148
transform 1 0 112700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1670771148
transform 1 0 116656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1670771148
transform 1 0 125856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1670771148
transform -1 0 125212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1670771148
transform 1 0 128248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B
timestamp 1670771148
transform -1 0 130916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1670771148
transform 1 0 114724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B
timestamp 1670771148
transform 1 0 113620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1670771148
transform 1 0 127604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B
timestamp 1670771148
transform -1 0 129444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1670771148
transform 1 0 131008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B
timestamp 1670771148
transform 1 0 129536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 1670771148
transform 1 0 114264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 1670771148
transform 1 0 113252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A
timestamp 1670771148
transform 1 0 133584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 1670771148
transform 1 0 132112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1670771148
transform 1 0 131376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B
timestamp 1670771148
transform -1 0 130364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1670771148
transform 1 0 132388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B
timestamp 1670771148
transform -1 0 131468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1670771148
transform -1 0 134320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B
timestamp 1670771148
transform -1 0 133768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A
timestamp 1670771148
transform -1 0 120060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A
timestamp 1670771148
transform -1 0 129628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B
timestamp 1670771148
transform -1 0 130364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1670771148
transform 1 0 126592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B
timestamp 1670771148
transform -1 0 127328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1670771148
transform -1 0 131744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B
timestamp 1670771148
transform -1 0 130364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1670771148
transform 1 0 124200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 1670771148
transform -1 0 123832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1670771148
transform 1 0 119232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B
timestamp 1670771148
transform -1 0 119784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1670771148
transform 1 0 127236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1670771148
transform -1 0 127788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1670771148
transform 1 0 127604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1670771148
transform -1 0 127328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1670771148
transform 1 0 123280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B
timestamp 1670771148
transform 1 0 121808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1670771148
transform 1 0 119876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B
timestamp 1670771148
transform 1 0 118588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1670771148
transform 1 0 126132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B
timestamp 1670771148
transform 1 0 125304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1670771148
transform 1 0 137264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1670771148
transform 1 0 131744 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B
timestamp 1670771148
transform -1 0 121440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B
timestamp 1670771148
transform 1 0 120152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1670771148
transform -1 0 138092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1670771148
transform -1 0 126040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1670771148
transform 1 0 124384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B
timestamp 1670771148
transform -1 0 126776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B
timestamp 1670771148
transform -1 0 123464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1670771148
transform 1 0 131192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1670771148
transform 1 0 135056 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1670771148
transform 1 0 125028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1670771148
transform -1 0 124568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1670771148
transform 1 0 130456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B
timestamp 1670771148
transform 1 0 128432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1670771148
transform 1 0 123832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1670771148
transform -1 0 130916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1670771148
transform -1 0 158424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B
timestamp 1670771148
transform -1 0 150236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1670771148
transform -1 0 117852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B
timestamp 1670771148
transform -1 0 116840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1670771148
transform 1 0 131376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1670771148
transform 1 0 131560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1670771148
transform 1 0 134688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1670771148
transform 1 0 134504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1670771148
transform 1 0 126960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1670771148
transform 1 0 126408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1670771148
transform 1 0 147568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1670771148
transform -1 0 145084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1670771148
transform 1 0 139380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B
timestamp 1670771148
transform 1 0 138000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1670771148
transform 1 0 132480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1670771148
transform -1 0 114908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1670771148
transform 1 0 119876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1670771148
transform 1 0 121256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1670771148
transform 1 0 123556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1670771148
transform -1 0 120152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B
timestamp 1670771148
transform -1 0 121256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1670771148
transform -1 0 124016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1670771148
transform 1 0 126408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1670771148
transform 1 0 129628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1670771148
transform -1 0 124844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1670771148
transform 1 0 118128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1670771148
transform -1 0 120888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1670771148
transform 1 0 126040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B
timestamp 1670771148
transform 1 0 129536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1670771148
transform 1 0 137264 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1670771148
transform 1 0 131376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1670771148
transform -1 0 128156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1670771148
transform 1 0 128708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B
timestamp 1670771148
transform -1 0 128708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1670771148
transform 1 0 125764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1670771148
transform 1 0 126684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1670771148
transform 1 0 131008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1670771148
transform 1 0 137632 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1670771148
transform -1 0 118864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B
timestamp 1670771148
transform -1 0 123740 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1670771148
transform 1 0 126408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B
timestamp 1670771148
transform -1 0 129168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1670771148
transform 1 0 126408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1670771148
transform 1 0 122452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1670771148
transform 1 0 123004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1670771148
transform 1 0 136344 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1670771148
transform 1 0 120152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1670771148
transform -1 0 116840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1670771148
transform -1 0 152352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1670771148
transform 1 0 122176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1670771148
transform -1 0 126592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1670771148
transform 1 0 121624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1670771148
transform 1 0 125488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B
timestamp 1670771148
transform -1 0 128064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1670771148
transform 1 0 136252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1670771148
transform 1 0 139840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1670771148
transform 1 0 132848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B
timestamp 1670771148
transform -1 0 132296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1670771148
transform 1 0 139840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1670771148
transform -1 0 157412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1670771148
transform 1 0 126960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B
timestamp 1670771148
transform 1 0 125304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1670771148
transform 1 0 124384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1670771148
transform 1 0 128984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1670771148
transform -1 0 116472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1670771148
transform -1 0 126040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1670771148
transform 1 0 139748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B
timestamp 1670771148
transform 1 0 139196 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1670771148
transform 1 0 150144 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1670771148
transform 1 0 120520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1670771148
transform -1 0 121992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1670771148
transform 1 0 133032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1670771148
transform 1 0 120796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__B
timestamp 1670771148
transform -1 0 121992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1670771148
transform -1 0 122912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1670771148
transform 1 0 124108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1670771148
transform 1 0 131928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1670771148
transform 1 0 132296 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1670771148
transform 1 0 125212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1670771148
transform 1 0 121348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1670771148
transform -1 0 122084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1670771148
transform 1 0 123188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1670771148
transform -1 0 136896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B
timestamp 1670771148
transform -1 0 137448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1670771148
transform 1 0 139840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1670771148
transform -1 0 138644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1670771148
transform -1 0 115920 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B
timestamp 1670771148
transform -1 0 124568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1670771148
transform -1 0 124660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1670771148
transform 1 0 132112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1670771148
transform 1 0 130272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1670771148
transform -1 0 132112 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B
timestamp 1670771148
transform 1 0 130824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1670771148
transform -1 0 124568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1670771148
transform -1 0 124016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B
timestamp 1670771148
transform -1 0 134136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 1670771148
transform -1 0 127880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B
timestamp 1670771148
transform -1 0 125488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1670771148
transform -1 0 120888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1670771148
transform -1 0 131744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1670771148
transform -1 0 120888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B
timestamp 1670771148
transform -1 0 127144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1670771148
transform -1 0 117668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B
timestamp 1670771148
transform -1 0 118864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1670771148
transform 1 0 134136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B
timestamp 1670771148
transform -1 0 134872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1670771148
transform 1 0 138644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1670771148
transform 1 0 139840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B
timestamp 1670771148
transform 1 0 140484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1670771148
transform 1 0 139840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1670771148
transform 1 0 140852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B
timestamp 1670771148
transform 1 0 139012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1670771148
transform 1 0 134136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1670771148
transform 1 0 134688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1670771148
transform 1 0 124384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1670771148
transform 1 0 130824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1670771148
transform -1 0 127144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1670771148
transform -1 0 140484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1670771148
transform 1 0 127880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1670771148
transform 1 0 111320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1670771148
transform 1 0 110768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1670771148
transform 1 0 110492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1670771148
transform 1 0 115368 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1670771148
transform 1 0 114724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B
timestamp 1670771148
transform 1 0 113068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1670771148
transform 1 0 112608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1670771148
transform -1 0 112240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1670771148
transform 1 0 104880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1670771148
transform -1 0 104420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1670771148
transform 1 0 113896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1670771148
transform 1 0 112700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1670771148
transform 1 0 109572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1670771148
transform -1 0 109756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1670771148
transform -1 0 107180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1670771148
transform -1 0 103960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1670771148
transform 1 0 61180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1670771148
transform 1 0 96600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1670771148
transform -1 0 113344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B
timestamp 1670771148
transform 1 0 112700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1670771148
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1670771148
transform 1 0 30820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1670771148
transform -1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A
timestamp 1670771148
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A
timestamp 1670771148
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B
timestamp 1670771148
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1670771148
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1670771148
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1670771148
transform 1 0 9844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A
timestamp 1670771148
transform -1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1670771148
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1670771148
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1670771148
transform 1 0 17572 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B
timestamp 1670771148
transform 1 0 18216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1670771148
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1670771148
transform -1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1670771148
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1670771148
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B
timestamp 1670771148
transform -1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__CLK
timestamp 1670771148
transform 1 0 21252 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__CLK
timestamp 1670771148
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__CLK
timestamp 1670771148
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__CLK
timestamp 1670771148
transform 1 0 23736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__CLK
timestamp 1670771148
transform 1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__CLK
timestamp 1670771148
transform 1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1670771148
transform 1 0 28980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__CLK
timestamp 1670771148
transform 1 0 21988 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1670771148
transform 1 0 23920 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1670771148
transform 1 0 26404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__CLK
timestamp 1670771148
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1670771148
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__CLK
timestamp 1670771148
transform 1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1670771148
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1670771148
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1670771148
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1670771148
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1670771148
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1670771148
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1670771148
transform -1 0 15180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1670771148
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1670771148
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1670771148
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1670771148
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1670771148
transform 1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1670771148
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1670771148
transform 1 0 26404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__CLK
timestamp 1670771148
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__CLK
timestamp 1670771148
transform 1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__CLK
timestamp 1670771148
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__CLK
timestamp 1670771148
transform -1 0 50508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__D
timestamp 1670771148
transform -1 0 48208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1670771148
transform -1 0 46828 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__CLK
timestamp 1670771148
transform 1 0 40664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__CLK
timestamp 1670771148
transform 1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__CLK
timestamp 1670771148
transform 1 0 48576 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1670771148
transform 1 0 39376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__CLK
timestamp 1670771148
transform 1 0 56120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__CLK
timestamp 1670771148
transform 1 0 35696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1670771148
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__CLK
timestamp 1670771148
transform 1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1670771148
transform 1 0 34776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1670771148
transform -1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1670771148
transform 1 0 38456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1670771148
transform -1 0 38640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__CLK
timestamp 1670771148
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1670771148
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__CLK
timestamp 1670771148
transform 1 0 30084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__CLK
timestamp 1670771148
transform 1 0 27232 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1670771148
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__CLK
timestamp 1670771148
transform 1 0 31004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__CLK
timestamp 1670771148
transform 1 0 37904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__CLK
timestamp 1670771148
transform -1 0 37904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__CLK
timestamp 1670771148
transform 1 0 42228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__CLK
timestamp 1670771148
transform 1 0 39928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1670771148
transform 1 0 40020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__CLK
timestamp 1670771148
transform -1 0 45264 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1670771148
transform 1 0 32200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__CLK
timestamp 1670771148
transform 1 0 45264 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1670771148
transform 1 0 47104 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__CLK
timestamp 1670771148
transform 1 0 54648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1670771148
transform 1 0 39376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1670771148
transform 1 0 39376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1670771148
transform -1 0 48024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1670771148
transform 1 0 39560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1670771148
transform -1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1670771148
transform 1 0 55568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1670771148
transform 1 0 65780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1670771148
transform 1 0 62192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1670771148
transform 1 0 58972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1670771148
transform 1 0 38732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1670771148
transform 1 0 65504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1670771148
transform 1 0 65228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1670771148
transform -1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1670771148
transform 1 0 44436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1670771148
transform -1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1670771148
transform 1 0 49680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1670771148
transform 1 0 74336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1670771148
transform 1 0 65780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1670771148
transform 1 0 53360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1670771148
transform -1 0 51704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1670771148
transform 1 0 55752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1670771148
transform 1 0 60628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1670771148
transform 1 0 66608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1670771148
transform 1 0 62560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1670771148
transform 1 0 55936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1670771148
transform 1 0 63204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1670771148
transform 1 0 62100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1670771148
transform 1 0 66976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1670771148
transform 1 0 78016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1670771148
transform 1 0 73784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1670771148
transform 1 0 65780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1670771148
transform 1 0 93196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__D
timestamp 1670771148
transform -1 0 94300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1670771148
transform -1 0 66240 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1670771148
transform 1 0 72036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1670771148
transform 1 0 87308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1670771148
transform 1 0 93748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1670771148
transform 1 0 74888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1670771148
transform 1 0 76084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1670771148
transform 1 0 88320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1670771148
transform 1 0 88228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1670771148
transform 1 0 80592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1670771148
transform 1 0 76728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1670771148
transform 1 0 96140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__D
timestamp 1670771148
transform 1 0 96692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1670771148
transform 1 0 81236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__D
timestamp 1670771148
transform 1 0 82892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1670771148
transform 1 0 81236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1670771148
transform 1 0 85744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1670771148
transform 1 0 88228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1670771148
transform 1 0 93196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__D
timestamp 1670771148
transform 1 0 92644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1670771148
transform 1 0 97244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1670771148
transform 1 0 101200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1670771148
transform 1 0 93380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1670771148
transform 1 0 77188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__D
timestamp 1670771148
transform 1 0 79764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1670771148
transform 1 0 75900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__D
timestamp 1670771148
transform -1 0 76636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1670771148
transform 1 0 114724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1670771148
transform 1 0 108836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1670771148
transform 1 0 97796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__D
timestamp 1670771148
transform -1 0 98348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1670771148
transform 1 0 74336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__D
timestamp 1670771148
transform -1 0 77372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1670771148
transform 1 0 88780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__D
timestamp 1670771148
transform -1 0 91080 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1670771148
transform 1 0 112884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1670771148
transform 1 0 117392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1670771148
transform 1 0 90712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__D
timestamp 1670771148
transform -1 0 92920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1670771148
transform 1 0 117300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__CLK
timestamp 1670771148
transform 1 0 104236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__D
timestamp 1670771148
transform 1 0 103316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1670771148
transform 1 0 101200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__D
timestamp 1670771148
transform 1 0 100648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__CLK
timestamp 1670771148
transform 1 0 100556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1670771148
transform 1 0 123648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__CLK
timestamp 1670771148
transform 1 0 104420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1670771148
transform -1 0 106628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1670771148
transform 1 0 102488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1670771148
transform 1 0 107548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__D
timestamp 1670771148
transform 1 0 106996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1670771148
transform 1 0 76636 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__D
timestamp 1670771148
transform 1 0 76268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1670771148
transform 1 0 104420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__D
timestamp 1670771148
transform 1 0 103408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1670771148
transform 1 0 99268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__D
timestamp 1670771148
transform 1 0 98256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1670771148
transform 1 0 99268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__D
timestamp 1670771148
transform 1 0 101844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1670771148
transform 1 0 94852 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__D
timestamp 1670771148
transform -1 0 94484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1670771148
transform 1 0 92184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__D
timestamp 1670771148
transform -1 0 94484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1670771148
transform 1 0 63664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__D
timestamp 1670771148
transform -1 0 62744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1670771148
transform 1 0 89700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__D
timestamp 1670771148
transform 1 0 88320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1670771148
transform 1 0 87676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__D
timestamp 1670771148
transform -1 0 87308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1670771148
transform 1 0 93472 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__D
timestamp 1670771148
transform -1 0 96416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1670771148
transform -1 0 73692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__D
timestamp 1670771148
transform -1 0 73048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1670771148
transform 1 0 96048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1670771148
transform -1 0 98716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1670771148
transform 1 0 134136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1670771148
transform 1 0 137908 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1670771148
transform 1 0 132112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1670771148
transform 1 0 147476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1670771148
transform -1 0 133768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1670771148
transform 1 0 122544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1670771148
transform 1 0 136804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__D
timestamp 1670771148
transform -1 0 137172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1670771148
transform 1 0 139656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__D
timestamp 1670771148
transform -1 0 139288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1670771148
transform 1 0 138460 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__D
timestamp 1670771148
transform -1 0 139472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__CLK
timestamp 1670771148
transform 1 0 135240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__CLK
timestamp 1670771148
transform 1 0 135608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1670771148
transform 1 0 137448 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1670771148
transform -1 0 151800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__CLK
timestamp 1670771148
transform 1 0 130180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1670771148
transform 1 0 134964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__CLK
timestamp 1670771148
transform 1 0 134136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1670771148
transform 1 0 117116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__D
timestamp 1670771148
transform 1 0 117300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__CLK
timestamp 1670771148
transform 1 0 125304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__D
timestamp 1670771148
transform -1 0 124936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1670771148
transform 1 0 110676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__D
timestamp 1670771148
transform -1 0 110308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__CLK
timestamp 1670771148
transform 1 0 119876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__D
timestamp 1670771148
transform 1 0 119232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__CLK
timestamp 1670771148
transform 1 0 110124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__D
timestamp 1670771148
transform -1 0 109756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__CLK
timestamp 1670771148
transform 1 0 117760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__CLK
timestamp 1670771148
transform 1 0 108836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__CLK
timestamp 1670771148
transform 1 0 121808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__CLK
timestamp 1670771148
transform 1 0 122452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__CLK
timestamp 1670771148
transform 1 0 135700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__D
timestamp 1670771148
transform -1 0 136160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__CLK
timestamp 1670771148
transform 1 0 137632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__CLK
timestamp 1670771148
transform 1 0 142416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__CLK
timestamp 1670771148
transform -1 0 158424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__CLK
timestamp 1670771148
transform 1 0 138092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__CLK
timestamp 1670771148
transform 1 0 141312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__D
timestamp 1670771148
transform -1 0 139472 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__CLK
timestamp 1670771148
transform 1 0 136528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1670771148
transform 1 0 129260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__D
timestamp 1670771148
transform -1 0 129260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__CLK
timestamp 1670771148
transform -1 0 110400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__CLK
timestamp 1670771148
transform 1 0 119232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1670771148
transform 1 0 134688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__CLK
timestamp 1670771148
transform 1 0 133584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__CLK
timestamp 1670771148
transform 1 0 147016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__CLK
timestamp 1670771148
transform 1 0 137080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__CLK
timestamp 1670771148
transform 1 0 140484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__D
timestamp 1670771148
transform -1 0 136528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1670771148
transform 1 0 152720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__D
timestamp 1670771148
transform -1 0 131744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__CLK
timestamp 1670771148
transform 1 0 136712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__CLK
timestamp 1670771148
transform 1 0 136896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__CLK
timestamp 1670771148
transform -1 0 158424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__CLK
timestamp 1670771148
transform 1 0 128984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__D
timestamp 1670771148
transform -1 0 128616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__CLK
timestamp 1670771148
transform 1 0 147568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__CLK
timestamp 1670771148
transform -1 0 158424 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__D
timestamp 1670771148
transform -1 0 158056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__CLK
timestamp 1670771148
transform 1 0 141864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__CLK
timestamp 1670771148
transform -1 0 147752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__CLK
timestamp 1670771148
transform 1 0 133124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__CLK
timestamp 1670771148
transform 1 0 152720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__CLK
timestamp 1670771148
transform 1 0 134688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__CLK
timestamp 1670771148
transform 1 0 133676 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__CLK
timestamp 1670771148
transform -1 0 152904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__CLK
timestamp 1670771148
transform 1 0 135608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__CLK
timestamp 1670771148
transform 1 0 135056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__CLK
timestamp 1670771148
transform 1 0 135700 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__CLK
timestamp 1670771148
transform -1 0 143244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__CLK
timestamp 1670771148
transform 1 0 142416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__CLK
timestamp 1670771148
transform 1 0 155296 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__CLK
timestamp 1670771148
transform 1 0 134228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__D
timestamp 1670771148
transform -1 0 136436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__CLK
timestamp 1670771148
transform 1 0 134136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__CLK
timestamp 1670771148
transform -1 0 150328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 1670771148
transform 1 0 134688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__CLK
timestamp 1670771148
transform 1 0 138184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__CLK
timestamp 1670771148
transform 1 0 150052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__CLK
timestamp 1670771148
transform 1 0 135792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__CLK
timestamp 1670771148
transform 1 0 121256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__CLK
timestamp 1670771148
transform 1 0 129720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__CLK
timestamp 1670771148
transform 1 0 124292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 1670771148
transform 1 0 133032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 1670771148
transform -1 0 142600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__CLK
timestamp 1670771148
transform 1 0 136804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 1670771148
transform 1 0 132112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__CLK
timestamp 1670771148
transform 1 0 127880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 1670771148
transform 1 0 136252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 1670771148
transform 1 0 155296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__CLK
timestamp 1670771148
transform 1 0 152720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__CLK
timestamp 1670771148
transform 1 0 148212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__CLK
timestamp 1670771148
transform -1 0 155480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__CLK
timestamp 1670771148
transform 1 0 136252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__CLK
timestamp 1670771148
transform 1 0 135792 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__CLK
timestamp 1670771148
transform 1 0 137264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 1670771148
transform 1 0 133400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 1670771148
transform 1 0 137172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 1670771148
transform 1 0 137908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 1670771148
transform 1 0 139196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__CLK
timestamp 1670771148
transform 1 0 137908 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 1670771148
transform 1 0 155296 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 1670771148
transform 1 0 137908 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__CLK
timestamp 1670771148
transform 1 0 131836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__D
timestamp 1670771148
transform 1 0 131284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__CLK
timestamp 1670771148
transform 1 0 106996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__D
timestamp 1670771148
transform -1 0 107088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__CLK
timestamp 1670771148
transform 1 0 109572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__CLK
timestamp 1670771148
transform 1 0 115552 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__CLK
timestamp 1670771148
transform 1 0 112792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__CLK
timestamp 1670771148
transform 1 0 112424 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__CLK
timestamp 1670771148
transform -1 0 95036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__CLK
timestamp 1670771148
transform 1 0 109572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 1670771148
transform 1 0 111412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__CLK
timestamp 1670771148
transform 1 0 96508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__CLK
timestamp 1670771148
transform 1 0 102672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__CLK
timestamp 1670771148
transform 1 0 78844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__CLK
timestamp 1670771148
transform 1 0 101200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__CLK
timestamp 1670771148
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__D
timestamp 1670771148
transform -1 0 28980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__CLK
timestamp 1670771148
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__CLK
timestamp 1670771148
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__CLK
timestamp 1670771148
transform 1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1670771148
transform -1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__D
timestamp 1670771148
transform 1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__D
timestamp 1670771148
transform 1 0 32752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__D
timestamp 1670771148
transform -1 0 29900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__D
timestamp 1670771148
transform -1 0 33028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__D
timestamp 1670771148
transform 1 0 32660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1670771148
transform 1 0 21160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__D
timestamp 1670771148
transform 1 0 35420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__D
timestamp 1670771148
transform -1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__D
timestamp 1670771148
transform -1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__D
timestamp 1670771148
transform -1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__D
timestamp 1670771148
transform -1 0 37996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__D
timestamp 1670771148
transform 1 0 28520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__D
timestamp 1670771148
transform -1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1670771148
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__D
timestamp 1670771148
transform -1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__D
timestamp 1670771148
transform -1 0 35052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__D
timestamp 1670771148
transform -1 0 49588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__D
timestamp 1670771148
transform 1 0 34960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__D
timestamp 1670771148
transform 1 0 50416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__D
timestamp 1670771148
transform -1 0 40296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__D
timestamp 1670771148
transform 1 0 44528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1670771148
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1670771148
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1670771148
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1670771148
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1670771148
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__D
timestamp 1670771148
transform 1 0 30544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__D
timestamp 1670771148
transform -1 0 32476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__D
timestamp 1670771148
transform 1 0 47288 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__D
timestamp 1670771148
transform 1 0 56304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__D
timestamp 1670771148
transform -1 0 44620 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__D
timestamp 1670771148
transform 1 0 44068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__D
timestamp 1670771148
transform -1 0 36984 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__D
timestamp 1670771148
transform -1 0 48760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__D
timestamp 1670771148
transform -1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1670771148
transform 1 0 62928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__D
timestamp 1670771148
transform -1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__D
timestamp 1670771148
transform -1 0 60076 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1670771148
transform 1 0 72772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__D
timestamp 1670771148
transform 1 0 72588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__D
timestamp 1670771148
transform -1 0 74796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1670771148
transform 1 0 68356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1670771148
transform 1 0 68356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__D
timestamp 1670771148
transform -1 0 65872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__D
timestamp 1670771148
transform -1 0 53360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__D
timestamp 1670771148
transform -1 0 52900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1670771148
transform 1 0 63572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__D
timestamp 1670771148
transform -1 0 53176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__D
timestamp 1670771148
transform 1 0 77924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1670771148
transform 1 0 66516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1670771148
transform 1 0 73600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1670771148
transform 1 0 68356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__D
timestamp 1670771148
transform 1 0 78844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__D
timestamp 1670771148
transform 1 0 83076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__D
timestamp 1670771148
transform -1 0 90988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__D
timestamp 1670771148
transform 1 0 81880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__D
timestamp 1670771148
transform 1 0 85928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__D
timestamp 1670771148
transform -1 0 77004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1670771148
transform 1 0 72864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__D
timestamp 1670771148
transform -1 0 73600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1670771148
transform 1 0 88412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__D
timestamp 1670771148
transform -1 0 89148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1670771148
transform 1 0 73140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__D
timestamp 1670771148
transform 1 0 74612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__D
timestamp 1670771148
transform 1 0 80960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1670771148
transform 1 0 85652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__D
timestamp 1670771148
transform -1 0 88228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1670771148
transform 1 0 70288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__D
timestamp 1670771148
transform 1 0 72312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1670771148
transform 1 0 78752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__D
timestamp 1670771148
transform 1 0 79120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1670771148
transform 1 0 69276 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__D
timestamp 1670771148
transform -1 0 71852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1670771148
transform 1 0 83168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__D
timestamp 1670771148
transform 1 0 85652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__D
timestamp 1670771148
transform -1 0 50600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__D
timestamp 1670771148
transform 1 0 90252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1670771148
transform 1 0 68356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__D
timestamp 1670771148
transform 1 0 70196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__D
timestamp 1670771148
transform 1 0 93380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__D
timestamp 1670771148
transform -1 0 91724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__D
timestamp 1670771148
transform 1 0 96692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__D
timestamp 1670771148
transform 1 0 61548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__D
timestamp 1670771148
transform 1 0 87952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1670771148
transform 1 0 71300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__D
timestamp 1670771148
transform 1 0 72864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1670771148
transform 1 0 69092 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__D
timestamp 1670771148
transform 1 0 71116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__D
timestamp 1670771148
transform 1 0 60720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__D
timestamp 1670771148
transform 1 0 90344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__D
timestamp 1670771148
transform -1 0 60076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1670771148
transform 1 0 80500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__D
timestamp 1670771148
transform 1 0 83168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__D
timestamp 1670771148
transform 1 0 88228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__D
timestamp 1670771148
transform -1 0 61732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__D
timestamp 1670771148
transform 1 0 65044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__D
timestamp 1670771148
transform -1 0 110308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1670771148
transform 1 0 68172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__D
timestamp 1670771148
transform 1 0 71024 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__D
timestamp 1670771148
transform -1 0 60812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__D
timestamp 1670771148
transform 1 0 59524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1670771148
transform 1 0 96048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__D
timestamp 1670771148
transform 1 0 98164 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1670771148
transform 1 0 140484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__D
timestamp 1670771148
transform 1 0 141036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1670771148
transform -1 0 152904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__D
timestamp 1670771148
transform 1 0 110308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1670771148
transform 1 0 95956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__D
timestamp 1670771148
transform 1 0 98348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__D
timestamp 1670771148
transform 1 0 92644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK
timestamp 1670771148
transform 1 0 76544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__D
timestamp 1670771148
transform 1 0 77740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__D
timestamp 1670771148
transform 1 0 93380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__D
timestamp 1670771148
transform 1 0 124108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1670771148
transform 1 0 97796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__D
timestamp 1670771148
transform 1 0 100188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__D
timestamp 1670771148
transform 1 0 125304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__D
timestamp 1670771148
transform 1 0 119232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__D
timestamp 1670771148
transform -1 0 123740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__D
timestamp 1670771148
transform 1 0 123004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1670771148
transform 1 0 88964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1670771148
transform 1 0 91356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__D
timestamp 1670771148
transform -1 0 126960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__D
timestamp 1670771148
transform 1 0 82984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1670771148
transform 1 0 95404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__D
timestamp 1670771148
transform -1 0 117024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__D
timestamp 1670771148
transform -1 0 130364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__D
timestamp 1670771148
transform 1 0 126960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__D
timestamp 1670771148
transform -1 0 126868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__D
timestamp 1670771148
transform -1 0 158056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__D
timestamp 1670771148
transform 1 0 109940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__D
timestamp 1670771148
transform 1 0 116564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__D
timestamp 1670771148
transform 1 0 111412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__D
timestamp 1670771148
transform 1 0 108192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__D
timestamp 1670771148
transform 1 0 137172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__CLK
timestamp 1670771148
transform -1 0 135884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__D
timestamp 1670771148
transform -1 0 136344 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__D
timestamp 1670771148
transform -1 0 123464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__CLK
timestamp 1670771148
transform 1 0 137356 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__D
timestamp 1670771148
transform 1 0 130824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__CLK
timestamp 1670771148
transform 1 0 141864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__CLK
timestamp 1670771148
transform 1 0 136344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__D
timestamp 1670771148
transform 1 0 127880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__CLK
timestamp 1670771148
transform 1 0 136068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__CLK
timestamp 1670771148
transform 1 0 139288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__CLK
timestamp 1670771148
transform -1 0 122912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1542__D
timestamp 1670771148
transform 1 0 136896 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__D
timestamp 1670771148
transform -1 0 133032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__D
timestamp 1670771148
transform 1 0 125948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__D
timestamp 1670771148
transform 1 0 123832 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1670771148
transform 1 0 126684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__D
timestamp 1670771148
transform 1 0 125028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__D
timestamp 1670771148
transform 1 0 118772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__D
timestamp 1670771148
transform 1 0 121624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__D
timestamp 1670771148
transform 1 0 131100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__D
timestamp 1670771148
transform 1 0 106444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__D
timestamp 1670771148
transform 1 0 127328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1553__D
timestamp 1670771148
transform -1 0 123832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__D
timestamp 1670771148
transform 1 0 115368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__D
timestamp 1670771148
transform 1 0 138736 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__D
timestamp 1670771148
transform 1 0 120704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__CLK
timestamp 1670771148
transform 1 0 140300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__D
timestamp 1670771148
transform 1 0 139840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__D
timestamp 1670771148
transform -1 0 127144 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__D
timestamp 1670771148
transform 1 0 123556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__CLK
timestamp 1670771148
transform 1 0 119876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__D
timestamp 1670771148
transform 1 0 120152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__D
timestamp 1670771148
transform -1 0 137172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__D
timestamp 1670771148
transform 1 0 129536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__D
timestamp 1670771148
transform 1 0 133124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__D
timestamp 1670771148
transform 1 0 131008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1571__D
timestamp 1670771148
transform -1 0 133860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__CLK
timestamp 1670771148
transform 1 0 139748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__D
timestamp 1670771148
transform 1 0 137356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__D
timestamp 1670771148
transform 1 0 128616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__D
timestamp 1670771148
transform -1 0 130364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__D
timestamp 1670771148
transform 1 0 133124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__D
timestamp 1670771148
transform -1 0 133676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__CLK
timestamp 1670771148
transform 1 0 138000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__D
timestamp 1670771148
transform 1 0 138368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__CLK
timestamp 1670771148
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__CLK
timestamp 1670771148
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__CLK
timestamp 1670771148
transform 1 0 17756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__CLK
timestamp 1670771148
transform 1 0 21252 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__CLK
timestamp 1670771148
transform 1 0 19412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__CLK
timestamp 1670771148
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__CLK
timestamp 1670771148
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__CLK
timestamp 1670771148
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__CLK
timestamp 1670771148
transform 1 0 22724 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__CLK
timestamp 1670771148
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__CLK
timestamp 1670771148
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__CLK
timestamp 1670771148
transform -1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__CLK
timestamp 1670771148
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_sclk_A
timestamp 1670771148
transform 1 0 80592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_sclk_A
timestamp 1670771148
transform 1 0 38088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_sclk_A
timestamp 1670771148
transform 1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_sclk_A
timestamp 1670771148
transform 1 0 68540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_sclk_A
timestamp 1670771148
transform 1 0 112148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_sclk_A
timestamp 1670771148
transform -1 0 144992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_sclk_A
timestamp 1670771148
transform 1 0 121624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_sclk_A
timestamp 1670771148
transform 1 0 138736 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_sclk_A
timestamp 1670771148
transform -1 0 132296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_sclk_A
timestamp 1670771148
transform 1 0 76176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_sclk_A
timestamp 1670771148
transform -1 0 27324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_sclk_A
timestamp 1670771148
transform 1 0 66056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout261_A
timestamp 1670771148
transform -1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout263_A
timestamp 1670771148
transform 1 0 24840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout265_A
timestamp 1670771148
transform -1 0 31096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout266_A
timestamp 1670771148
transform -1 0 40296 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout267_A
timestamp 1670771148
transform 1 0 38824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout268_A
timestamp 1670771148
transform 1 0 12512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout271_A
timestamp 1670771148
transform -1 0 45632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout273_A
timestamp 1670771148
transform 1 0 55660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout274_A
timestamp 1670771148
transform -1 0 67436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout275_A
timestamp 1670771148
transform 1 0 73784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout276_A
timestamp 1670771148
transform -1 0 69000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout277_A
timestamp 1670771148
transform -1 0 48392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout279_A
timestamp 1670771148
transform 1 0 84824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout280_A
timestamp 1670771148
transform 1 0 86388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout281_A
timestamp 1670771148
transform 1 0 119140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout282_A
timestamp 1670771148
transform 1 0 103684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout284_A
timestamp 1670771148
transform 1 0 125028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout285_A
timestamp 1670771148
transform -1 0 129444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout286_A
timestamp 1670771148
transform 1 0 130732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout287_A
timestamp 1670771148
transform 1 0 138644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout288_A
timestamp 1670771148
transform 1 0 132480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout290_A
timestamp 1670771148
transform -1 0 152904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout291_A
timestamp 1670771148
transform -1 0 139472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout292_A
timestamp 1670771148
transform -1 0 85008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1670771148
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1670771148
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1670771148
transform -1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_A
timestamp 1670771148
transform -1 0 66148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1670771148
transform -1 0 67804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output13_A
timestamp 1670771148
transform -1 0 67252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output15_A
timestamp 1670771148
transform -1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output17_A
timestamp 1670771148
transform 1 0 70932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output18_A
timestamp 1670771148
transform 1 0 71576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1670771148
transform 1 0 79948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1670771148
transform -1 0 9936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1670771148
transform -1 0 84732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1670771148
transform -1 0 84456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1670771148
transform -1 0 87308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1670771148
transform -1 0 89884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1670771148
transform -1 0 95036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1670771148
transform -1 0 96324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1670771148
transform -1 0 97428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1670771148
transform -1 0 95772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1670771148
transform -1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1670771148
transform -1 0 95588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1670771148
transform -1 0 98900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1670771148
transform 1 0 99268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1670771148
transform 1 0 95956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1670771148
transform 1 0 99820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1670771148
transform -1 0 99452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1670771148
transform -1 0 100004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1670771148
transform 1 0 101844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1670771148
transform 1 0 101200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1670771148
transform 1 0 103776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1670771148
transform 1 0 106904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1670771148
transform 1 0 103408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1670771148
transform 1 0 105616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1670771148
transform -1 0 106352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1670771148
transform 1 0 108928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1670771148
transform -1 0 104972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1670771148
transform 1 0 108560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1670771148
transform 1 0 109940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1670771148
transform 1 0 113436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1670771148
transform 1 0 113252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1670771148
transform 1 0 114540 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1670771148
transform -1 0 114172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1670771148
transform 1 0 112976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1670771148
transform 1 0 114724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1670771148
transform 1 0 115644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1670771148
transform -1 0 118036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1670771148
transform -1 0 119140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1670771148
transform -1 0 124476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1670771148
transform 1 0 119876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1670771148
transform 1 0 123096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1670771148
transform 1 0 125028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1670771148
transform 1 0 126132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1670771148
transform 1 0 125580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1670771148
transform 1 0 123096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1670771148
transform 1 0 125580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1670771148
transform 1 0 124384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1670771148
transform 1 0 129444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1670771148
transform -1 0 129076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1670771148
transform -1 0 128524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1670771148
transform 1 0 129996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1670771148
transform 1 0 130548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1670771148
transform 1 0 131652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output129_A
timestamp 1670771148
transform 1 0 131284 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1670771148
transform 1 0 131836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output134_A
timestamp 1670771148
transform 1 0 132756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1670771148
transform 1 0 133308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1670771148
transform -1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output143_A
timestamp 1670771148
transform -1 0 136252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1670771148
transform -1 0 135700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1670771148
transform -1 0 136252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1670771148
transform -1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1670771148
transform -1 0 138644 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1670771148
transform -1 0 143244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1670771148
transform -1 0 135700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output156_A
timestamp 1670771148
transform -1 0 136988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output157_A
timestamp 1670771148
transform 1 0 136252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output158_A
timestamp 1670771148
transform -1 0 136804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output163_A
timestamp 1670771148
transform -1 0 153548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1670771148
transform -1 0 157964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1670771148
transform -1 0 131192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1670771148
transform 1 0 125856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1670771148
transform -1 0 118404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1670771148
transform -1 0 115000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1670771148
transform -1 0 115368 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1670771148
transform -1 0 115552 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1670771148
transform 1 0 114080 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1670771148
transform -1 0 116288 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output177_A
timestamp 1670771148
transform 1 0 22908 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output182_A
timestamp 1670771148
transform -1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output183_A
timestamp 1670771148
transform -1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output185_A
timestamp 1670771148
transform -1 0 26128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output186_A
timestamp 1670771148
transform -1 0 26220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1670771148
transform -1 0 25576 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1670771148
transform -1 0 24840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output193_A
timestamp 1670771148
transform -1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output197_A
timestamp 1670771148
transform 1 0 33396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output201_A
timestamp 1670771148
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1670771148
transform -1 0 36432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1670771148
transform -1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1670771148
transform -1 0 42780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output228_A
timestamp 1670771148
transform -1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1670771148
transform -1 0 49312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output236_A
timestamp 1670771148
transform -1 0 53912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output237_A
timestamp 1670771148
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1670771148
transform -1 0 47288 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1670771148
transform 1 0 50600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1670771148
transform -1 0 10580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output259_A
timestamp 1670771148
transform -1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output260_A
timestamp 1670771148
transform -1 0 116840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1670771148
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1670771148
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1670771148
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61
timestamp 1670771148
transform 1 0 6716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1670771148
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1670771148
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1670771148
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1670771148
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1670771148
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122
timestamp 1670771148
transform 1 0 12328 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 13064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1670771148
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1670771148
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1670771148
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1670771148
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1670771148
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1670771148
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1670771148
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1670771148
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1670771148
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1670771148
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1670771148
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1670771148
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1670771148
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1670771148
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1670771148
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1670771148
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_271
timestamp 1670771148
transform 1 0 26036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1670771148
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1670771148
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1670771148
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1670771148
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1670771148
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1670771148
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_329
timestamp 1670771148
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1670771148
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_337
timestamp 1670771148
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1670771148
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1670771148
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1670771148
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1670771148
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1670771148
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1670771148
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1670771148
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1670771148
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1670771148
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1670771148
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1670771148
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_461
timestamp 1670771148
transform 1 0 43516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_469
timestamp 1670771148
transform 1 0 44252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1670771148
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1670771148
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1670771148
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_492
timestamp 1670771148
transform 1 0 46368 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1670771148
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1670771148
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1670771148
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1670771148
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1670771148
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1670771148
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1670771148
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1670771148
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1670771148
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1670771148
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1670771148
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1670771148
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1670771148
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 1670771148
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_625
timestamp 1670771148
transform 1 0 58604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1670771148
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 1670771148
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_649
timestamp 1670771148
transform 1 0 60812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_661
timestamp 1670771148
transform 1 0 61916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1670771148
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_673
timestamp 1670771148
transform 1 0 63020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_677
timestamp 1670771148
transform 1 0 63388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_694
timestamp 1670771148
transform 1 0 64952 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_701
timestamp 1670771148
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_705
timestamp 1670771148
transform 1 0 65964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_717
timestamp 1670771148
transform 1 0 67068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1670771148
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1670771148
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1670771148
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1670771148
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1670771148
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1670771148
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1670771148
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_785
timestamp 1670771148
transform 1 0 73324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_790
timestamp 1670771148
transform 1 0 73784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_810
timestamp 1670771148
transform 1 0 75624 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1670771148
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1670771148
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1670771148
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1670771148
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1670771148
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1670771148
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_869
timestamp 1670771148
transform 1 0 81052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_889
timestamp 1670771148
transform 1 0 82892 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 1670771148
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1670771148
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1670771148
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1670771148
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1670771148
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1670771148
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1670771148
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1670771148
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1670771148
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1670771148
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1670771148
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1670771148
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1670771148
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1670771148
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1670771148
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1670771148
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1670771148
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1670771148
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1670771148
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1670771148
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1670771148
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1670771148
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1670771148
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1670771148
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1670771148
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1670771148
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1670771148
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1670771148
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1149
timestamp 1670771148
transform 1 0 106812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1670771148
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1177
timestamp 1670771148
transform 1 0 109388 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1181
timestamp 1670771148
transform 1 0 109756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1193
timestamp 1670771148
transform 1 0 110860 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1670771148
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1670771148
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1219
timestamp 1670771148
transform 1 0 113252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1228
timestamp 1670771148
transform 1 0 114080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1233
timestamp 1670771148
transform 1 0 114540 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1237
timestamp 1670771148
transform 1 0 114908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1249
timestamp 1670771148
transform 1 0 116012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1670771148
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1261
timestamp 1670771148
transform 1 0 117116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1280
timestamp 1670771148
transform 1 0 118864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1286
timestamp 1670771148
transform 1 0 119416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1289
timestamp 1670771148
transform 1 0 119692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1293
timestamp 1670771148
transform 1 0 120060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1299
timestamp 1670771148
transform 1 0 120612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1302
timestamp 1670771148
transform 1 0 120888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1308
timestamp 1670771148
transform 1 0 121440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1314
timestamp 1670771148
transform 1 0 121992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1317
timestamp 1670771148
transform 1 0 122268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1321
timestamp 1670771148
transform 1 0 122636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1324
timestamp 1670771148
transform 1 0 122912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1330
timestamp 1670771148
transform 1 0 123464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1336
timestamp 1670771148
transform 1 0 124016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1342
timestamp 1670771148
transform 1 0 124568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1345
timestamp 1670771148
transform 1 0 124844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1349
timestamp 1670771148
transform 1 0 125212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1352
timestamp 1670771148
transform 1 0 125488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1358
timestamp 1670771148
transform 1 0 126040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1364
timestamp 1670771148
transform 1 0 126592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1370
timestamp 1670771148
transform 1 0 127144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1373
timestamp 1670771148
transform 1 0 127420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1377
timestamp 1670771148
transform 1 0 127788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1380
timestamp 1670771148
transform 1 0 128064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1386
timestamp 1670771148
transform 1 0 128616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1392
timestamp 1670771148
transform 1 0 129168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1398
timestamp 1670771148
transform 1 0 129720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1401
timestamp 1670771148
transform 1 0 129996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1408
timestamp 1670771148
transform 1 0 130640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1414
timestamp 1670771148
transform 1 0 131192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1420
timestamp 1670771148
transform 1 0 131744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1426
timestamp 1670771148
transform 1 0 132296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1429
timestamp 1670771148
transform 1 0 132572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1435
timestamp 1670771148
transform 1 0 133124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1452
timestamp 1670771148
transform 1 0 134688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1457
timestamp 1670771148
transform 1 0 135148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1475
timestamp 1670771148
transform 1 0 136804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1670771148
transform 1 0 137356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1485
timestamp 1670771148
transform 1 0 137724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1490
timestamp 1670771148
transform 1 0 138184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1499
timestamp 1670771148
transform 1 0 139012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1505
timestamp 1670771148
transform 1 0 139564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1511
timestamp 1670771148
transform 1 0 140116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1513
timestamp 1670771148
transform 1 0 140300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1532
timestamp 1670771148
transform 1 0 142048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1538
timestamp 1670771148
transform 1 0 142600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1541
timestamp 1670771148
transform 1 0 142876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1545
timestamp 1670771148
transform 1 0 143244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1566
timestamp 1670771148
transform 1 0 145176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1569
timestamp 1670771148
transform 1 0 145452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1587
timestamp 1670771148
transform 1 0 147108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1594
timestamp 1670771148
transform 1 0 147752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1597
timestamp 1670771148
transform 1 0 148028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1615
timestamp 1670771148
transform 1 0 149684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1670771148
transform 1 0 150236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1625
timestamp 1670771148
transform 1 0 150604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1632
timestamp 1670771148
transform 1 0 151248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1638
timestamp 1670771148
transform 1 0 151800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1644
timestamp 1670771148
transform 1 0 152352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1650
timestamp 1670771148
transform 1 0 152904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1653
timestamp 1670771148
transform 1 0 153180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1657
timestamp 1670771148
transform 1 0 153548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1668
timestamp 1670771148
transform 1 0 154560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1670771148
transform 1 0 155388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1681
timestamp 1670771148
transform 1 0 155756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1686
timestamp 1670771148
transform 1 0 156216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1693
timestamp 1670771148
transform 1 0 156860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1699
timestamp 1670771148
transform 1 0 157412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1670771148
transform 1 0 157964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1709
timestamp 1670771148
transform 1 0 158332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1670771148
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7
timestamp 1670771148
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1670771148
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1670771148
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_43
timestamp 1670771148
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_49
timestamp 1670771148
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1670771148
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1670771148
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1670771148
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1670771148
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1670771148
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp 1670771148
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1670771148
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1670771148
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1670771148
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1670771148
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1670771148
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1670771148
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 1670771148
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1670771148
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1670771148
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_180
timestamp 1670771148
transform 1 0 17664 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1670771148
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1670771148
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_212
timestamp 1670771148
transform 1 0 20608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1670771148
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1670771148
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1670771148
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_255
timestamp 1670771148
transform 1 0 24564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_267
timestamp 1670771148
transform 1 0 25668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1670771148
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1670771148
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1670771148
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_305
timestamp 1670771148
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_313
timestamp 1670771148
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1670771148
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1670771148
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_344
timestamp 1670771148
transform 1 0 32752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1670771148
transform 1 0 33304 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_356
timestamp 1670771148
transform 1 0 33856 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_368
timestamp 1670771148
transform 1 0 34960 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_380
timestamp 1670771148
transform 1 0 36064 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1670771148
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1670771148
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_417
timestamp 1670771148
transform 1 0 39468 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_423
timestamp 1670771148
transform 1 0 40020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1670771148
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1670771148
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1670771148
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_461
timestamp 1670771148
transform 1 0 43516 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_469
timestamp 1670771148
transform 1 0 44252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1670771148
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_493
timestamp 1670771148
transform 1 0 46460 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_499
timestamp 1670771148
transform 1 0 47012 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1670771148
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1670771148
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_523
timestamp 1670771148
transform 1 0 49220 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_543
timestamp 1670771148
transform 1 0 51060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1670771148
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1670771148
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1670771148
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1670771148
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_585
timestamp 1670771148
transform 1 0 54924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_591
timestamp 1670771148
transform 1 0 55476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_594
timestamp 1670771148
transform 1 0 55752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1670771148
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1670771148
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1670771148
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1670771148
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1670771148
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_665
timestamp 1670771148
transform 1 0 62284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_670
timestamp 1670771148
transform 1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_673
timestamp 1670771148
transform 1 0 63020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_691
timestamp 1670771148
transform 1 0 64676 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_699
timestamp 1670771148
transform 1 0 65412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_704
timestamp 1670771148
transform 1 0 65872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1670771148
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_729
timestamp 1670771148
transform 1 0 68172 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_733
timestamp 1670771148
transform 1 0 68540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_745
timestamp 1670771148
transform 1 0 69644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_757
timestamp 1670771148
transform 1 0 70748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_769
timestamp 1670771148
transform 1 0 71852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_777
timestamp 1670771148
transform 1 0 72588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_781
timestamp 1670771148
transform 1 0 72956 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1670771148
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1670771148
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1670771148
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1670771148
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1670771148
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1670771148
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1670771148
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1670771148
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_865
timestamp 1670771148
transform 1 0 80684 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_873
timestamp 1670771148
transform 1 0 81420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_885
timestamp 1670771148
transform 1 0 82524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_891
timestamp 1670771148
transform 1 0 83076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1670771148
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1670771148
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1670771148
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1670771148
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1670771148
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1670771148
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1670771148
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1670771148
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1670771148
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1670771148
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1670771148
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1670771148
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1670771148
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1670771148
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1670771148
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1035
timestamp 1670771148
transform 1 0 96324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1047
timestamp 1670771148
transform 1 0 97428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1059
timestamp 1670771148
transform 1 0 98532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1670771148
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1670771148
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1670771148
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1670771148
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1670771148
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1670771148
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1670771148
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1670771148
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1670771148
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1670771148
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1670771148
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1670771148
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1670771148
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1177
timestamp 1670771148
transform 1 0 109388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1181
timestamp 1670771148
transform 1 0 109756 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1187
timestamp 1670771148
transform 1 0 110308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1199
timestamp 1670771148
transform 1 0 111412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1211
timestamp 1670771148
transform 1 0 112516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1223
timestamp 1670771148
transform 1 0 113620 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1230
timestamp 1670771148
transform 1 0 114264 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1233
timestamp 1670771148
transform 1 0 114540 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1237
timestamp 1670771148
transform 1 0 114908 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1246
timestamp 1670771148
transform 1 0 115736 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1260
timestamp 1670771148
transform 1 0 117024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1264
timestamp 1670771148
transform 1 0 117392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1267
timestamp 1670771148
transform 1 0 117668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1274
timestamp 1670771148
transform 1 0 118312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1280
timestamp 1670771148
transform 1 0 118864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1286
timestamp 1670771148
transform 1 0 119416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1289
timestamp 1670771148
transform 1 0 119692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1294
timestamp 1670771148
transform 1 0 120152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1300
timestamp 1670771148
transform 1 0 120704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1306
timestamp 1670771148
transform 1 0 121256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1312
timestamp 1670771148
transform 1 0 121808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1318
timestamp 1670771148
transform 1 0 122360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1324
timestamp 1670771148
transform 1 0 122912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1330
timestamp 1670771148
transform 1 0 123464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1336
timestamp 1670771148
transform 1 0 124016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1342
timestamp 1670771148
transform 1 0 124568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1345
timestamp 1670771148
transform 1 0 124844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1349
timestamp 1670771148
transform 1 0 125212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1360
timestamp 1670771148
transform 1 0 126224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1364
timestamp 1670771148
transform 1 0 126592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1367
timestamp 1670771148
transform 1 0 126868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1374
timestamp 1670771148
transform 1 0 127512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1380
timestamp 1670771148
transform 1 0 128064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1384
timestamp 1670771148
transform 1 0 128432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1387
timestamp 1670771148
transform 1 0 128708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1393
timestamp 1670771148
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1670771148
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1401
timestamp 1670771148
transform 1 0 129996 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1405
timestamp 1670771148
transform 1 0 130364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1414
timestamp 1670771148
transform 1 0 131192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1438
timestamp 1670771148
transform 1 0 133400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1448
timestamp 1670771148
transform 1 0 134320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1454
timestamp 1670771148
transform 1 0 134872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1457
timestamp 1670771148
transform 1 0 135148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1476
timestamp 1670771148
transform 1 0 136896 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1496
timestamp 1670771148
transform 1 0 138736 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1504
timestamp 1670771148
transform 1 0 139472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1510
timestamp 1670771148
transform 1 0 140024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1513
timestamp 1670771148
transform 1 0 140300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1517
timestamp 1670771148
transform 1 0 140668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1523
timestamp 1670771148
transform 1 0 141220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1526
timestamp 1670771148
transform 1 0 141496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1532
timestamp 1670771148
transform 1 0 142048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1538
timestamp 1670771148
transform 1 0 142600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1545
timestamp 1670771148
transform 1 0 143244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1565
timestamp 1670771148
transform 1 0 145084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1569
timestamp 1670771148
transform 1 0 145452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1587
timestamp 1670771148
transform 1 0 147108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1607
timestamp 1670771148
transform 1 0 148948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1616
timestamp 1670771148
transform 1 0 149776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1622
timestamp 1670771148
transform 1 0 150328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1625
timestamp 1670771148
transform 1 0 150604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1632
timestamp 1670771148
transform 1 0 151248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1644
timestamp 1670771148
transform 1 0 152352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1650
timestamp 1670771148
transform 1 0 152904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1659
timestamp 1670771148
transform 1 0 153732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1663
timestamp 1670771148
transform 1 0 154100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1669
timestamp 1670771148
transform 1 0 154652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1678
timestamp 1670771148
transform 1 0 155480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1681
timestamp 1670771148
transform 1 0 155756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1687
timestamp 1670771148
transform 1 0 156308 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1691
timestamp 1670771148
transform 1 0 156676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1698
timestamp 1670771148
transform 1 0 157320 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1709
timestamp 1670771148
transform 1 0 158332 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1670771148
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1670771148
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1670771148
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1670771148
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1670771148
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1670771148
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1670771148
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1670771148
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1670771148
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1670771148
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1670771148
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1670771148
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_121
timestamp 1670771148
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1670771148
transform 1 0 12972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1670771148
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1670771148
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1670771148
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_148
timestamp 1670771148
transform 1 0 14720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1670771148
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_162
timestamp 1670771148
transform 1 0 16008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1670771148
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1670771148
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1670771148
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1670771148
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1670771148
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1670771148
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_225
timestamp 1670771148
transform 1 0 21804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1670771148
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1670771148
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1670771148
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1670771148
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_268
timestamp 1670771148
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_280
timestamp 1670771148
transform 1 0 26864 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_292
timestamp 1670771148
transform 1 0 27968 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1670771148
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1670771148
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_317
timestamp 1670771148
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1670771148
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1670771148
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1670771148
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1670771148
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1670771148
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_383
timestamp 1670771148
transform 1 0 36340 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_386
timestamp 1670771148
transform 1 0 36616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1670771148
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1670771148
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1670771148
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1670771148
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1670771148
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1670771148
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1670771148
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1670771148
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_469
timestamp 1670771148
transform 1 0 44252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1670771148
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1670771148
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_495
timestamp 1670771148
transform 1 0 46644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_507
timestamp 1670771148
transform 1 0 47748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_513
timestamp 1670771148
transform 1 0 48300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_530
timestamp 1670771148
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1670771148
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1670771148
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1670771148
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_569
timestamp 1670771148
transform 1 0 53452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_573
timestamp 1670771148
transform 1 0 53820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_585
timestamp 1670771148
transform 1 0 54924 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1670771148
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_601
timestamp 1670771148
transform 1 0 56396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_625
timestamp 1670771148
transform 1 0 58604 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_631
timestamp 1670771148
transform 1 0 59156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1670771148
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_645
timestamp 1670771148
transform 1 0 60444 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_655
timestamp 1670771148
transform 1 0 61364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_668
timestamp 1670771148
transform 1 0 62560 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_674
timestamp 1670771148
transform 1 0 63112 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_686
timestamp 1670771148
transform 1 0 64216 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_692
timestamp 1670771148
transform 1 0 64768 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_696
timestamp 1670771148
transform 1 0 65136 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1670771148
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1670771148
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1670771148
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1670771148
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1670771148
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1670771148
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1670771148
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_769
timestamp 1670771148
transform 1 0 71852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_779
timestamp 1670771148
transform 1 0 72772 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_799
timestamp 1670771148
transform 1 0 74612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1670771148
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_813
timestamp 1670771148
transform 1 0 75900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_831
timestamp 1670771148
transform 1 0 77556 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1670771148
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1670771148
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1670771148
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1670771148
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1670771148
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1670771148
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1670771148
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1670771148
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1670771148
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1670771148
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1670771148
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1670771148
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_951
timestamp 1670771148
transform 1 0 88596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_971
timestamp 1670771148
transform 1 0 90436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1670771148
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1670771148
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1670771148
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1005
timestamp 1670771148
transform 1 0 93564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1013
timestamp 1670771148
transform 1 0 94300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1031
timestamp 1670771148
transform 1 0 95956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1670771148
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1037
timestamp 1670771148
transform 1 0 96508 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1041
timestamp 1670771148
transform 1 0 96876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1053
timestamp 1670771148
transform 1 0 97980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1059
timestamp 1670771148
transform 1 0 98532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1077
timestamp 1670771148
transform 1 0 100188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1083
timestamp 1670771148
transform 1 0 100740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1670771148
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1093
timestamp 1670771148
transform 1 0 101660 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1111
timestamp 1670771148
transform 1 0 103316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1123
timestamp 1670771148
transform 1 0 104420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1135
timestamp 1670771148
transform 1 0 105524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1670771148
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1670771148
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1161
timestamp 1670771148
transform 1 0 107916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1181
timestamp 1670771148
transform 1 0 109756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1187
timestamp 1670771148
transform 1 0 110308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1193
timestamp 1670771148
transform 1 0 110860 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1201
timestamp 1670771148
transform 1 0 111596 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1670771148
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1670771148
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1670771148
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1241
timestamp 1670771148
transform 1 0 115276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1258
timestamp 1670771148
transform 1 0 116840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1261
timestamp 1670771148
transform 1 0 117116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1267
timestamp 1670771148
transform 1 0 117668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1284
timestamp 1670771148
transform 1 0 119232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1304
timestamp 1670771148
transform 1 0 121072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1314
timestamp 1670771148
transform 1 0 121992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1317
timestamp 1670771148
transform 1 0 122268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1321
timestamp 1670771148
transform 1 0 122636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1327
timestamp 1670771148
transform 1 0 123188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1333
timestamp 1670771148
transform 1 0 123740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1353
timestamp 1670771148
transform 1 0 125580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1359
timestamp 1670771148
transform 1 0 126132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1370
timestamp 1670771148
transform 1 0 127144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1373
timestamp 1670771148
transform 1 0 127420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1391
timestamp 1670771148
transform 1 0 129076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1411
timestamp 1670771148
transform 1 0 130916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1417
timestamp 1670771148
transform 1 0 131468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1423
timestamp 1670771148
transform 1 0 132020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1670771148
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1429
timestamp 1670771148
transform 1 0 132572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1436
timestamp 1670771148
transform 1 0 133216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1442
timestamp 1670771148
transform 1 0 133768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1448
timestamp 1670771148
transform 1 0 134320 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1454
timestamp 1670771148
transform 1 0 134872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1460
timestamp 1670771148
transform 1 0 135424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1466
timestamp 1670771148
transform 1 0 135976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1472
timestamp 1670771148
transform 1 0 136528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1478
timestamp 1670771148
transform 1 0 137080 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1485
timestamp 1670771148
transform 1 0 137724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1489
timestamp 1670771148
transform 1 0 138092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1509
timestamp 1670771148
transform 1 0 139932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1515
timestamp 1670771148
transform 1 0 140484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1521
timestamp 1670771148
transform 1 0 141036 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1529
timestamp 1670771148
transform 1 0 141772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1532
timestamp 1670771148
transform 1 0 142048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1538
timestamp 1670771148
transform 1 0 142600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1541
timestamp 1670771148
transform 1 0 142876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1547
timestamp 1670771148
transform 1 0 143428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1551
timestamp 1670771148
transform 1 0 143796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1571
timestamp 1670771148
transform 1 0 145636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1594
timestamp 1670771148
transform 1 0 147752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1597
timestamp 1670771148
transform 1 0 148028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1601
timestamp 1670771148
transform 1 0 148396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1618
timestamp 1670771148
transform 1 0 149960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1639
timestamp 1670771148
transform 1 0 151892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1650
timestamp 1670771148
transform 1 0 152904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1653
timestamp 1670771148
transform 1 0 153180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1675
timestamp 1670771148
transform 1 0 155204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1684
timestamp 1670771148
transform 1 0 156032 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1695
timestamp 1670771148
transform 1 0 157044 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1702
timestamp 1670771148
transform 1 0 157688 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1709
timestamp 1670771148
transform 1 0 158332 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1670771148
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1670771148
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1670771148
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1670771148
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1670771148
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1670771148
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1670771148
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp 1670771148
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp 1670771148
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_79
timestamp 1670771148
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_91
timestamp 1670771148
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1670771148
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1670771148
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1670771148
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1670771148
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1670771148
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1670771148
transform 1 0 13156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1670771148
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1670771148
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1670771148
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1670771148
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1670771148
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_173
timestamp 1670771148
transform 1 0 17020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_179
timestamp 1670771148
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_183
timestamp 1670771148
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1670771148
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_211
timestamp 1670771148
transform 1 0 20516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_217
timestamp 1670771148
transform 1 0 21068 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1670771148
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1670771148
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1670771148
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1670771148
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1670771148
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1670771148
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1670771148
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1670771148
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1670771148
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1670771148
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_317
timestamp 1670771148
transform 1 0 30268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_320
timestamp 1670771148
transform 1 0 30544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1670771148
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1670771148
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_343
timestamp 1670771148
transform 1 0 32660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_346
timestamp 1670771148
transform 1 0 32936 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_358
timestamp 1670771148
transform 1 0 34040 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_370
timestamp 1670771148
transform 1 0 35144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_382
timestamp 1670771148
transform 1 0 36248 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1670771148
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1670771148
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1670771148
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1670771148
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1670771148
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_441
timestamp 1670771148
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1670771148
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1670771148
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_467
timestamp 1670771148
transform 1 0 44068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_479
timestamp 1670771148
transform 1 0 45172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_491
timestamp 1670771148
transform 1 0 46276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1670771148
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1670771148
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_510
timestamp 1670771148
transform 1 0 48024 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_522
timestamp 1670771148
transform 1 0 49128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_534
timestamp 1670771148
transform 1 0 50232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_538
timestamp 1670771148
transform 1 0 50600 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_542
timestamp 1670771148
transform 1 0 50968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1670771148
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1670771148
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_573
timestamp 1670771148
transform 1 0 53820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_577
timestamp 1670771148
transform 1 0 54188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_594
timestamp 1670771148
transform 1 0 55752 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_600
timestamp 1670771148
transform 1 0 56304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_612
timestamp 1670771148
transform 1 0 57408 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1670771148
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1670771148
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_641
timestamp 1670771148
transform 1 0 60076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_660
timestamp 1670771148
transform 1 0 61824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_666
timestamp 1670771148
transform 1 0 62376 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1670771148
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1670771148
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1670771148
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1670771148
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1670771148
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1670771148
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1670771148
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1670771148
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1670771148
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1670771148
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1670771148
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1670771148
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1670771148
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_797
timestamp 1670771148
transform 1 0 74428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_817
timestamp 1670771148
transform 1 0 76268 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_823
timestamp 1670771148
transform 1 0 76820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_835
timestamp 1670771148
transform 1 0 77924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1670771148
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_841
timestamp 1670771148
transform 1 0 78476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_849
timestamp 1670771148
transform 1 0 79212 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_854
timestamp 1670771148
transform 1 0 79672 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_866
timestamp 1670771148
transform 1 0 80776 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_878
timestamp 1670771148
transform 1 0 81880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_890
timestamp 1670771148
transform 1 0 82984 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1670771148
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1670771148
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1670771148
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1670771148
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1670771148
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1670771148
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1670771148
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1670771148
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1670771148
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1670771148
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1670771148
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1670771148
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1670771148
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1670771148
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1670771148
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1670771148
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1670771148
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1670771148
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1670771148
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1670771148
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1670771148
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1670771148
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1670771148
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1670771148
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1121
timestamp 1670771148
transform 1 0 104236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1141
timestamp 1670771148
transform 1 0 106076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1147
timestamp 1670771148
transform 1 0 106628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1155
timestamp 1670771148
transform 1 0 107364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1174
timestamp 1670771148
transform 1 0 109112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1177
timestamp 1670771148
transform 1 0 109388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1195
timestamp 1670771148
transform 1 0 111044 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1670771148
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1670771148
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1670771148
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1670771148
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1670771148
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1670771148
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1670771148
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1269
timestamp 1670771148
transform 1 0 117852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1278
timestamp 1670771148
transform 1 0 118680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1286
timestamp 1670771148
transform 1 0 119416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1289
timestamp 1670771148
transform 1 0 119692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1293
timestamp 1670771148
transform 1 0 120060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1303
timestamp 1670771148
transform 1 0 120980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1309
timestamp 1670771148
transform 1 0 121532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1315
timestamp 1670771148
transform 1 0 122084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1335
timestamp 1670771148
transform 1 0 123924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1341
timestamp 1670771148
transform 1 0 124476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1345
timestamp 1670771148
transform 1 0 124844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1352
timestamp 1670771148
transform 1 0 125488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1374
timestamp 1670771148
transform 1 0 127512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1380
timestamp 1670771148
transform 1 0 128064 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1386
timestamp 1670771148
transform 1 0 128616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1389
timestamp 1670771148
transform 1 0 128892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1395
timestamp 1670771148
transform 1 0 129444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1670771148
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1401
timestamp 1670771148
transform 1 0 129996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1419
timestamp 1670771148
transform 1 0 131652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1439
timestamp 1670771148
transform 1 0 133492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1445
timestamp 1670771148
transform 1 0 134044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1448
timestamp 1670771148
transform 1 0 134320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1454
timestamp 1670771148
transform 1 0 134872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1457
timestamp 1670771148
transform 1 0 135148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1463
timestamp 1670771148
transform 1 0 135700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1466
timestamp 1670771148
transform 1 0 135976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1472
timestamp 1670771148
transform 1 0 136528 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1478
timestamp 1670771148
transform 1 0 137080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1484
timestamp 1670771148
transform 1 0 137632 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1504
timestamp 1670771148
transform 1 0 139472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1510
timestamp 1670771148
transform 1 0 140024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1513
timestamp 1670771148
transform 1 0 140300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1517
timestamp 1670771148
transform 1 0 140668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1523
timestamp 1670771148
transform 1 0 141220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1545
timestamp 1670771148
transform 1 0 143244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1565
timestamp 1670771148
transform 1 0 145084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1569
timestamp 1670771148
transform 1 0 145452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1576
timestamp 1670771148
transform 1 0 146096 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1598
timestamp 1670771148
transform 1 0 148120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1618
timestamp 1670771148
transform 1 0 149960 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1625
timestamp 1670771148
transform 1 0 150604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1644
timestamp 1670771148
transform 1 0 152352 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1650
timestamp 1670771148
transform 1 0 152904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1670
timestamp 1670771148
transform 1 0 154744 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1677
timestamp 1670771148
transform 1 0 155388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1681
timestamp 1670771148
transform 1 0 155756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1688
timestamp 1670771148
transform 1 0 156400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1695
timestamp 1670771148
transform 1 0 157044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1702
timestamp 1670771148
transform 1 0 157688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1709
timestamp 1670771148
transform 1 0 158332 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1670771148
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1670771148
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1670771148
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1670771148
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1670771148
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1670771148
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_51
timestamp 1670771148
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_63
timestamp 1670771148
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1670771148
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1670771148
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1670771148
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1670771148
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_109
timestamp 1670771148
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_117
timestamp 1670771148
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1670771148
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1670771148
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1670771148
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1670771148
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 1670771148
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1670771148
transform 1 0 15272 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_160
timestamp 1670771148
transform 1 0 15824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1670771148
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_183
timestamp 1670771148
transform 1 0 17940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp 1670771148
transform 1 0 18676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1670771148
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1670771148
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1670771148
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_236
timestamp 1670771148
transform 1 0 22816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1670771148
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1670771148
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1670771148
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_261
timestamp 1670771148
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_264
timestamp 1670771148
transform 1 0 25392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_273
timestamp 1670771148
transform 1 0 26220 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_279
timestamp 1670771148
transform 1 0 26772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_291
timestamp 1670771148
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1670771148
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1670771148
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1670771148
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_318
timestamp 1670771148
transform 1 0 30360 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_325
timestamp 1670771148
transform 1 0 31004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1670771148
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1670771148
transform 1 0 33212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1670771148
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1670771148
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1670771148
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1670771148
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1670771148
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1670771148
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1670771148
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1670771148
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1670771148
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_445
timestamp 1670771148
transform 1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_449
timestamp 1670771148
transform 1 0 42412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1670771148
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1670771148
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1670771148
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_492
timestamp 1670771148
transform 1 0 46368 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_504
timestamp 1670771148
transform 1 0 47472 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_516
timestamp 1670771148
transform 1 0 48576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1670771148
transform 1 0 49680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_533
timestamp 1670771148
transform 1 0 50140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_538
timestamp 1670771148
transform 1 0 50600 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_558
timestamp 1670771148
transform 1 0 52440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_570
timestamp 1670771148
transform 1 0 53544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_582
timestamp 1670771148
transform 1 0 54648 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1670771148
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1670771148
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1670771148
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1670771148
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1670771148
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1670771148
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1670771148
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1670771148
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1670771148
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1670771148
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1670771148
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1670771148
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1670771148
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1670771148
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1670771148
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1670771148
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1670771148
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1670771148
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1670771148
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1670771148
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_781
timestamp 1670771148
transform 1 0 72956 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_786
timestamp 1670771148
transform 1 0 73416 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_798
timestamp 1670771148
transform 1 0 74520 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_810
timestamp 1670771148
transform 1 0 75624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_813
timestamp 1670771148
transform 1 0 75900 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_819
timestamp 1670771148
transform 1 0 76452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_831
timestamp 1670771148
transform 1 0 77556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_843
timestamp 1670771148
transform 1 0 78660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_855
timestamp 1670771148
transform 1 0 79764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1670771148
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_869
timestamp 1670771148
transform 1 0 81052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_875
timestamp 1670771148
transform 1 0 81604 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_884
timestamp 1670771148
transform 1 0 82432 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_896
timestamp 1670771148
transform 1 0 83536 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_907
timestamp 1670771148
transform 1 0 84548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_919
timestamp 1670771148
transform 1 0 85652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1670771148
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1670771148
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_937
timestamp 1670771148
transform 1 0 87308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_945
timestamp 1670771148
transform 1 0 88044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_949
timestamp 1670771148
transform 1 0 88412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_969
timestamp 1670771148
transform 1 0 90252 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_977
timestamp 1670771148
transform 1 0 90988 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1670771148
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_993
timestamp 1670771148
transform 1 0 92460 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_998
timestamp 1670771148
transform 1 0 92920 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1010
timestamp 1670771148
transform 1 0 94024 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1022
timestamp 1670771148
transform 1 0 95128 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1030
timestamp 1670771148
transform 1 0 95864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1034
timestamp 1670771148
transform 1 0 96232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1037
timestamp 1670771148
transform 1 0 96508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1055
timestamp 1670771148
transform 1 0 98164 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1670771148
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1670771148
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1670771148
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1670771148
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1670771148
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1670771148
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1117
timestamp 1670771148
transform 1 0 103868 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1125
timestamp 1670771148
transform 1 0 104604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1137
timestamp 1670771148
transform 1 0 105708 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1145
timestamp 1670771148
transform 1 0 106444 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1670771148
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1161
timestamp 1670771148
transform 1 0 107916 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1181
timestamp 1670771148
transform 1 0 109756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1193
timestamp 1670771148
transform 1 0 110860 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1201
timestamp 1670771148
transform 1 0 111596 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1670771148
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1217
timestamp 1670771148
transform 1 0 113068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1221
timestamp 1670771148
transform 1 0 113436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1238
timestamp 1670771148
transform 1 0 115000 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1244
timestamp 1670771148
transform 1 0 115552 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1256
timestamp 1670771148
transform 1 0 116656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1261
timestamp 1670771148
transform 1 0 117116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1267
timestamp 1670771148
transform 1 0 117668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1270
timestamp 1670771148
transform 1 0 117944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1278
timestamp 1670771148
transform 1 0 118680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1284
timestamp 1670771148
transform 1 0 119232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1290
timestamp 1670771148
transform 1 0 119784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1296
timestamp 1670771148
transform 1 0 120336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1302
timestamp 1670771148
transform 1 0 120888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1308
timestamp 1670771148
transform 1 0 121440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1314
timestamp 1670771148
transform 1 0 121992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1317
timestamp 1670771148
transform 1 0 122268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1323
timestamp 1670771148
transform 1 0 122820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1340
timestamp 1670771148
transform 1 0 124384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1346
timestamp 1670771148
transform 1 0 124936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1352
timestamp 1670771148
transform 1 0 125488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1358
timestamp 1670771148
transform 1 0 126040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1364
timestamp 1670771148
transform 1 0 126592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1370
timestamp 1670771148
transform 1 0 127144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1373
timestamp 1670771148
transform 1 0 127420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1377
timestamp 1670771148
transform 1 0 127788 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1394
timestamp 1670771148
transform 1 0 129352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1400
timestamp 1670771148
transform 1 0 129904 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1408
timestamp 1670771148
transform 1 0 130640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1414
timestamp 1670771148
transform 1 0 131192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1420
timestamp 1670771148
transform 1 0 131744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1426
timestamp 1670771148
transform 1 0 132296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1429
timestamp 1670771148
transform 1 0 132572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1437
timestamp 1670771148
transform 1 0 133308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1457
timestamp 1670771148
transform 1 0 135148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1465
timestamp 1670771148
transform 1 0 135884 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1482
timestamp 1670771148
transform 1 0 137448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1485
timestamp 1670771148
transform 1 0 137724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1489
timestamp 1670771148
transform 1 0 138092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1495
timestamp 1670771148
transform 1 0 138644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1501
timestamp 1670771148
transform 1 0 139196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1508
timestamp 1670771148
transform 1 0 139840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1517
timestamp 1670771148
transform 1 0 140668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1537
timestamp 1670771148
transform 1 0 142508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1541
timestamp 1670771148
transform 1 0 142876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1548
timestamp 1670771148
transform 1 0 143520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1572
timestamp 1670771148
transform 1 0 145728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1592
timestamp 1670771148
transform 1 0 147568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1597
timestamp 1670771148
transform 1 0 148028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1615
timestamp 1670771148
transform 1 0 149684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1635
timestamp 1670771148
transform 1 0 151524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1644
timestamp 1670771148
transform 1 0 152352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1650
timestamp 1670771148
transform 1 0 152904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1653
timestamp 1670771148
transform 1 0 153180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1662
timestamp 1670771148
transform 1 0 154008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1669
timestamp 1670771148
transform 1 0 154652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1673
timestamp 1670771148
transform 1 0 155020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1679
timestamp 1670771148
transform 1 0 155572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1686
timestamp 1670771148
transform 1 0 156216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1693
timestamp 1670771148
transform 1 0 156860 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1700
timestamp 1670771148
transform 1 0 157504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1706
timestamp 1670771148
transform 1 0 158056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1709
timestamp 1670771148
transform 1 0 158332 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1670771148
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1670771148
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1670771148
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1670771148
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1670771148
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1670771148
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_61
timestamp 1670771148
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_73
timestamp 1670771148
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_85
timestamp 1670771148
transform 1 0 8924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1670771148
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1670771148
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1670771148
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1670771148
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_147
timestamp 1670771148
transform 1 0 14628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_156
timestamp 1670771148
transform 1 0 15456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1670771148
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1670771148
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_173
timestamp 1670771148
transform 1 0 17020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1670771148
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_187
timestamp 1670771148
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp 1670771148
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1670771148
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1670771148
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1670771148
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1670771148
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_233
timestamp 1670771148
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1670771148
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1670771148
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1670771148
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1670771148
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_285
timestamp 1670771148
transform 1 0 27324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_297
timestamp 1670771148
transform 1 0 28428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_314
timestamp 1670771148
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1670771148
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1670771148
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_349
timestamp 1670771148
transform 1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_357
timestamp 1670771148
transform 1 0 33948 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1670771148
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_365
timestamp 1670771148
transform 1 0 34684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_368
timestamp 1670771148
transform 1 0 34960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1670771148
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1670771148
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1670771148
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1670771148
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1670771148
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1670771148
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1670771148
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1670771148
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1670771148
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_473
timestamp 1670771148
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_479
timestamp 1670771148
transform 1 0 45172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_482
timestamp 1670771148
transform 1 0 45448 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_494
timestamp 1670771148
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1670771148
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1670771148
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_513
timestamp 1670771148
transform 1 0 48300 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_518
timestamp 1670771148
transform 1 0 48760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_530
timestamp 1670771148
transform 1 0 49864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_542
timestamp 1670771148
transform 1 0 50968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_554
timestamp 1670771148
transform 1 0 52072 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_561
timestamp 1670771148
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_579
timestamp 1670771148
transform 1 0 54372 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_587
timestamp 1670771148
transform 1 0 55108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_606
timestamp 1670771148
transform 1 0 56856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1670771148
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1670771148
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1670771148
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_641
timestamp 1670771148
transform 1 0 60076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_649
timestamp 1670771148
transform 1 0 60812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_667
timestamp 1670771148
transform 1 0 62468 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1670771148
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_673
timestamp 1670771148
transform 1 0 63020 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_677
timestamp 1670771148
transform 1 0 63388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_689
timestamp 1670771148
transform 1 0 64492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_703
timestamp 1670771148
transform 1 0 65780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_715
timestamp 1670771148
transform 1 0 66884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1670771148
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1670771148
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1670771148
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1670771148
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1670771148
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1670771148
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1670771148
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_785
timestamp 1670771148
transform 1 0 73324 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_789
timestamp 1670771148
transform 1 0 73692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_801
timestamp 1670771148
transform 1 0 74796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_804
timestamp 1670771148
transform 1 0 75072 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_828
timestamp 1670771148
transform 1 0 77280 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_841
timestamp 1670771148
transform 1 0 78476 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_848
timestamp 1670771148
transform 1 0 79120 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_860
timestamp 1670771148
transform 1 0 80224 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_872
timestamp 1670771148
transform 1 0 81328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_876
timestamp 1670771148
transform 1 0 81696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_879
timestamp 1670771148
transform 1 0 81972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_888
timestamp 1670771148
transform 1 0 82800 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1670771148
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1670771148
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1670771148
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1670771148
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1670771148
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1670771148
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1670771148
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_965
timestamp 1670771148
transform 1 0 89884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_973
timestamp 1670771148
transform 1 0 90620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_976
timestamp 1670771148
transform 1 0 90896 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_996
timestamp 1670771148
transform 1 0 92736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1003
timestamp 1670771148
transform 1 0 93380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1670771148
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1670771148
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1670771148
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1670771148
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1670771148
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1670771148
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1670771148
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1670771148
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1670771148
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1670771148
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1670771148
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1670771148
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1670771148
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1121
timestamp 1670771148
transform 1 0 104236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1141
timestamp 1670771148
transform 1 0 106076 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1147
timestamp 1670771148
transform 1 0 106628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1159
timestamp 1670771148
transform 1 0 107732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1171
timestamp 1670771148
transform 1 0 108836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1670771148
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1670771148
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1670771148
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1201
timestamp 1670771148
transform 1 0 111596 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1210
timestamp 1670771148
transform 1 0 112424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1222
timestamp 1670771148
transform 1 0 113528 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1230
timestamp 1670771148
transform 1 0 114264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1233
timestamp 1670771148
transform 1 0 114540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1240
timestamp 1670771148
transform 1 0 115184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1246
timestamp 1670771148
transform 1 0 115736 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1268
timestamp 1670771148
transform 1 0 117760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1279
timestamp 1670771148
transform 1 0 118772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1283
timestamp 1670771148
transform 1 0 119140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1286
timestamp 1670771148
transform 1 0 119416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1289
timestamp 1670771148
transform 1 0 119692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1307
timestamp 1670771148
transform 1 0 121348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1327
timestamp 1670771148
transform 1 0 123188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1333
timestamp 1670771148
transform 1 0 123740 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1336
timestamp 1670771148
transform 1 0 124016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1342
timestamp 1670771148
transform 1 0 124568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1345
timestamp 1670771148
transform 1 0 124844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1357
timestamp 1670771148
transform 1 0 125948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1363
timestamp 1670771148
transform 1 0 126500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1366
timestamp 1670771148
transform 1 0 126776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1372
timestamp 1670771148
transform 1 0 127328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1381
timestamp 1670771148
transform 1 0 128156 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1389
timestamp 1670771148
transform 1 0 128892 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1392
timestamp 1670771148
transform 1 0 129168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1398
timestamp 1670771148
transform 1 0 129720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1401
timestamp 1670771148
transform 1 0 129996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1406
timestamp 1670771148
transform 1 0 130456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1412
timestamp 1670771148
transform 1 0 131008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1418
timestamp 1670771148
transform 1 0 131560 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1424
timestamp 1670771148
transform 1 0 132112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1430
timestamp 1670771148
transform 1 0 132664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1436
timestamp 1670771148
transform 1 0 133216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1442
timestamp 1670771148
transform 1 0 133768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1448
timestamp 1670771148
transform 1 0 134320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1454
timestamp 1670771148
transform 1 0 134872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1457
timestamp 1670771148
transform 1 0 135148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1465
timestamp 1670771148
transform 1 0 135884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1471
timestamp 1670771148
transform 1 0 136436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1478
timestamp 1670771148
transform 1 0 137080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1488
timestamp 1670771148
transform 1 0 138000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1495
timestamp 1670771148
transform 1 0 138644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1503
timestamp 1670771148
transform 1 0 139380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1510
timestamp 1670771148
transform 1 0 140024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1513
timestamp 1670771148
transform 1 0 140300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1532
timestamp 1670771148
transform 1 0 142048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1552
timestamp 1670771148
transform 1 0 143888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1565
timestamp 1670771148
transform 1 0 145084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1569
timestamp 1670771148
transform 1 0 145452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1587
timestamp 1670771148
transform 1 0 147108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1607
timestamp 1670771148
transform 1 0 148948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1619
timestamp 1670771148
transform 1 0 150052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1670771148
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1625
timestamp 1670771148
transform 1 0 150604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1643
timestamp 1670771148
transform 1 0 152260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1652
timestamp 1670771148
transform 1 0 153088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1659
timestamp 1670771148
transform 1 0 153732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1667
timestamp 1670771148
transform 1 0 154468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1670771148
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1670771148
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1681
timestamp 1670771148
transform 1 0 155756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1688
timestamp 1670771148
transform 1 0 156400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1695
timestamp 1670771148
transform 1 0 157044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1702
timestamp 1670771148
transform 1 0 157688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1709
timestamp 1670771148
transform 1 0 158332 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1670771148
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1670771148
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1670771148
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1670771148
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1670771148
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_54
timestamp 1670771148
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1670771148
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1670771148
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1670771148
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1670771148
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1670771148
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1670771148
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_117
timestamp 1670771148
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_132
timestamp 1670771148
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1670771148
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1670771148
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1670771148
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1670771148
transform 1 0 16560 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1670771148
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_185
timestamp 1670771148
transform 1 0 18124 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1670771148
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1670771148
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_204
timestamp 1670771148
transform 1 0 19872 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_216
timestamp 1670771148
transform 1 0 20976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_224
timestamp 1670771148
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_227
timestamp 1670771148
transform 1 0 21988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_239
timestamp 1670771148
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1670771148
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1670771148
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_258
timestamp 1670771148
transform 1 0 24840 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_270
timestamp 1670771148
transform 1 0 25944 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_282
timestamp 1670771148
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1670771148
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1670771148
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1670771148
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1670771148
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_319
timestamp 1670771148
transform 1 0 30452 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_325
timestamp 1670771148
transform 1 0 31004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_337
timestamp 1670771148
transform 1 0 32108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_340
timestamp 1670771148
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_352
timestamp 1670771148
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1670771148
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1670771148
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1670771148
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_402
timestamp 1670771148
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_408
timestamp 1670771148
transform 1 0 38640 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1670771148
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1670771148
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1670771148
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_457
timestamp 1670771148
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1670771148
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_477
timestamp 1670771148
transform 1 0 44988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_481
timestamp 1670771148
transform 1 0 45356 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_487
timestamp 1670771148
transform 1 0 45908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_499
timestamp 1670771148
transform 1 0 47012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_504
timestamp 1670771148
transform 1 0 47472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_524
timestamp 1670771148
transform 1 0 49312 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1670771148
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_545
timestamp 1670771148
transform 1 0 51244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_553
timestamp 1670771148
transform 1 0 51980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_571
timestamp 1670771148
transform 1 0 53636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_578
timestamp 1670771148
transform 1 0 54280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_584
timestamp 1670771148
transform 1 0 54832 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1670771148
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1670771148
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_613
timestamp 1670771148
transform 1 0 57500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_621
timestamp 1670771148
transform 1 0 58236 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_626
timestamp 1670771148
transform 1 0 58696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_638
timestamp 1670771148
transform 1 0 59800 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1670771148
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1670771148
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1670771148
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_681
timestamp 1670771148
transform 1 0 63756 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_698
timestamp 1670771148
transform 1 0 65320 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_701
timestamp 1670771148
transform 1 0 65596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_708
timestamp 1670771148
transform 1 0 66240 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_714
timestamp 1670771148
transform 1 0 66792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_726
timestamp 1670771148
transform 1 0 67896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_730
timestamp 1670771148
transform 1 0 68264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_733
timestamp 1670771148
transform 1 0 68540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_753
timestamp 1670771148
transform 1 0 70380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1670771148
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_769
timestamp 1670771148
transform 1 0 71852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_777
timestamp 1670771148
transform 1 0 72588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_783
timestamp 1670771148
transform 1 0 73140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_789
timestamp 1670771148
transform 1 0 73692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_809
timestamp 1670771148
transform 1 0 75532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_813
timestamp 1670771148
transform 1 0 75900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_818
timestamp 1670771148
transform 1 0 76360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_842
timestamp 1670771148
transform 1 0 78568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_846
timestamp 1670771148
transform 1 0 78936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_863
timestamp 1670771148
transform 1 0 80500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1670771148
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_869
timestamp 1670771148
transform 1 0 81052 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_891
timestamp 1670771148
transform 1 0 83076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_903
timestamp 1670771148
transform 1 0 84180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_915
timestamp 1670771148
transform 1 0 85284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1670771148
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1670771148
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1670771148
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1670771148
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1670771148
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1670771148
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1670771148
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_981
timestamp 1670771148
transform 1 0 91356 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_987
timestamp 1670771148
transform 1 0 91908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_999
timestamp 1670771148
transform 1 0 93012 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1005
timestamp 1670771148
transform 1 0 93564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1025
timestamp 1670771148
transform 1 0 95404 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1033
timestamp 1670771148
transform 1 0 96140 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1670771148
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1670771148
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1061
timestamp 1670771148
transform 1 0 98716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1069
timestamp 1670771148
transform 1 0 99452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1090
timestamp 1670771148
transform 1 0 101384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1093
timestamp 1670771148
transform 1 0 101660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1097
timestamp 1670771148
transform 1 0 102028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1109
timestamp 1670771148
transform 1 0 103132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1121
timestamp 1670771148
transform 1 0 104236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1133
timestamp 1670771148
transform 1 0 105340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1145
timestamp 1670771148
transform 1 0 106444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1149
timestamp 1670771148
transform 1 0 106812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1167
timestamp 1670771148
transform 1 0 108468 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1670771148
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1670771148
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1670771148
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1670771148
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1670771148
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1670771148
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1229
timestamp 1670771148
transform 1 0 114172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1232
timestamp 1670771148
transform 1 0 114448 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1240
timestamp 1670771148
transform 1 0 115184 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1258
timestamp 1670771148
transform 1 0 116840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1261
timestamp 1670771148
transform 1 0 117116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1265
timestamp 1670771148
transform 1 0 117484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1273
timestamp 1670771148
transform 1 0 118220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1277
timestamp 1670771148
transform 1 0 118588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1297
timestamp 1670771148
transform 1 0 120428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1306
timestamp 1670771148
transform 1 0 121256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1312
timestamp 1670771148
transform 1 0 121808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1317
timestamp 1670771148
transform 1 0 122268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1321
timestamp 1670771148
transform 1 0 122636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1327
timestamp 1670771148
transform 1 0 123188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1333
timestamp 1670771148
transform 1 0 123740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1343
timestamp 1670771148
transform 1 0 124660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1349
timestamp 1670771148
transform 1 0 125212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1356
timestamp 1670771148
transform 1 0 125856 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1364
timestamp 1670771148
transform 1 0 126592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1370
timestamp 1670771148
transform 1 0 127144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1373
timestamp 1670771148
transform 1 0 127420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1391
timestamp 1670771148
transform 1 0 129076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1399
timestamp 1670771148
transform 1 0 129812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1407
timestamp 1670771148
transform 1 0 130548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1413
timestamp 1670771148
transform 1 0 131100 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1416
timestamp 1670771148
transform 1 0 131376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1424
timestamp 1670771148
transform 1 0 132112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1429
timestamp 1670771148
transform 1 0 132572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1434
timestamp 1670771148
transform 1 0 133032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1440
timestamp 1670771148
transform 1 0 133584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1446
timestamp 1670771148
transform 1 0 134136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1452
timestamp 1670771148
transform 1 0 134688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1458
timestamp 1670771148
transform 1 0 135240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1464
timestamp 1670771148
transform 1 0 135792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1470
timestamp 1670771148
transform 1 0 136344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1476
timestamp 1670771148
transform 1 0 136896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1482
timestamp 1670771148
transform 1 0 137448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1485
timestamp 1670771148
transform 1 0 137724 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1489
timestamp 1670771148
transform 1 0 138092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1509
timestamp 1670771148
transform 1 0 139932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1516
timestamp 1670771148
transform 1 0 140576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1536
timestamp 1670771148
transform 1 0 142416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1541
timestamp 1670771148
transform 1 0 142876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1559
timestamp 1670771148
transform 1 0 144532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1579
timestamp 1670771148
transform 1 0 146372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1588
timestamp 1670771148
transform 1 0 147200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1594
timestamp 1670771148
transform 1 0 147752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1597
timestamp 1670771148
transform 1 0 148028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1615
timestamp 1670771148
transform 1 0 149684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1624
timestamp 1670771148
transform 1 0 150512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1631
timestamp 1670771148
transform 1 0 151156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1635
timestamp 1670771148
transform 1 0 151524 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1639
timestamp 1670771148
transform 1 0 151892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1646
timestamp 1670771148
transform 1 0 152536 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1653
timestamp 1670771148
transform 1 0 153180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1657
timestamp 1670771148
transform 1 0 153548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1663
timestamp 1670771148
transform 1 0 154100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1672
timestamp 1670771148
transform 1 0 154928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1681
timestamp 1670771148
transform 1 0 155756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1690
timestamp 1670771148
transform 1 0 156584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1697
timestamp 1670771148
transform 1 0 157228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1704
timestamp 1670771148
transform 1 0 157872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1709
timestamp 1670771148
transform 1 0 158332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1670771148
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 1670771148
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_14
timestamp 1670771148
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1670771148
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_38
timestamp 1670771148
transform 1 0 4600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1670771148
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1670771148
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1670771148
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1670771148
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1670771148
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1670771148
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1670771148
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1670771148
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1670771148
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1670771148
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1670771148
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_137
timestamp 1670771148
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1670771148
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1670771148
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1670771148
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1670771148
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1670771148
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1670771148
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1670771148
transform 1 0 17296 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_180
timestamp 1670771148
transform 1 0 17664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1670771148
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1670771148
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_199
timestamp 1670771148
transform 1 0 19412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_207
timestamp 1670771148
transform 1 0 20148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1670771148
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1670771148
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1670771148
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_232
timestamp 1670771148
transform 1 0 22448 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_244
timestamp 1670771148
transform 1 0 23552 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_263
timestamp 1670771148
transform 1 0 25300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1670771148
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1670771148
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 1670771148
transform 1 0 28060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_303
timestamp 1670771148
transform 1 0 28980 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_323
timestamp 1670771148
transform 1 0 30820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1670771148
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp 1670771148
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_356
timestamp 1670771148
transform 1 0 33856 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_362
timestamp 1670771148
transform 1 0 34408 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_374
timestamp 1670771148
transform 1 0 35512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1670771148
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1670771148
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_401
timestamp 1670771148
transform 1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_421
timestamp 1670771148
transform 1 0 39836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_430
timestamp 1670771148
transform 1 0 40664 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_436
timestamp 1670771148
transform 1 0 41216 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1670771148
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_461
timestamp 1670771148
transform 1 0 43516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_469
timestamp 1670771148
transform 1 0 44252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_489
timestamp 1670771148
transform 1 0 46092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_496
timestamp 1670771148
transform 1 0 46736 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1670771148
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1670771148
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1670771148
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_543
timestamp 1670771148
transform 1 0 51060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_552
timestamp 1670771148
transform 1 0 51888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_558
timestamp 1670771148
transform 1 0 52440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_561
timestamp 1670771148
transform 1 0 52716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_565
timestamp 1670771148
transform 1 0 53084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_569
timestamp 1670771148
transform 1 0 53452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_575
timestamp 1670771148
transform 1 0 54004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_592
timestamp 1670771148
transform 1 0 55568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_600
timestamp 1670771148
transform 1 0 56304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_605
timestamp 1670771148
transform 1 0 56764 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_613
timestamp 1670771148
transform 1 0 57500 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1670771148
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_629
timestamp 1670771148
transform 1 0 58972 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_639
timestamp 1670771148
transform 1 0 59892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_651
timestamp 1670771148
transform 1 0 60996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_663
timestamp 1670771148
transform 1 0 62100 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1670771148
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_673
timestamp 1670771148
transform 1 0 63020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_681
timestamp 1670771148
transform 1 0 63756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_701
timestamp 1670771148
transform 1 0 65596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_707
timestamp 1670771148
transform 1 0 66148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_715
timestamp 1670771148
transform 1 0 66884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1670771148
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1670771148
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1670771148
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_743
timestamp 1670771148
transform 1 0 69460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_763
timestamp 1670771148
transform 1 0 71300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_769
timestamp 1670771148
transform 1 0 71852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_777
timestamp 1670771148
transform 1 0 72588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_782
timestamp 1670771148
transform 1 0 73048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_785
timestamp 1670771148
transform 1 0 73324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_789
timestamp 1670771148
transform 1 0 73692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_792
timestamp 1670771148
transform 1 0 73968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_800
timestamp 1670771148
transform 1 0 74704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_819
timestamp 1670771148
transform 1 0 76452 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_825
timestamp 1670771148
transform 1 0 77004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_837
timestamp 1670771148
transform 1 0 78108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_841
timestamp 1670771148
transform 1 0 78476 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_847
timestamp 1670771148
transform 1 0 79028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_859
timestamp 1670771148
transform 1 0 80132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_871
timestamp 1670771148
transform 1 0 81236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_883
timestamp 1670771148
transform 1 0 82340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1670771148
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1670771148
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_909
timestamp 1670771148
transform 1 0 84732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_917
timestamp 1670771148
transform 1 0 85468 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_921
timestamp 1670771148
transform 1 0 85836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_941
timestamp 1670771148
transform 1 0 87676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_947
timestamp 1670771148
transform 1 0 88228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1670771148
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_953
timestamp 1670771148
transform 1 0 88780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_957
timestamp 1670771148
transform 1 0 89148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_977
timestamp 1670771148
transform 1 0 90988 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_983
timestamp 1670771148
transform 1 0 91540 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_992
timestamp 1670771148
transform 1 0 92368 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1004
timestamp 1670771148
transform 1 0 93472 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1670771148
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1670771148
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1033
timestamp 1670771148
transform 1 0 96140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1039
timestamp 1670771148
transform 1 0 96692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1060
timestamp 1670771148
transform 1 0 98624 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1670771148
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1077
timestamp 1670771148
transform 1 0 100188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1083
timestamp 1670771148
transform 1 0 100740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1086
timestamp 1670771148
transform 1 0 101016 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1096
timestamp 1670771148
transform 1 0 101936 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1108
timestamp 1670771148
transform 1 0 103040 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1121
timestamp 1670771148
transform 1 0 104236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1129
timestamp 1670771148
transform 1 0 104972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1147
timestamp 1670771148
transform 1 0 106628 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1171
timestamp 1670771148
transform 1 0 108836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1670771148
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1177
timestamp 1670771148
transform 1 0 109388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1181
timestamp 1670771148
transform 1 0 109756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1189
timestamp 1670771148
transform 1 0 110492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1193
timestamp 1670771148
transform 1 0 110860 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1199
timestamp 1670771148
transform 1 0 111412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1211
timestamp 1670771148
transform 1 0 112516 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1221
timestamp 1670771148
transform 1 0 113436 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1230
timestamp 1670771148
transform 1 0 114264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1233
timestamp 1670771148
transform 1 0 114540 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1251
timestamp 1670771148
transform 1 0 116196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1257
timestamp 1670771148
transform 1 0 116748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1263
timestamp 1670771148
transform 1 0 117300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1271
timestamp 1670771148
transform 1 0 118036 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1274
timestamp 1670771148
transform 1 0 118312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1280
timestamp 1670771148
transform 1 0 118864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1286
timestamp 1670771148
transform 1 0 119416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1289
timestamp 1670771148
transform 1 0 119692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1307
timestamp 1670771148
transform 1 0 121348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1327
timestamp 1670771148
transform 1 0 123188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1333
timestamp 1670771148
transform 1 0 123740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1339
timestamp 1670771148
transform 1 0 124292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1342
timestamp 1670771148
transform 1 0 124568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1345
timestamp 1670771148
transform 1 0 124844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1351
timestamp 1670771148
transform 1 0 125396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1368
timestamp 1670771148
transform 1 0 126960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1374
timestamp 1670771148
transform 1 0 127512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1380
timestamp 1670771148
transform 1 0 128064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1386
timestamp 1670771148
transform 1 0 128616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1392
timestamp 1670771148
transform 1 0 129168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1398
timestamp 1670771148
transform 1 0 129720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1401
timestamp 1670771148
transform 1 0 129996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1405
timestamp 1670771148
transform 1 0 130364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1409
timestamp 1670771148
transform 1 0 130732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1412
timestamp 1670771148
transform 1 0 131008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1418
timestamp 1670771148
transform 1 0 131560 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1424
timestamp 1670771148
transform 1 0 132112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1430
timestamp 1670771148
transform 1 0 132664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1436
timestamp 1670771148
transform 1 0 133216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1442
timestamp 1670771148
transform 1 0 133768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1448
timestamp 1670771148
transform 1 0 134320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1454
timestamp 1670771148
transform 1 0 134872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1457
timestamp 1670771148
transform 1 0 135148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1465
timestamp 1670771148
transform 1 0 135884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1471
timestamp 1670771148
transform 1 0 136436 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1477
timestamp 1670771148
transform 1 0 136988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1483
timestamp 1670771148
transform 1 0 137540 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1486
timestamp 1670771148
transform 1 0 137816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1492
timestamp 1670771148
transform 1 0 138368 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1498
timestamp 1670771148
transform 1 0 138920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1504
timestamp 1670771148
transform 1 0 139472 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1510
timestamp 1670771148
transform 1 0 140024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1513
timestamp 1670771148
transform 1 0 140300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1517
timestamp 1670771148
transform 1 0 140668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1543
timestamp 1670771148
transform 1 0 143060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1563
timestamp 1670771148
transform 1 0 144900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1670771148
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1569
timestamp 1670771148
transform 1 0 145452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1587
timestamp 1670771148
transform 1 0 147108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1607
timestamp 1670771148
transform 1 0 148948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1615
timestamp 1670771148
transform 1 0 149684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1622
timestamp 1670771148
transform 1 0 150328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1625
timestamp 1670771148
transform 1 0 150604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1630
timestamp 1670771148
transform 1 0 151064 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1639
timestamp 1670771148
transform 1 0 151892 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1650
timestamp 1670771148
transform 1 0 152904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1656
timestamp 1670771148
transform 1 0 153456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1661
timestamp 1670771148
transform 1 0 153916 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1669
timestamp 1670771148
transform 1 0 154652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1675
timestamp 1670771148
transform 1 0 155204 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1670771148
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1681
timestamp 1670771148
transform 1 0 155756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1688
timestamp 1670771148
transform 1 0 156400 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1695
timestamp 1670771148
transform 1 0 157044 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1702
timestamp 1670771148
transform 1 0 157688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1709
timestamp 1670771148
transform 1 0 158332 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1670771148
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1670771148
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1670771148
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1670771148
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_40
timestamp 1670771148
transform 1 0 4784 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1670771148
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1670771148
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1670771148
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1670771148
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1670771148
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1670771148
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_118
timestamp 1670771148
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1670771148
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_130
timestamp 1670771148
transform 1 0 13064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1670771148
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1670771148
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1670771148
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_156
timestamp 1670771148
transform 1 0 15456 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_180
timestamp 1670771148
transform 1 0 17664 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_186
timestamp 1670771148
transform 1 0 18216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1670771148
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1670771148
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1670771148
transform 1 0 19596 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1670771148
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_222
timestamp 1670771148
transform 1 0 21528 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_231
timestamp 1670771148
transform 1 0 22356 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_237
timestamp 1670771148
transform 1 0 22908 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp 1670771148
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1670771148
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1670771148
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1670771148
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_274
timestamp 1670771148
transform 1 0 26312 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_283
timestamp 1670771148
transform 1 0 27140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_295
timestamp 1670771148
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1670771148
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1670771148
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1670771148
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_333
timestamp 1670771148
transform 1 0 31740 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_341
timestamp 1670771148
transform 1 0 32476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_345
timestamp 1670771148
transform 1 0 32844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_351
timestamp 1670771148
transform 1 0 33396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1670771148
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1670771148
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1670771148
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_369
timestamp 1670771148
transform 1 0 35052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_381
timestamp 1670771148
transform 1 0 36156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_386
timestamp 1670771148
transform 1 0 36616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_392
timestamp 1670771148
transform 1 0 37168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_398
timestamp 1670771148
transform 1 0 37720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_418
timestamp 1670771148
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1670771148
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1670771148
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1670771148
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_457
timestamp 1670771148
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_466
timestamp 1670771148
transform 1 0 43976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_472
timestamp 1670771148
transform 1 0 44528 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1670771148
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1670771148
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1670771148
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1670771148
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1670771148
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1670771148
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_533
timestamp 1670771148
transform 1 0 50140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_537
timestamp 1670771148
transform 1 0 50508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_540
timestamp 1670771148
transform 1 0 50784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_550
timestamp 1670771148
transform 1 0 51704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_556
timestamp 1670771148
transform 1 0 52256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_562
timestamp 1670771148
transform 1 0 52808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_570
timestamp 1670771148
transform 1 0 53544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_576
timestamp 1670771148
transform 1 0 54096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_582
timestamp 1670771148
transform 1 0 54648 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_589
timestamp 1670771148
transform 1 0 55292 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_593
timestamp 1670771148
transform 1 0 55660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_605
timestamp 1670771148
transform 1 0 56764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_613
timestamp 1670771148
transform 1 0 57500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_616
timestamp 1670771148
transform 1 0 57776 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_628
timestamp 1670771148
transform 1 0 58880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1670771148
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1670771148
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1670771148
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1670771148
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_669
timestamp 1670771148
transform 1 0 62652 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_677
timestamp 1670771148
transform 1 0 63388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_696
timestamp 1670771148
transform 1 0 65136 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_701
timestamp 1670771148
transform 1 0 65596 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_705
timestamp 1670771148
transform 1 0 65964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_727
timestamp 1670771148
transform 1 0 67988 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_733
timestamp 1670771148
transform 1 0 68540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_745
timestamp 1670771148
transform 1 0 69644 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_753
timestamp 1670771148
transform 1 0 70380 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1670771148
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_769
timestamp 1670771148
transform 1 0 71852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_773
timestamp 1670771148
transform 1 0 72220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_790
timestamp 1670771148
transform 1 0 73784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_810
timestamp 1670771148
transform 1 0 75624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_813
timestamp 1670771148
transform 1 0 75900 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_817
timestamp 1670771148
transform 1 0 76268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_829
timestamp 1670771148
transform 1 0 77372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_841
timestamp 1670771148
transform 1 0 78476 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_847
timestamp 1670771148
transform 1 0 79028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_859
timestamp 1670771148
transform 1 0 80132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1670771148
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_869
timestamp 1670771148
transform 1 0 81052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_887
timestamp 1670771148
transform 1 0 82708 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1670771148
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1670771148
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_917
timestamp 1670771148
transform 1 0 85468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_922
timestamp 1670771148
transform 1 0 85928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_925
timestamp 1670771148
transform 1 0 86204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_943
timestamp 1670771148
transform 1 0 87860 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1670771148
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1670771148
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1670771148
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1670771148
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_981
timestamp 1670771148
transform 1 0 91356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1003
timestamp 1670771148
transform 1 0 93380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1009
timestamp 1670771148
transform 1 0 93932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1021
timestamp 1670771148
transform 1 0 95036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1033
timestamp 1670771148
transform 1 0 96140 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1670771148
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1670771148
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1670771148
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1670771148
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1670771148
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1670771148
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1670771148
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1670771148
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1670771148
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1670771148
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1670771148
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1670771148
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1149
timestamp 1670771148
transform 1 0 106812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1167
timestamp 1670771148
transform 1 0 108468 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1670771148
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1185
timestamp 1670771148
transform 1 0 110124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1191
timestamp 1670771148
transform 1 0 110676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1200
timestamp 1670771148
transform 1 0 111504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1205
timestamp 1670771148
transform 1 0 111964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1213
timestamp 1670771148
transform 1 0 112700 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1216
timestamp 1670771148
transform 1 0 112976 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1228
timestamp 1670771148
transform 1 0 114080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1232
timestamp 1670771148
transform 1 0 114448 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1238
timestamp 1670771148
transform 1 0 115000 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1244
timestamp 1670771148
transform 1 0 115552 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1258
timestamp 1670771148
transform 1 0 116840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1261
timestamp 1670771148
transform 1 0 117116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1269
timestamp 1670771148
transform 1 0 117852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1275
timestamp 1670771148
transform 1 0 118404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1281
timestamp 1670771148
transform 1 0 118956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1290
timestamp 1670771148
transform 1 0 119784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1311
timestamp 1670771148
transform 1 0 121716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1670771148
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1317
timestamp 1670771148
transform 1 0 122268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1324
timestamp 1670771148
transform 1 0 122912 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1346
timestamp 1670771148
transform 1 0 124936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1352
timestamp 1670771148
transform 1 0 125488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1358
timestamp 1670771148
transform 1 0 126040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1364
timestamp 1670771148
transform 1 0 126592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1370
timestamp 1670771148
transform 1 0 127144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1373
timestamp 1670771148
transform 1 0 127420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1377
timestamp 1670771148
transform 1 0 127788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1399
timestamp 1670771148
transform 1 0 129812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1405
timestamp 1670771148
transform 1 0 130364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1411
timestamp 1670771148
transform 1 0 130916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1417
timestamp 1670771148
transform 1 0 131468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1420
timestamp 1670771148
transform 1 0 131744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1426
timestamp 1670771148
transform 1 0 132296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1429
timestamp 1670771148
transform 1 0 132572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1437
timestamp 1670771148
transform 1 0 133308 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1443
timestamp 1670771148
transform 1 0 133860 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1449
timestamp 1670771148
transform 1 0 134412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1455
timestamp 1670771148
transform 1 0 134964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1473
timestamp 1670771148
transform 1 0 136620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1479
timestamp 1670771148
transform 1 0 137172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1670771148
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1485
timestamp 1670771148
transform 1 0 137724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1491
timestamp 1670771148
transform 1 0 138276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1497
timestamp 1670771148
transform 1 0 138828 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1503
timestamp 1670771148
transform 1 0 139380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1507
timestamp 1670771148
transform 1 0 139748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1514
timestamp 1670771148
transform 1 0 140392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1534
timestamp 1670771148
transform 1 0 142232 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1541
timestamp 1670771148
transform 1 0 142876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1559
timestamp 1670771148
transform 1 0 144532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1567
timestamp 1670771148
transform 1 0 145268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1584
timestamp 1670771148
transform 1 0 146832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1593
timestamp 1670771148
transform 1 0 147660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1597
timestamp 1670771148
transform 1 0 148028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1615
timestamp 1670771148
transform 1 0 149684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1623
timestamp 1670771148
transform 1 0 150420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1630
timestamp 1670771148
transform 1 0 151064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1637
timestamp 1670771148
transform 1 0 151708 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1644
timestamp 1670771148
transform 1 0 152352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1650
timestamp 1670771148
transform 1 0 152904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1653
timestamp 1670771148
transform 1 0 153180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1672
timestamp 1670771148
transform 1 0 154928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1681
timestamp 1670771148
transform 1 0 155756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1690
timestamp 1670771148
transform 1 0 156584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1697
timestamp 1670771148
transform 1 0 157228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1704
timestamp 1670771148
transform 1 0 157872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1709
timestamp 1670771148
transform 1 0 158332 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1670771148
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1670771148
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1670771148
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1670771148
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1670771148
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_48
timestamp 1670771148
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1670771148
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1670771148
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1670771148
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1670771148
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1670771148
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1670771148
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1670771148
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1670771148
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1670771148
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_128
timestamp 1670771148
transform 1 0 12880 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1670771148
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_144
timestamp 1670771148
transform 1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1670771148
transform 1 0 14904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1670771148
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_157
timestamp 1670771148
transform 1 0 15548 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1670771148
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1670771148
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1670771148
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_173
timestamp 1670771148
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1670771148
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1670771148
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_195
timestamp 1670771148
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_207
timestamp 1670771148
transform 1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1670771148
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1670771148
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1670771148
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_229
timestamp 1670771148
transform 1 0 22172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_241
timestamp 1670771148
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_253
timestamp 1670771148
transform 1 0 24380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1670771148
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1670771148
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1670771148
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1670771148
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_305
timestamp 1670771148
transform 1 0 29164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_311
timestamp 1670771148
transform 1 0 29716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp 1670771148
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_325
timestamp 1670771148
transform 1 0 31004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1670771148
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1670771148
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1670771148
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_361
timestamp 1670771148
transform 1 0 34316 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_381
timestamp 1670771148
transform 1 0 36156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1670771148
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1670771148
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_399
timestamp 1670771148
transform 1 0 37812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1670771148
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_408
timestamp 1670771148
transform 1 0 38640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_412
timestamp 1670771148
transform 1 0 39008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_429
timestamp 1670771148
transform 1 0 40572 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_435
timestamp 1670771148
transform 1 0 41124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_439
timestamp 1670771148
transform 1 0 41492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1670771148
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_449
timestamp 1670771148
transform 1 0 42412 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_457
timestamp 1670771148
transform 1 0 43148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_469
timestamp 1670771148
transform 1 0 44252 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_477
timestamp 1670771148
transform 1 0 44988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_480
timestamp 1670771148
transform 1 0 45264 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_488
timestamp 1670771148
transform 1 0 46000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_494
timestamp 1670771148
transform 1 0 46552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1670771148
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1670771148
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_517
timestamp 1670771148
transform 1 0 48668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_525
timestamp 1670771148
transform 1 0 49404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_533
timestamp 1670771148
transform 1 0 50140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_537
timestamp 1670771148
transform 1 0 50508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_541
timestamp 1670771148
transform 1 0 50876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_558
timestamp 1670771148
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_561
timestamp 1670771148
transform 1 0 52716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_565
timestamp 1670771148
transform 1 0 53084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_568
timestamp 1670771148
transform 1 0 53360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_574
timestamp 1670771148
transform 1 0 53912 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_582
timestamp 1670771148
transform 1 0 54648 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1670771148
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1670771148
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_609
timestamp 1670771148
transform 1 0 57132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1670771148
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1670771148
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_622
timestamp 1670771148
transform 1 0 58328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_628
timestamp 1670771148
transform 1 0 58880 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_636
timestamp 1670771148
transform 1 0 59616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_639
timestamp 1670771148
transform 1 0 59892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_645
timestamp 1670771148
transform 1 0 60444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_649
timestamp 1670771148
transform 1 0 60812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_661
timestamp 1670771148
transform 1 0 61916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_667
timestamp 1670771148
transform 1 0 62468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_670
timestamp 1670771148
transform 1 0 62744 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_673
timestamp 1670771148
transform 1 0 63020 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_678
timestamp 1670771148
transform 1 0 63480 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_693
timestamp 1670771148
transform 1 0 64860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_699
timestamp 1670771148
transform 1 0 65412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_705
timestamp 1670771148
transform 1 0 65964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_708
timestamp 1670771148
transform 1 0 66240 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_714
timestamp 1670771148
transform 1 0 66792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_718
timestamp 1670771148
transform 1 0 67160 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_726
timestamp 1670771148
transform 1 0 67896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_729
timestamp 1670771148
transform 1 0 68172 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_733
timestamp 1670771148
transform 1 0 68540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_745
timestamp 1670771148
transform 1 0 69644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_757
timestamp 1670771148
transform 1 0 70748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_782
timestamp 1670771148
transform 1 0 73048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_785
timestamp 1670771148
transform 1 0 73324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_791
timestamp 1670771148
transform 1 0 73876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_809
timestamp 1670771148
transform 1 0 75532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_815
timestamp 1670771148
transform 1 0 76084 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1670771148
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1670771148
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1670771148
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_841
timestamp 1670771148
transform 1 0 78476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_864
timestamp 1670771148
transform 1 0 80592 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_886
timestamp 1670771148
transform 1 0 82616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_892
timestamp 1670771148
transform 1 0 83168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_897
timestamp 1670771148
transform 1 0 83628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_905
timestamp 1670771148
transform 1 0 84364 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1670771148
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_921
timestamp 1670771148
transform 1 0 85836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_924
timestamp 1670771148
transform 1 0 86112 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_938
timestamp 1670771148
transform 1 0 87400 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_950
timestamp 1670771148
transform 1 0 88504 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1670771148
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1670771148
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_977
timestamp 1670771148
transform 1 0 90988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_999
timestamp 1670771148
transform 1 0 93012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1670771148
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1670771148
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1021
timestamp 1670771148
transform 1 0 95036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1041
timestamp 1670771148
transform 1 0 96876 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1047
timestamp 1670771148
transform 1 0 97428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1059
timestamp 1670771148
transform 1 0 98532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1670771148
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1670771148
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1670771148
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1670771148
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1670771148
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1670771148
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1670771148
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1670771148
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1670771148
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1670771148
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1670771148
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1670771148
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1670771148
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1177
timestamp 1670771148
transform 1 0 109388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1185
timestamp 1670771148
transform 1 0 110124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1194
timestamp 1670771148
transform 1 0 110952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1214
timestamp 1670771148
transform 1 0 112792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1220
timestamp 1670771148
transform 1 0 113344 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1229
timestamp 1670771148
transform 1 0 114172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1670771148
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1245
timestamp 1670771148
transform 1 0 115644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1253
timestamp 1670771148
transform 1 0 116380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1258
timestamp 1670771148
transform 1 0 116840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1266
timestamp 1670771148
transform 1 0 117576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1286
timestamp 1670771148
transform 1 0 119416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1289
timestamp 1670771148
transform 1 0 119692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1308
timestamp 1670771148
transform 1 0 121440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1328
timestamp 1670771148
transform 1 0 123280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1334
timestamp 1670771148
transform 1 0 123832 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1342
timestamp 1670771148
transform 1 0 124568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1345
timestamp 1670771148
transform 1 0 124844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1351
timestamp 1670771148
transform 1 0 125396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1354
timestamp 1670771148
transform 1 0 125672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1360
timestamp 1670771148
transform 1 0 126224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1366
timestamp 1670771148
transform 1 0 126776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1372
timestamp 1670771148
transform 1 0 127328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1381
timestamp 1670771148
transform 1 0 128156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1389
timestamp 1670771148
transform 1 0 128892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1395
timestamp 1670771148
transform 1 0 129444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1670771148
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1401
timestamp 1670771148
transform 1 0 129996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1406
timestamp 1670771148
transform 1 0 130456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1412
timestamp 1670771148
transform 1 0 131008 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1422
timestamp 1670771148
transform 1 0 131928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1428
timestamp 1670771148
transform 1 0 132480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1434
timestamp 1670771148
transform 1 0 133032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1454
timestamp 1670771148
transform 1 0 134872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1457
timestamp 1670771148
transform 1 0 135148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1462
timestamp 1670771148
transform 1 0 135608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1468
timestamp 1670771148
transform 1 0 136160 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1474
timestamp 1670771148
transform 1 0 136712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1480
timestamp 1670771148
transform 1 0 137264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1486
timestamp 1670771148
transform 1 0 137816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1495
timestamp 1670771148
transform 1 0 138644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1504
timestamp 1670771148
transform 1 0 139472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1510
timestamp 1670771148
transform 1 0 140024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1513
timestamp 1670771148
transform 1 0 140300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1522
timestamp 1670771148
transform 1 0 141128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1546
timestamp 1670771148
transform 1 0 143336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1566
timestamp 1670771148
transform 1 0 145176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1569
timestamp 1670771148
transform 1 0 145452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1575
timestamp 1670771148
transform 1 0 146004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1593
timestamp 1670771148
transform 1 0 147660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1615
timestamp 1670771148
transform 1 0 149684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1621
timestamp 1670771148
transform 1 0 150236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1625
timestamp 1670771148
transform 1 0 150604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1643
timestamp 1670771148
transform 1 0 152260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1657
timestamp 1670771148
transform 1 0 153548 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1668
timestamp 1670771148
transform 1 0 154560 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1677
timestamp 1670771148
transform 1 0 155388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1681
timestamp 1670771148
transform 1 0 155756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1688
timestamp 1670771148
transform 1 0 156400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1697
timestamp 1670771148
transform 1 0 157228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1704
timestamp 1670771148
transform 1 0 157872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1710
timestamp 1670771148
transform 1 0 158424 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1670771148
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1670771148
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1670771148
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1670771148
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_37
timestamp 1670771148
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1670771148
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_51
timestamp 1670771148
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_59
timestamp 1670771148
transform 1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1670771148
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1670771148
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1670771148
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1670771148
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1670771148
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1670771148
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1670771148
transform 1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1670771148
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1670771148
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1670771148
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_146
timestamp 1670771148
transform 1 0 14536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_155
timestamp 1670771148
transform 1 0 15364 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1670771148
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1670771148
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1670771148
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1670771148
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_201
timestamp 1670771148
transform 1 0 19596 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1670771148
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_227
timestamp 1670771148
transform 1 0 21988 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_231
timestamp 1670771148
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1670771148
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1670771148
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1670771148
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1670771148
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_272
timestamp 1670771148
transform 1 0 26128 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_284
timestamp 1670771148
transform 1 0 27232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_296
timestamp 1670771148
transform 1 0 28336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1670771148
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_321
timestamp 1670771148
transform 1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_327
timestamp 1670771148
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_334
timestamp 1670771148
transform 1 0 31832 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_342
timestamp 1670771148
transform 1 0 32568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1670771148
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1670771148
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_371
timestamp 1670771148
transform 1 0 35236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_375
timestamp 1670771148
transform 1 0 35604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_383
timestamp 1670771148
transform 1 0 36340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_390
timestamp 1670771148
transform 1 0 36984 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_396
timestamp 1670771148
transform 1 0 37536 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_399
timestamp 1670771148
transform 1 0 37812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_408
timestamp 1670771148
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_412
timestamp 1670771148
transform 1 0 39008 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1670771148
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1670771148
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_428
timestamp 1670771148
transform 1 0 40480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_434
timestamp 1670771148
transform 1 0 41032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_454
timestamp 1670771148
transform 1 0 42872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_474
timestamp 1670771148
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp 1670771148
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_482
timestamp 1670771148
transform 1 0 45448 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_491
timestamp 1670771148
transform 1 0 46276 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_497
timestamp 1670771148
transform 1 0 46828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_506
timestamp 1670771148
transform 1 0 47656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1670771148
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_518
timestamp 1670771148
transform 1 0 48760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_524
timestamp 1670771148
transform 1 0 49312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_530
timestamp 1670771148
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_533
timestamp 1670771148
transform 1 0 50140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_538
timestamp 1670771148
transform 1 0 50600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_558
timestamp 1670771148
transform 1 0 52440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_565
timestamp 1670771148
transform 1 0 53084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_573
timestamp 1670771148
transform 1 0 53820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_579
timestamp 1670771148
transform 1 0 54372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_586
timestamp 1670771148
transform 1 0 55016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_589
timestamp 1670771148
transform 1 0 55292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_593
timestamp 1670771148
transform 1 0 55660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_596
timestamp 1670771148
transform 1 0 55936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1670771148
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_608
timestamp 1670771148
transform 1 0 57040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_628
timestamp 1670771148
transform 1 0 58880 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_634
timestamp 1670771148
transform 1 0 59432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1670771148
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1670771148
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_645
timestamp 1670771148
transform 1 0 60444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_649
timestamp 1670771148
transform 1 0 60812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_669
timestamp 1670771148
transform 1 0 62652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_675
timestamp 1670771148
transform 1 0 63204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_692
timestamp 1670771148
transform 1 0 64768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_698
timestamp 1670771148
transform 1 0 65320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_701
timestamp 1670771148
transform 1 0 65596 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_707
timestamp 1670771148
transform 1 0 66148 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_715
timestamp 1670771148
transform 1 0 66884 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_718
timestamp 1670771148
transform 1 0 67160 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_738
timestamp 1670771148
transform 1 0 69000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_750
timestamp 1670771148
transform 1 0 70104 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1670771148
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_769
timestamp 1670771148
transform 1 0 71852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_773
timestamp 1670771148
transform 1 0 72220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_793
timestamp 1670771148
transform 1 0 74060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_802
timestamp 1670771148
transform 1 0 74888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_810
timestamp 1670771148
transform 1 0 75624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_813
timestamp 1670771148
transform 1 0 75900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_818
timestamp 1670771148
transform 1 0 76360 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_824
timestamp 1670771148
transform 1 0 76912 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_836
timestamp 1670771148
transform 1 0 78016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_848
timestamp 1670771148
transform 1 0 79120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_860
timestamp 1670771148
transform 1 0 80224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_866
timestamp 1670771148
transform 1 0 80776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_869
timestamp 1670771148
transform 1 0 81052 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_891
timestamp 1670771148
transform 1 0 83076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_903
timestamp 1670771148
transform 1 0 84180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_922
timestamp 1670771148
transform 1 0 85928 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_925
timestamp 1670771148
transform 1 0 86204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_934
timestamp 1670771148
transform 1 0 87032 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_943
timestamp 1670771148
transform 1 0 87860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_955
timestamp 1670771148
transform 1 0 88964 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_967
timestamp 1670771148
transform 1 0 90068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_972
timestamp 1670771148
transform 1 0 90528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_978
timestamp 1670771148
transform 1 0 91080 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_981
timestamp 1670771148
transform 1 0 91356 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_999
timestamp 1670771148
transform 1 0 93012 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1005
timestamp 1670771148
transform 1 0 93564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1011
timestamp 1670771148
transform 1 0 94116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1019
timestamp 1670771148
transform 1 0 94852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1025
timestamp 1670771148
transform 1 0 95404 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1033
timestamp 1670771148
transform 1 0 96140 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1670771148
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1049
timestamp 1670771148
transform 1 0 97612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1053
timestamp 1670771148
transform 1 0 97980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1073
timestamp 1670771148
transform 1 0 99820 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1079
timestamp 1670771148
transform 1 0 100372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1670771148
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1670771148
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1670771148
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1670771148
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1129
timestamp 1670771148
transform 1 0 104972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1140
timestamp 1670771148
transform 1 0 105984 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1670771148
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1670771148
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1173
timestamp 1670771148
transform 1 0 109020 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1190
timestamp 1670771148
transform 1 0 110584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1670771148
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1670771148
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1205
timestamp 1670771148
transform 1 0 111964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1211
timestamp 1670771148
transform 1 0 112516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1217
timestamp 1670771148
transform 1 0 113068 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1223
timestamp 1670771148
transform 1 0 113620 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1240
timestamp 1670771148
transform 1 0 115184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1246
timestamp 1670771148
transform 1 0 115736 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1252
timestamp 1670771148
transform 1 0 116288 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1258
timestamp 1670771148
transform 1 0 116840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1261
timestamp 1670771148
transform 1 0 117116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1270
timestamp 1670771148
transform 1 0 117944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1276
timestamp 1670771148
transform 1 0 118496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1282
timestamp 1670771148
transform 1 0 119048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1306
timestamp 1670771148
transform 1 0 121256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1312
timestamp 1670771148
transform 1 0 121808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1317
timestamp 1670771148
transform 1 0 122268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1323
timestamp 1670771148
transform 1 0 122820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1329
timestamp 1670771148
transform 1 0 123372 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1345
timestamp 1670771148
transform 1 0 124844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1349
timestamp 1670771148
transform 1 0 125212 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1352
timestamp 1670771148
transform 1 0 125488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1358
timestamp 1670771148
transform 1 0 126040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1364
timestamp 1670771148
transform 1 0 126592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1370
timestamp 1670771148
transform 1 0 127144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1373
timestamp 1670771148
transform 1 0 127420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1391
timestamp 1670771148
transform 1 0 129076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1397
timestamp 1670771148
transform 1 0 129628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1403
timestamp 1670771148
transform 1 0 130180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1412
timestamp 1670771148
transform 1 0 131008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1418
timestamp 1670771148
transform 1 0 131560 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1426
timestamp 1670771148
transform 1 0 132296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1429
timestamp 1670771148
transform 1 0 132572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1441
timestamp 1670771148
transform 1 0 133676 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1465
timestamp 1670771148
transform 1 0 135884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1471
timestamp 1670771148
transform 1 0 136436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1479
timestamp 1670771148
transform 1 0 137172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1482
timestamp 1670771148
transform 1 0 137448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1485
timestamp 1670771148
transform 1 0 137724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1490
timestamp 1670771148
transform 1 0 138184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1494
timestamp 1670771148
transform 1 0 138552 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1512
timestamp 1670771148
transform 1 0 140208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1521
timestamp 1670771148
transform 1 0 141036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1528
timestamp 1670771148
transform 1 0 141680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1538
timestamp 1670771148
transform 1 0 142600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1541
timestamp 1670771148
transform 1 0 142876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1559
timestamp 1670771148
transform 1 0 144532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1579
timestamp 1670771148
transform 1 0 146372 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1592
timestamp 1670771148
transform 1 0 147568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1597
timestamp 1670771148
transform 1 0 148028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1615
timestamp 1670771148
transform 1 0 149684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1623
timestamp 1670771148
transform 1 0 150420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1637
timestamp 1670771148
transform 1 0 151708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1646
timestamp 1670771148
transform 1 0 152536 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1653
timestamp 1670771148
transform 1 0 153180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1660
timestamp 1670771148
transform 1 0 153824 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1666
timestamp 1670771148
transform 1 0 154376 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1684
timestamp 1670771148
transform 1 0 156032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1693
timestamp 1670771148
transform 1 0 156860 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1700
timestamp 1670771148
transform 1 0 157504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1706
timestamp 1670771148
transform 1 0 158056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1709
timestamp 1670771148
transform 1 0 158332 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1670771148
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1670771148
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1670771148
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1670771148
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1670771148
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_46
timestamp 1670771148
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1670771148
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1670771148
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1670771148
transform 1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_70
timestamp 1670771148
transform 1 0 7544 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_82
timestamp 1670771148
transform 1 0 8648 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_94
timestamp 1670771148
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1670771148
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1670771148
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1670771148
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_138
timestamp 1670771148
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1670771148
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1670771148
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1670771148
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1670771148
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_176
timestamp 1670771148
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_183
timestamp 1670771148
transform 1 0 17940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1670771148
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1670771148
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_201
timestamp 1670771148
transform 1 0 19596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1670771148
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1670771148
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1670771148
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1670771148
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1670771148
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1670771148
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1670771148
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1670771148
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1670771148
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_299
timestamp 1670771148
transform 1 0 28612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1670771148
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_311
timestamp 1670771148
transform 1 0 29716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_317
timestamp 1670771148
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_326
timestamp 1670771148
transform 1 0 31096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1670771148
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_337
timestamp 1670771148
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_343
timestamp 1670771148
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_346
timestamp 1670771148
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_353
timestamp 1670771148
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_373
timestamp 1670771148
transform 1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_379
timestamp 1670771148
transform 1 0 35972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1670771148
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_393
timestamp 1670771148
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_404
timestamp 1670771148
transform 1 0 38272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_424
timestamp 1670771148
transform 1 0 40112 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_432
timestamp 1670771148
transform 1 0 40848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1670771148
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1670771148
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1670771148
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_467
timestamp 1670771148
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_474
timestamp 1670771148
transform 1 0 44712 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_496
timestamp 1670771148
transform 1 0 46736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1670771148
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_505
timestamp 1670771148
transform 1 0 47564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_511
timestamp 1670771148
transform 1 0 48116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_514
timestamp 1670771148
transform 1 0 48392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_521
timestamp 1670771148
transform 1 0 49036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_541
timestamp 1670771148
transform 1 0 50876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_549
timestamp 1670771148
transform 1 0 51612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1670771148
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_561
timestamp 1670771148
transform 1 0 52716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_567
timestamp 1670771148
transform 1 0 53268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_570
timestamp 1670771148
transform 1 0 53544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_590
timestamp 1670771148
transform 1 0 55384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_598
timestamp 1670771148
transform 1 0 56120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_605
timestamp 1670771148
transform 1 0 56764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1670771148
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_617
timestamp 1670771148
transform 1 0 57868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_635
timestamp 1670771148
transform 1 0 59524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_641
timestamp 1670771148
transform 1 0 60076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_650
timestamp 1670771148
transform 1 0 60904 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_656
timestamp 1670771148
transform 1 0 61456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_670
timestamp 1670771148
transform 1 0 62744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_673
timestamp 1670771148
transform 1 0 63020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_679
timestamp 1670771148
transform 1 0 63572 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_682
timestamp 1670771148
transform 1 0 63848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_706
timestamp 1670771148
transform 1 0 66056 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_714
timestamp 1670771148
transform 1 0 66792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_717
timestamp 1670771148
transform 1 0 67068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_726
timestamp 1670771148
transform 1 0 67896 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_729
timestamp 1670771148
transform 1 0 68172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_747
timestamp 1670771148
transform 1 0 69828 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1670771148
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1670771148
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1670771148
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1670771148
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_785
timestamp 1670771148
transform 1 0 73324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_789
timestamp 1670771148
transform 1 0 73692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_797
timestamp 1670771148
transform 1 0 74428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_801
timestamp 1670771148
transform 1 0 74796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_818
timestamp 1670771148
transform 1 0 76360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_838
timestamp 1670771148
transform 1 0 78200 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1670771148
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1670771148
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1670771148
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1670771148
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1670771148
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1670771148
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_897
timestamp 1670771148
transform 1 0 83628 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_902
timestamp 1670771148
transform 1 0 84088 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_914
timestamp 1670771148
transform 1 0 85192 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_926
timestamp 1670771148
transform 1 0 86296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_930
timestamp 1670771148
transform 1 0 86664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_947
timestamp 1670771148
transform 1 0 88228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1670771148
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_953
timestamp 1670771148
transform 1 0 88780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_971
timestamp 1670771148
transform 1 0 90436 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_991
timestamp 1670771148
transform 1 0 92276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_997
timestamp 1670771148
transform 1 0 92828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1003
timestamp 1670771148
transform 1 0 93380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1670771148
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1009
timestamp 1670771148
transform 1 0 93932 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1016
timestamp 1670771148
transform 1 0 94576 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1028
timestamp 1670771148
transform 1 0 95680 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1040
timestamp 1670771148
transform 1 0 96784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1052
timestamp 1670771148
transform 1 0 97888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1670771148
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1670771148
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1670771148
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1670771148
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1670771148
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1670771148
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1670771148
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1670771148
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1670771148
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1670771148
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1145
timestamp 1670771148
transform 1 0 106444 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1153
timestamp 1670771148
transform 1 0 107180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1161
timestamp 1670771148
transform 1 0 107916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1166
timestamp 1670771148
transform 1 0 108376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1173
timestamp 1670771148
transform 1 0 109020 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1177
timestamp 1670771148
transform 1 0 109388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1195
timestamp 1670771148
transform 1 0 111044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1201
timestamp 1670771148
transform 1 0 111596 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1209
timestamp 1670771148
transform 1 0 112332 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1215
timestamp 1670771148
transform 1 0 112884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1227
timestamp 1670771148
transform 1 0 113988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1670771148
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1233
timestamp 1670771148
transform 1 0 114540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1239
timestamp 1670771148
transform 1 0 115092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1242
timestamp 1670771148
transform 1 0 115368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1248
timestamp 1670771148
transform 1 0 115920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1254
timestamp 1670771148
transform 1 0 116472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1260
timestamp 1670771148
transform 1 0 117024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1266
timestamp 1670771148
transform 1 0 117576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1275
timestamp 1670771148
transform 1 0 118404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1284
timestamp 1670771148
transform 1 0 119232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1289
timestamp 1670771148
transform 1 0 119692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1293
timestamp 1670771148
transform 1 0 120060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1313
timestamp 1670771148
transform 1 0 121900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1317
timestamp 1670771148
transform 1 0 122268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1321
timestamp 1670771148
transform 1 0 122636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1341
timestamp 1670771148
transform 1 0 124476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1345
timestamp 1670771148
transform 1 0 124844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1349
timestamp 1670771148
transform 1 0 125212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1367
timestamp 1670771148
transform 1 0 126868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1373
timestamp 1670771148
transform 1 0 127420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1381
timestamp 1670771148
transform 1 0 128156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1395
timestamp 1670771148
transform 1 0 129444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1670771148
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1401
timestamp 1670771148
transform 1 0 129996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1408
timestamp 1670771148
transform 1 0 130640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1414
timestamp 1670771148
transform 1 0 131192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1434
timestamp 1670771148
transform 1 0 133032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1454
timestamp 1670771148
transform 1 0 134872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1457
timestamp 1670771148
transform 1 0 135148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1465
timestamp 1670771148
transform 1 0 135884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1471
timestamp 1670771148
transform 1 0 136436 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1477
timestamp 1670771148
transform 1 0 136988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1483
timestamp 1670771148
transform 1 0 137540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1489
timestamp 1670771148
transform 1 0 138092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1495
timestamp 1670771148
transform 1 0 138644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1501
timestamp 1670771148
transform 1 0 139196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1504
timestamp 1670771148
transform 1 0 139472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1510
timestamp 1670771148
transform 1 0 140024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1513
timestamp 1670771148
transform 1 0 140300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1518
timestamp 1670771148
transform 1 0 140760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1525
timestamp 1670771148
transform 1 0 141404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1545
timestamp 1670771148
transform 1 0 143244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1565
timestamp 1670771148
transform 1 0 145084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1569
timestamp 1670771148
transform 1 0 145452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1587
timestamp 1670771148
transform 1 0 147108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1607
timestamp 1670771148
transform 1 0 148948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1616
timestamp 1670771148
transform 1 0 149776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1622
timestamp 1670771148
transform 1 0 150328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1625
timestamp 1670771148
transform 1 0 150604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1630
timestamp 1670771148
transform 1 0 151064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1644
timestamp 1670771148
transform 1 0 152352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1654
timestamp 1670771148
transform 1 0 153272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1663
timestamp 1670771148
transform 1 0 154100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1672
timestamp 1670771148
transform 1 0 154928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1678
timestamp 1670771148
transform 1 0 155480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1681
timestamp 1670771148
transform 1 0 155756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1688
timestamp 1670771148
transform 1 0 156400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1697
timestamp 1670771148
transform 1 0 157228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1705
timestamp 1670771148
transform 1 0 157964 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1710
timestamp 1670771148
transform 1 0 158424 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1670771148
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1670771148
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1670771148
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1670771148
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_47
timestamp 1670771148
transform 1 0 5428 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1670771148
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1670771148
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1670771148
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1670771148
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1670771148
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1670771148
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_103
timestamp 1670771148
transform 1 0 10580 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_106
timestamp 1670771148
transform 1 0 10856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_115
timestamp 1670771148
transform 1 0 11684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1670771148
transform 1 0 12236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1670771148
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1670771148
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1670771148
transform 1 0 14720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1670771148
transform 1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1670771148
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1670771148
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1670771148
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1670771148
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1670771148
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1670771148
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1670771148
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1670771148
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1670771148
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1670771148
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1670771148
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1670771148
transform 1 0 26220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_277
timestamp 1670771148
transform 1 0 26588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_286
timestamp 1670771148
transform 1 0 27416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1670771148
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1670771148
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_327
timestamp 1670771148
transform 1 0 31188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_349
timestamp 1670771148
transform 1 0 33212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1670771148
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1670771148
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_371
timestamp 1670771148
transform 1 0 35236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_388
timestamp 1670771148
transform 1 0 36800 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_408
timestamp 1670771148
transform 1 0 38640 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1670771148
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_421
timestamp 1670771148
transform 1 0 39836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_443
timestamp 1670771148
transform 1 0 41860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_449
timestamp 1670771148
transform 1 0 42412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_466
timestamp 1670771148
transform 1 0 43976 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1670771148
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1670771148
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_482
timestamp 1670771148
transform 1 0 45448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_502
timestamp 1670771148
transform 1 0 47288 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1670771148
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_518
timestamp 1670771148
transform 1 0 48760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_524
timestamp 1670771148
transform 1 0 49312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_530
timestamp 1670771148
transform 1 0 49864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_533
timestamp 1670771148
transform 1 0 50140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_555
timestamp 1670771148
transform 1 0 52164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_563
timestamp 1670771148
transform 1 0 52900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_571
timestamp 1670771148
transform 1 0 53636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_577
timestamp 1670771148
transform 1 0 54188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_583
timestamp 1670771148
transform 1 0 54740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1670771148
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_589
timestamp 1670771148
transform 1 0 55292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_595
timestamp 1670771148
transform 1 0 55844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_602
timestamp 1670771148
transform 1 0 56488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_611
timestamp 1670771148
transform 1 0 57316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_631
timestamp 1670771148
transform 1 0 59156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1670771148
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1670771148
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_645
timestamp 1670771148
transform 1 0 60444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_650
timestamp 1670771148
transform 1 0 60904 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_656
timestamp 1670771148
transform 1 0 61456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_659
timestamp 1670771148
transform 1 0 61732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_680
timestamp 1670771148
transform 1 0 63664 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_688
timestamp 1670771148
transform 1 0 64400 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_691
timestamp 1670771148
transform 1 0 64676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_695
timestamp 1670771148
transform 1 0 65044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_698
timestamp 1670771148
transform 1 0 65320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_701
timestamp 1670771148
transform 1 0 65596 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_719
timestamp 1670771148
transform 1 0 67252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_727
timestamp 1670771148
transform 1 0 67988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_732
timestamp 1670771148
transform 1 0 68448 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_738
timestamp 1670771148
transform 1 0 69000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_750
timestamp 1670771148
transform 1 0 70104 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1670771148
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1670771148
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1670771148
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_793
timestamp 1670771148
transform 1 0 74060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_798
timestamp 1670771148
transform 1 0 74520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1670771148
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1670771148
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_813
timestamp 1670771148
transform 1 0 75900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_820
timestamp 1670771148
transform 1 0 76544 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_826
timestamp 1670771148
transform 1 0 77096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_838
timestamp 1670771148
transform 1 0 78200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_850
timestamp 1670771148
transform 1 0 79304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_862
timestamp 1670771148
transform 1 0 80408 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1670771148
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1670771148
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1670771148
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1670771148
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1670771148
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1670771148
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_925
timestamp 1670771148
transform 1 0 86204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_943
timestamp 1670771148
transform 1 0 87860 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_949
timestamp 1670771148
transform 1 0 88412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_955
timestamp 1670771148
transform 1 0 88964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_976
timestamp 1670771148
transform 1 0 90896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_981
timestamp 1670771148
transform 1 0 91356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_999
timestamp 1670771148
transform 1 0 93012 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1019
timestamp 1670771148
transform 1 0 94852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1031
timestamp 1670771148
transform 1 0 95956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1034
timestamp 1670771148
transform 1 0 96232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1037
timestamp 1670771148
transform 1 0 96508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1055
timestamp 1670771148
transform 1 0 98164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1061
timestamp 1670771148
transform 1 0 98716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1067
timestamp 1670771148
transform 1 0 99268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1084
timestamp 1670771148
transform 1 0 100832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1090
timestamp 1670771148
transform 1 0 101384 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1670771148
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1670771148
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1117
timestamp 1670771148
transform 1 0 103868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1123
timestamp 1670771148
transform 1 0 104420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1127
timestamp 1670771148
transform 1 0 104788 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1130
timestamp 1670771148
transform 1 0 105064 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1142
timestamp 1670771148
transform 1 0 106168 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1149
timestamp 1670771148
transform 1 0 106812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1160
timestamp 1670771148
transform 1 0 107824 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1167
timestamp 1670771148
transform 1 0 108468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1179
timestamp 1670771148
transform 1 0 109572 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1191
timestamp 1670771148
transform 1 0 110676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1196
timestamp 1670771148
transform 1 0 111136 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1205
timestamp 1670771148
transform 1 0 111964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1213
timestamp 1670771148
transform 1 0 112700 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1219
timestamp 1670771148
transform 1 0 113252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1231
timestamp 1670771148
transform 1 0 114356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1235
timestamp 1670771148
transform 1 0 114724 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1238
timestamp 1670771148
transform 1 0 115000 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1244
timestamp 1670771148
transform 1 0 115552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1250
timestamp 1670771148
transform 1 0 116104 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1258
timestamp 1670771148
transform 1 0 116840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1261
timestamp 1670771148
transform 1 0 117116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1265
timestamp 1670771148
transform 1 0 117484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1269
timestamp 1670771148
transform 1 0 117852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1273
timestamp 1670771148
transform 1 0 118220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1279
timestamp 1670771148
transform 1 0 118772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1285
timestamp 1670771148
transform 1 0 119324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1290
timestamp 1670771148
transform 1 0 119784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1296
timestamp 1670771148
transform 1 0 120336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1302
timestamp 1670771148
transform 1 0 120888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1308
timestamp 1670771148
transform 1 0 121440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1314
timestamp 1670771148
transform 1 0 121992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1317
timestamp 1670771148
transform 1 0 122268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1324
timestamp 1670771148
transform 1 0 122912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1330
timestamp 1670771148
transform 1 0 123464 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1336
timestamp 1670771148
transform 1 0 124016 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1339
timestamp 1670771148
transform 1 0 124292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1345
timestamp 1670771148
transform 1 0 124844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1351
timestamp 1670771148
transform 1 0 125396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1357
timestamp 1670771148
transform 1 0 125948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1363
timestamp 1670771148
transform 1 0 126500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1369
timestamp 1670771148
transform 1 0 127052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1373
timestamp 1670771148
transform 1 0 127420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1377
timestamp 1670771148
transform 1 0 127788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1385
timestamp 1670771148
transform 1 0 128524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1388
timestamp 1670771148
transform 1 0 128800 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1408
timestamp 1670771148
transform 1 0 130640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1414
timestamp 1670771148
transform 1 0 131192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1420
timestamp 1670771148
transform 1 0 131744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1426
timestamp 1670771148
transform 1 0 132296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1429
timestamp 1670771148
transform 1 0 132572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1436
timestamp 1670771148
transform 1 0 133216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1442
timestamp 1670771148
transform 1 0 133768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1448
timestamp 1670771148
transform 1 0 134320 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1458
timestamp 1670771148
transform 1 0 135240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1466
timestamp 1670771148
transform 1 0 135976 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1472
timestamp 1670771148
transform 1 0 136528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1482
timestamp 1670771148
transform 1 0 137448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1485
timestamp 1670771148
transform 1 0 137724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1491
timestamp 1670771148
transform 1 0 138276 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1497
timestamp 1670771148
transform 1 0 138828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1503
timestamp 1670771148
transform 1 0 139380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1509
timestamp 1670771148
transform 1 0 139932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1516
timestamp 1670771148
transform 1 0 140576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1524
timestamp 1670771148
transform 1 0 141312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1538
timestamp 1670771148
transform 1 0 142600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1541
timestamp 1670771148
transform 1 0 142876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1559
timestamp 1670771148
transform 1 0 144532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1565
timestamp 1670771148
transform 1 0 145084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1587
timestamp 1670771148
transform 1 0 147108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1593
timestamp 1670771148
transform 1 0 147660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1597
timestamp 1670771148
transform 1 0 148028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1601
timestamp 1670771148
transform 1 0 148396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1621
timestamp 1670771148
transform 1 0 150236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1630
timestamp 1670771148
transform 1 0 151064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1639
timestamp 1670771148
transform 1 0 151892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1648
timestamp 1670771148
transform 1 0 152720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1653
timestamp 1670771148
transform 1 0 153180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1660
timestamp 1670771148
transform 1 0 153824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1669
timestamp 1670771148
transform 1 0 154652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1678
timestamp 1670771148
transform 1 0 155480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1687
timestamp 1670771148
transform 1 0 156308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1696
timestamp 1670771148
transform 1 0 157136 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1703
timestamp 1670771148
transform 1 0 157780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1707
timestamp 1670771148
transform 1 0 158148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1709
timestamp 1670771148
transform 1 0 158332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1670771148
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1670771148
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_19
timestamp 1670771148
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1670771148
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 1670771148
transform 1 0 5336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1670771148
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1670771148
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1670771148
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1670771148
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1670771148
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1670771148
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1670771148
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1670771148
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1670771148
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1670771148
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_127
timestamp 1670771148
transform 1 0 12788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1670771148
transform 1 0 14996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_160
timestamp 1670771148
transform 1 0 15824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1670771148
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1670771148
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1670771148
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1670771148
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1670771148
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1670771148
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1670771148
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1670771148
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1670771148
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1670771148
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1670771148
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_257
timestamp 1670771148
transform 1 0 24748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1670771148
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1670771148
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_281
timestamp 1670771148
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1670771148
transform 1 0 28704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_320
timestamp 1670771148
transform 1 0 30544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_326
timestamp 1670771148
transform 1 0 31096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1670771148
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_337
timestamp 1670771148
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1670771148
transform 1 0 34132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_383
timestamp 1670771148
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_387
timestamp 1670771148
transform 1 0 36708 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1670771148
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_393
timestamp 1670771148
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_412
timestamp 1670771148
transform 1 0 39008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_420
timestamp 1670771148
transform 1 0 39744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_426
timestamp 1670771148
transform 1 0 40296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1670771148
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1670771148
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_453
timestamp 1670771148
transform 1 0 42780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_473
timestamp 1670771148
transform 1 0 44620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_480
timestamp 1670771148
transform 1 0 45264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_484
timestamp 1670771148
transform 1 0 45632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_487
timestamp 1670771148
transform 1 0 45908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_493
timestamp 1670771148
transform 1 0 46460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1670771148
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_505
timestamp 1670771148
transform 1 0 47564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_511
timestamp 1670771148
transform 1 0 48116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_517
timestamp 1670771148
transform 1 0 48668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_525
timestamp 1670771148
transform 1 0 49404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_533
timestamp 1670771148
transform 1 0 50140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_550
timestamp 1670771148
transform 1 0 51704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_558
timestamp 1670771148
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_561
timestamp 1670771148
transform 1 0 52716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_579
timestamp 1670771148
transform 1 0 54372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_590
timestamp 1670771148
transform 1 0 55384 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_599
timestamp 1670771148
transform 1 0 56212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_607
timestamp 1670771148
transform 1 0 56948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1670771148
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_617
timestamp 1670771148
transform 1 0 57868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_625
timestamp 1670771148
transform 1 0 58604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_649
timestamp 1670771148
transform 1 0 60812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_659
timestamp 1670771148
transform 1 0 61732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1670771148
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1670771148
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_673
timestamp 1670771148
transform 1 0 63020 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_682
timestamp 1670771148
transform 1 0 63848 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_690
timestamp 1670771148
transform 1 0 64584 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_696
timestamp 1670771148
transform 1 0 65136 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_702
timestamp 1670771148
transform 1 0 65688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_708
timestamp 1670771148
transform 1 0 66240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_714
timestamp 1670771148
transform 1 0 66792 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_720
timestamp 1670771148
transform 1 0 67344 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_724
timestamp 1670771148
transform 1 0 67712 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1670771148
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1670771148
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1670771148
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1670771148
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_777
timestamp 1670771148
transform 1 0 72588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_782
timestamp 1670771148
transform 1 0 73048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_785
timestamp 1670771148
transform 1 0 73324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_792
timestamp 1670771148
transform 1 0 73968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_798
timestamp 1670771148
transform 1 0 74520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_801
timestamp 1670771148
transform 1 0 74796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_821
timestamp 1670771148
transform 1 0 76636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_828
timestamp 1670771148
transform 1 0 77280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_834
timestamp 1670771148
transform 1 0 77832 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1670771148
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_853
timestamp 1670771148
transform 1 0 79580 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_857
timestamp 1670771148
transform 1 0 79948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_869
timestamp 1670771148
transform 1 0 81052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_881
timestamp 1670771148
transform 1 0 82156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_889
timestamp 1670771148
transform 1 0 82892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_894
timestamp 1670771148
transform 1 0 83352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_897
timestamp 1670771148
transform 1 0 83628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_915
timestamp 1670771148
transform 1 0 85284 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1670771148
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1670771148
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_945
timestamp 1670771148
transform 1 0 88044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_950
timestamp 1670771148
transform 1 0 88504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_953
timestamp 1670771148
transform 1 0 88780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_972
timestamp 1670771148
transform 1 0 90528 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_992
timestamp 1670771148
transform 1 0 92368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1006
timestamp 1670771148
transform 1 0 93656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1009
timestamp 1670771148
transform 1 0 93932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1030
timestamp 1670771148
transform 1 0 95864 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1036
timestamp 1670771148
transform 1 0 96416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1048
timestamp 1670771148
transform 1 0 97520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1053
timestamp 1670771148
transform 1 0 97980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1062
timestamp 1670771148
transform 1 0 98808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1065
timestamp 1670771148
transform 1 0 99084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1084
timestamp 1670771148
transform 1 0 100832 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1090
timestamp 1670771148
transform 1 0 101384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1102
timestamp 1670771148
transform 1 0 102488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1110
timestamp 1670771148
transform 1 0 103224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1670771148
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1670771148
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1121
timestamp 1670771148
transform 1 0 104236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1128
timestamp 1670771148
transform 1 0 104880 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1137
timestamp 1670771148
transform 1 0 105708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1149
timestamp 1670771148
transform 1 0 106812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1155
timestamp 1670771148
transform 1 0 107364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1163
timestamp 1670771148
transform 1 0 108100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1670771148
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1670771148
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1177
timestamp 1670771148
transform 1 0 109388 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1185
timestamp 1670771148
transform 1 0 110124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1197
timestamp 1670771148
transform 1 0 111228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1670771148
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1215
timestamp 1670771148
transform 1 0 112884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1224
timestamp 1670771148
transform 1 0 113712 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1230
timestamp 1670771148
transform 1 0 114264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1233
timestamp 1670771148
transform 1 0 114540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1237
timestamp 1670771148
transform 1 0 114908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1241
timestamp 1670771148
transform 1 0 115276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1259
timestamp 1670771148
transform 1 0 116932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1263
timestamp 1670771148
transform 1 0 117300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1266
timestamp 1670771148
transform 1 0 117576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1272
timestamp 1670771148
transform 1 0 118128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1275
timestamp 1670771148
transform 1 0 118404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1281
timestamp 1670771148
transform 1 0 118956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1287
timestamp 1670771148
transform 1 0 119508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1289
timestamp 1670771148
transform 1 0 119692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1293
timestamp 1670771148
transform 1 0 120060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1301
timestamp 1670771148
transform 1 0 120796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1304
timestamp 1670771148
transform 1 0 121072 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1328
timestamp 1670771148
transform 1 0 123280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1334
timestamp 1670771148
transform 1 0 123832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1342
timestamp 1670771148
transform 1 0 124568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1345
timestamp 1670771148
transform 1 0 124844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1349
timestamp 1670771148
transform 1 0 125212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1355
timestamp 1670771148
transform 1 0 125764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1361
timestamp 1670771148
transform 1 0 126316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1367
timestamp 1670771148
transform 1 0 126868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1375
timestamp 1670771148
transform 1 0 127604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1378
timestamp 1670771148
transform 1 0 127880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1398
timestamp 1670771148
transform 1 0 129720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1401
timestamp 1670771148
transform 1 0 129996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1405
timestamp 1670771148
transform 1 0 130364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1413
timestamp 1670771148
transform 1 0 131100 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1430
timestamp 1670771148
transform 1 0 132664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1454
timestamp 1670771148
transform 1 0 134872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1457
timestamp 1670771148
transform 1 0 135148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1461
timestamp 1670771148
transform 1 0 135516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1464
timestamp 1670771148
transform 1 0 135792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1468
timestamp 1670771148
transform 1 0 136160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1471
timestamp 1670771148
transform 1 0 136436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1477
timestamp 1670771148
transform 1 0 136988 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1483
timestamp 1670771148
transform 1 0 137540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1503
timestamp 1670771148
transform 1 0 139380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1509
timestamp 1670771148
transform 1 0 139932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1513
timestamp 1670771148
transform 1 0 140300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1517
timestamp 1670771148
transform 1 0 140668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1523
timestamp 1670771148
transform 1 0 141220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1529
timestamp 1670771148
transform 1 0 141772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1546
timestamp 1670771148
transform 1 0 143336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1566
timestamp 1670771148
transform 1 0 145176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1569
timestamp 1670771148
transform 1 0 145452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1588
timestamp 1670771148
transform 1 0 147200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1608
timestamp 1670771148
transform 1 0 149040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1617
timestamp 1670771148
transform 1 0 149868 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1623
timestamp 1670771148
transform 1 0 150420 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1625
timestamp 1670771148
transform 1 0 150604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1631
timestamp 1670771148
transform 1 0 151156 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1648
timestamp 1670771148
transform 1 0 152720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1657
timestamp 1670771148
transform 1 0 153548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1666
timestamp 1670771148
transform 1 0 154376 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1675
timestamp 1670771148
transform 1 0 155204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1679
timestamp 1670771148
transform 1 0 155572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1681
timestamp 1670771148
transform 1 0 155756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1688
timestamp 1670771148
transform 1 0 156400 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1697
timestamp 1670771148
transform 1 0 157228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1704
timestamp 1670771148
transform 1 0 157872 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1710
timestamp 1670771148
transform 1 0 158424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1670771148
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1670771148
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1670771148
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1670771148
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1670771148
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1670771148
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1670771148
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1670771148
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1670771148
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1670771148
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1670771148
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1670771148
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1670771148
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_108
timestamp 1670771148
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_117
timestamp 1670771148
transform 1 0 11868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_123
timestamp 1670771148
transform 1 0 12420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1670771148
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1670771148
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1670771148
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1670771148
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1670771148
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_163
timestamp 1670771148
transform 1 0 16100 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1670771148
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_173
timestamp 1670771148
transform 1 0 17020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1670771148
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1670771148
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1670771148
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1670771148
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1670771148
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1670771148
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_208
timestamp 1670771148
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_220
timestamp 1670771148
transform 1 0 21344 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1670771148
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1670771148
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_253
timestamp 1670771148
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_261
timestamp 1670771148
transform 1 0 25116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_266
timestamp 1670771148
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1670771148
transform 1 0 27416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1670771148
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1670771148
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_328
timestamp 1670771148
transform 1 0 31280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1670771148
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 1670771148
transform 1 0 32844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_349
timestamp 1670771148
transform 1 0 33212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_355
timestamp 1670771148
transform 1 0 33764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1670771148
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1670771148
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_369
timestamp 1670771148
transform 1 0 35052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_375
timestamp 1670771148
transform 1 0 35604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_378
timestamp 1670771148
transform 1 0 35880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_398
timestamp 1670771148
transform 1 0 37720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_404
timestamp 1670771148
transform 1 0 38272 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_412
timestamp 1670771148
transform 1 0 39008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1670771148
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_421
timestamp 1670771148
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_427
timestamp 1670771148
transform 1 0 40388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_434
timestamp 1670771148
transform 1 0 41032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_454
timestamp 1670771148
transform 1 0 42872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1670771148
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_477
timestamp 1670771148
transform 1 0 44988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_481
timestamp 1670771148
transform 1 0 45356 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_484
timestamp 1670771148
transform 1 0 45632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_492
timestamp 1670771148
transform 1 0 46368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_501
timestamp 1670771148
transform 1 0 47196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_505
timestamp 1670771148
transform 1 0 47564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_510
timestamp 1670771148
transform 1 0 48024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_530
timestamp 1670771148
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_533
timestamp 1670771148
transform 1 0 50140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_539
timestamp 1670771148
transform 1 0 50692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_547
timestamp 1670771148
transform 1 0 51428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_556
timestamp 1670771148
transform 1 0 52256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_576
timestamp 1670771148
transform 1 0 54096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_585
timestamp 1670771148
transform 1 0 54924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_589
timestamp 1670771148
transform 1 0 55292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_593
timestamp 1670771148
transform 1 0 55660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_601
timestamp 1670771148
transform 1 0 56396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_610
timestamp 1670771148
transform 1 0 57224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_618
timestamp 1670771148
transform 1 0 57960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_626
timestamp 1670771148
transform 1 0 58696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_631
timestamp 1670771148
transform 1 0 59156 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_637
timestamp 1670771148
transform 1 0 59708 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_642
timestamp 1670771148
transform 1 0 60168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_645
timestamp 1670771148
transform 1 0 60444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_663
timestamp 1670771148
transform 1 0 62100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_669
timestamp 1670771148
transform 1 0 62652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_678
timestamp 1670771148
transform 1 0 63480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_698
timestamp 1670771148
transform 1 0 65320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_701
timestamp 1670771148
transform 1 0 65596 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_719
timestamp 1670771148
transform 1 0 67252 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_731
timestamp 1670771148
transform 1 0 68356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_743
timestamp 1670771148
transform 1 0 69460 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_746
timestamp 1670771148
transform 1 0 69736 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_754
timestamp 1670771148
transform 1 0 70472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_757
timestamp 1670771148
transform 1 0 70748 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_763
timestamp 1670771148
transform 1 0 71300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_775
timestamp 1670771148
transform 1 0 72404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_779
timestamp 1670771148
transform 1 0 72772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_785
timestamp 1670771148
transform 1 0 73324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1670771148
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1670771148
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_813
timestamp 1670771148
transform 1 0 75900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_820
timestamp 1670771148
transform 1 0 76544 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_826
timestamp 1670771148
transform 1 0 77096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_829
timestamp 1670771148
transform 1 0 77372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_835
timestamp 1670771148
transform 1 0 77924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_855
timestamp 1670771148
transform 1 0 79764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_863
timestamp 1670771148
transform 1 0 80500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_866
timestamp 1670771148
transform 1 0 80776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_869
timestamp 1670771148
transform 1 0 81052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_887
timestamp 1670771148
transform 1 0 82708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_893
timestamp 1670771148
transform 1 0 83260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_904
timestamp 1670771148
transform 1 0 84272 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_912
timestamp 1670771148
transform 1 0 85008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_920
timestamp 1670771148
transform 1 0 85744 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1670771148
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_939
timestamp 1670771148
transform 1 0 87492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_959
timestamp 1670771148
transform 1 0 89332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_965
timestamp 1670771148
transform 1 0 89884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_971
timestamp 1670771148
transform 1 0 90436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_977
timestamp 1670771148
transform 1 0 90988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_981
timestamp 1670771148
transform 1 0 91356 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_985
timestamp 1670771148
transform 1 0 91724 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_989
timestamp 1670771148
transform 1 0 92092 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_992
timestamp 1670771148
transform 1 0 92368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1013
timestamp 1670771148
transform 1 0 94300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1017
timestamp 1670771148
transform 1 0 94668 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1034
timestamp 1670771148
transform 1 0 96232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1037
timestamp 1670771148
transform 1 0 96508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1045
timestamp 1670771148
transform 1 0 97244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1054
timestamp 1670771148
transform 1 0 98072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1078
timestamp 1670771148
transform 1 0 100280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1084
timestamp 1670771148
transform 1 0 100832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1090
timestamp 1670771148
transform 1 0 101384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1093
timestamp 1670771148
transform 1 0 101660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1111
timestamp 1670771148
transform 1 0 103316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1117
timestamp 1670771148
transform 1 0 103868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1123
timestamp 1670771148
transform 1 0 104420 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1670771148
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1670771148
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1670771148
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1149
timestamp 1670771148
transform 1 0 106812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1153
timestamp 1670771148
transform 1 0 107180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1159
timestamp 1670771148
transform 1 0 107732 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1165
timestamp 1670771148
transform 1 0 108284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1182
timestamp 1670771148
transform 1 0 109848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1188
timestamp 1670771148
transform 1 0 110400 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1194
timestamp 1670771148
transform 1 0 110952 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1200
timestamp 1670771148
transform 1 0 111504 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1205
timestamp 1670771148
transform 1 0 111964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1209
timestamp 1670771148
transform 1 0 112332 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1212
timestamp 1670771148
transform 1 0 112608 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1218
timestamp 1670771148
transform 1 0 113160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1222
timestamp 1670771148
transform 1 0 113528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1225
timestamp 1670771148
transform 1 0 113804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1234
timestamp 1670771148
transform 1 0 114632 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1242
timestamp 1670771148
transform 1 0 115368 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1246
timestamp 1670771148
transform 1 0 115736 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1255
timestamp 1670771148
transform 1 0 116564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1670771148
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1261
timestamp 1670771148
transform 1 0 117116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1279
timestamp 1670771148
transform 1 0 118772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1287
timestamp 1670771148
transform 1 0 119508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1293
timestamp 1670771148
transform 1 0 120060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1297
timestamp 1670771148
transform 1 0 120428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1300
timestamp 1670771148
transform 1 0 120704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1309
timestamp 1670771148
transform 1 0 121532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1315
timestamp 1670771148
transform 1 0 122084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1317
timestamp 1670771148
transform 1 0 122268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1322
timestamp 1670771148
transform 1 0 122728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1328
timestamp 1670771148
transform 1 0 123280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1336
timestamp 1670771148
transform 1 0 124016 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1342
timestamp 1670771148
transform 1 0 124568 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1364
timestamp 1670771148
transform 1 0 126592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1370
timestamp 1670771148
transform 1 0 127144 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1373
timestamp 1670771148
transform 1 0 127420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1377
timestamp 1670771148
transform 1 0 127788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1381
timestamp 1670771148
transform 1 0 128156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1384
timestamp 1670771148
transform 1 0 128432 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1402
timestamp 1670771148
transform 1 0 130088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1416
timestamp 1670771148
transform 1 0 131376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1426
timestamp 1670771148
transform 1 0 132296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1429
timestamp 1670771148
transform 1 0 132572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1435
timestamp 1670771148
transform 1 0 133124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1441
timestamp 1670771148
transform 1 0 133676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1462
timestamp 1670771148
transform 1 0 135608 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1482
timestamp 1670771148
transform 1 0 137448 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1485
timestamp 1670771148
transform 1 0 137724 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1492
timestamp 1670771148
transform 1 0 138368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1498
timestamp 1670771148
transform 1 0 138920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1504
timestamp 1670771148
transform 1 0 139472 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1510
timestamp 1670771148
transform 1 0 140024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1517
timestamp 1670771148
transform 1 0 140668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1538
timestamp 1670771148
transform 1 0 142600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1541
timestamp 1670771148
transform 1 0 142876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1545
timestamp 1670771148
transform 1 0 143244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1562
timestamp 1670771148
transform 1 0 144808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1582
timestamp 1670771148
transform 1 0 146648 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1588
timestamp 1670771148
transform 1 0 147200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1594
timestamp 1670771148
transform 1 0 147752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1597
timestamp 1670771148
transform 1 0 148028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1615
timestamp 1670771148
transform 1 0 149684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1635
timestamp 1670771148
transform 1 0 151524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1644
timestamp 1670771148
transform 1 0 152352 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1650
timestamp 1670771148
transform 1 0 152904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1653
timestamp 1670771148
transform 1 0 153180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1676
timestamp 1670771148
transform 1 0 155296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1685
timestamp 1670771148
transform 1 0 156124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1694
timestamp 1670771148
transform 1 0 156952 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1701
timestamp 1670771148
transform 1 0 157596 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1707
timestamp 1670771148
transform 1 0 158148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1709
timestamp 1670771148
transform 1 0 158332 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1670771148
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1670771148
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1670771148
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_45
timestamp 1670771148
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1670771148
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1670771148
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1670771148
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_69
timestamp 1670771148
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_79
timestamp 1670771148
transform 1 0 8372 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1670771148
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1670771148
transform 1 0 10120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1670771148
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1670771148
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1670771148
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1670771148
transform 1 0 13248 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_140
timestamp 1670771148
transform 1 0 13984 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1670771148
transform 1 0 14536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1670771148
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1670771148
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_161
timestamp 1670771148
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1670771148
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1670771148
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_173
timestamp 1670771148
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1670771148
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_199
timestamp 1670771148
transform 1 0 19412 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1670771148
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1670771148
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1670771148
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1670771148
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_229
timestamp 1670771148
transform 1 0 22172 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_239
timestamp 1670771148
transform 1 0 23092 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1670771148
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_248
timestamp 1670771148
transform 1 0 23920 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_256
timestamp 1670771148
transform 1 0 24656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1670771148
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1670771148
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_272
timestamp 1670771148
transform 1 0 26128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1670771148
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1670771148
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1670771148
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_306
timestamp 1670771148
transform 1 0 29256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1670771148
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_337
timestamp 1670771148
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_342
timestamp 1670771148
transform 1 0 32568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_350
timestamp 1670771148
transform 1 0 33304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_359
timestamp 1670771148
transform 1 0 34132 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_367
timestamp 1670771148
transform 1 0 34868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_370
timestamp 1670771148
transform 1 0 35144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1670771148
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1670771148
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_397
timestamp 1670771148
transform 1 0 37628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_409
timestamp 1670771148
transform 1 0 38732 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_412
timestamp 1670771148
transform 1 0 39008 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_418
timestamp 1670771148
transform 1 0 39560 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_424
timestamp 1670771148
transform 1 0 40112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_431
timestamp 1670771148
transform 1 0 40756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_438
timestamp 1670771148
transform 1 0 41400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1670771148
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1670771148
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_467
timestamp 1670771148
transform 1 0 44068 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_473
timestamp 1670771148
transform 1 0 44620 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_481
timestamp 1670771148
transform 1 0 45356 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_485
timestamp 1670771148
transform 1 0 45724 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_502
timestamp 1670771148
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_505
timestamp 1670771148
transform 1 0 47564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_510
timestamp 1670771148
transform 1 0 48024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_530
timestamp 1670771148
transform 1 0 49864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_537
timestamp 1670771148
transform 1 0 50508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_545
timestamp 1670771148
transform 1 0 51244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_554
timestamp 1670771148
transform 1 0 52072 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_561
timestamp 1670771148
transform 1 0 52716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_573
timestamp 1670771148
transform 1 0 53820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_577
timestamp 1670771148
transform 1 0 54188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_594
timestamp 1670771148
transform 1 0 55752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_614
timestamp 1670771148
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_617
timestamp 1670771148
transform 1 0 57868 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_628
timestamp 1670771148
transform 1 0 58880 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_648
timestamp 1670771148
transform 1 0 60720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_668
timestamp 1670771148
transform 1 0 62560 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_673
timestamp 1670771148
transform 1 0 63020 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_679
timestamp 1670771148
transform 1 0 63572 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_685
timestamp 1670771148
transform 1 0 64124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_692
timestamp 1670771148
transform 1 0 64768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_698
timestamp 1670771148
transform 1 0 65320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_702
timestamp 1670771148
transform 1 0 65688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_719
timestamp 1670771148
transform 1 0 67252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_723
timestamp 1670771148
transform 1 0 67620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_726
timestamp 1670771148
transform 1 0 67896 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1670771148
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_735
timestamp 1670771148
transform 1 0 68724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_741
timestamp 1670771148
transform 1 0 69276 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_761
timestamp 1670771148
transform 1 0 71116 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_767
timestamp 1670771148
transform 1 0 71668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_770
timestamp 1670771148
transform 1 0 71944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_779
timestamp 1670771148
transform 1 0 72772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1670771148
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_785
timestamp 1670771148
transform 1 0 73324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_792
timestamp 1670771148
transform 1 0 73968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_800
timestamp 1670771148
transform 1 0 74704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_817
timestamp 1670771148
transform 1 0 76268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_821
timestamp 1670771148
transform 1 0 76636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_838
timestamp 1670771148
transform 1 0 78200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_841
timestamp 1670771148
transform 1 0 78476 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_847
timestamp 1670771148
transform 1 0 79028 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_850
timestamp 1670771148
transform 1 0 79304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_870
timestamp 1670771148
transform 1 0 81144 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_881
timestamp 1670771148
transform 1 0 82156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_890
timestamp 1670771148
transform 1 0 82984 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1670771148
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_909
timestamp 1670771148
transform 1 0 84732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_913
timestamp 1670771148
transform 1 0 85100 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_931
timestamp 1670771148
transform 1 0 86756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_937
timestamp 1670771148
transform 1 0 87308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_943
timestamp 1670771148
transform 1 0 87860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_947
timestamp 1670771148
transform 1 0 88228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_950
timestamp 1670771148
transform 1 0 88504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_953
timestamp 1670771148
transform 1 0 88780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_959
timestamp 1670771148
transform 1 0 89332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_965
timestamp 1670771148
transform 1 0 89884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_989
timestamp 1670771148
transform 1 0 92092 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_997
timestamp 1670771148
transform 1 0 92828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1003
timestamp 1670771148
transform 1 0 93380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1670771148
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1009
timestamp 1670771148
transform 1 0 93932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1015
timestamp 1670771148
transform 1 0 94484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1021
timestamp 1670771148
transform 1 0 95036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1027
timestamp 1670771148
transform 1 0 95588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1033
timestamp 1670771148
transform 1 0 96140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1037
timestamp 1670771148
transform 1 0 96508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1040
timestamp 1670771148
transform 1 0 96784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1052
timestamp 1670771148
transform 1 0 97888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1058
timestamp 1670771148
transform 1 0 98440 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1670771148
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1077
timestamp 1670771148
transform 1 0 100188 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1083
timestamp 1670771148
transform 1 0 100740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1100
timestamp 1670771148
transform 1 0 102304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1106
timestamp 1670771148
transform 1 0 102856 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1110
timestamp 1670771148
transform 1 0 103224 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1115
timestamp 1670771148
transform 1 0 103684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1119
timestamp 1670771148
transform 1 0 104052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1121
timestamp 1670771148
transform 1 0 104236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1125
timestamp 1670771148
transform 1 0 104604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1129
timestamp 1670771148
transform 1 0 104972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1146
timestamp 1670771148
transform 1 0 106536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1152
timestamp 1670771148
transform 1 0 107088 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1158
timestamp 1670771148
transform 1 0 107640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1164
timestamp 1670771148
transform 1 0 108192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1170
timestamp 1670771148
transform 1 0 108744 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1177
timestamp 1670771148
transform 1 0 109388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1181
timestamp 1670771148
transform 1 0 109756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1187
timestamp 1670771148
transform 1 0 110308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1193
timestamp 1670771148
transform 1 0 110860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1202
timestamp 1670771148
transform 1 0 111688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1208
timestamp 1670771148
transform 1 0 112240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1214
timestamp 1670771148
transform 1 0 112792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1222
timestamp 1670771148
transform 1 0 113528 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1226
timestamp 1670771148
transform 1 0 113896 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1233
timestamp 1670771148
transform 1 0 114540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1237
timestamp 1670771148
transform 1 0 114908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1243
timestamp 1670771148
transform 1 0 115460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1264
timestamp 1670771148
transform 1 0 117392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1284
timestamp 1670771148
transform 1 0 119232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1289
timestamp 1670771148
transform 1 0 119692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1299
timestamp 1670771148
transform 1 0 120612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1319
timestamp 1670771148
transform 1 0 122452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1327
timestamp 1670771148
transform 1 0 123188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1333
timestamp 1670771148
transform 1 0 123740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1339
timestamp 1670771148
transform 1 0 124292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1343
timestamp 1670771148
transform 1 0 124660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1345
timestamp 1670771148
transform 1 0 124844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1349
timestamp 1670771148
transform 1 0 125212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1352
timestamp 1670771148
transform 1 0 125488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1361
timestamp 1670771148
transform 1 0 126316 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1368
timestamp 1670771148
transform 1 0 126960 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1376
timestamp 1670771148
transform 1 0 127696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1381
timestamp 1670771148
transform 1 0 128156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1395
timestamp 1670771148
transform 1 0 129444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1399
timestamp 1670771148
transform 1 0 129812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1401
timestamp 1670771148
transform 1 0 129996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1405
timestamp 1670771148
transform 1 0 130364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1411
timestamp 1670771148
transform 1 0 130916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1431
timestamp 1670771148
transform 1 0 132756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1437
timestamp 1670771148
transform 1 0 133308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1443
timestamp 1670771148
transform 1 0 133860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1451
timestamp 1670771148
transform 1 0 134596 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1454
timestamp 1670771148
transform 1 0 134872 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1457
timestamp 1670771148
transform 1 0 135148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1463
timestamp 1670771148
transform 1 0 135700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1469
timestamp 1670771148
transform 1 0 136252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1475
timestamp 1670771148
transform 1 0 136804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1496
timestamp 1670771148
transform 1 0 138736 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1502
timestamp 1670771148
transform 1 0 139288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1508
timestamp 1670771148
transform 1 0 139840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1513
timestamp 1670771148
transform 1 0 140300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1519
timestamp 1670771148
transform 1 0 140852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1523
timestamp 1670771148
transform 1 0 141220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1549
timestamp 1670771148
transform 1 0 143612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1558
timestamp 1670771148
transform 1 0 144440 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1564
timestamp 1670771148
transform 1 0 144992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1569
timestamp 1670771148
transform 1 0 145452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1587
timestamp 1670771148
transform 1 0 147108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1607
timestamp 1670771148
transform 1 0 148948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1615
timestamp 1670771148
transform 1 0 149684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1622
timestamp 1670771148
transform 1 0 150328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1625
timestamp 1670771148
transform 1 0 150604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1643
timestamp 1670771148
transform 1 0 152260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1663
timestamp 1670771148
transform 1 0 154100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1672
timestamp 1670771148
transform 1 0 154928 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1678
timestamp 1670771148
transform 1 0 155480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1681
timestamp 1670771148
transform 1 0 155756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1688
timestamp 1670771148
transform 1 0 156400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1697
timestamp 1670771148
transform 1 0 157228 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1704
timestamp 1670771148
transform 1 0 157872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1710
timestamp 1670771148
transform 1 0 158424 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1670771148
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1670771148
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1670771148
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1670771148
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 1670771148
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1670771148
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1670771148
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1670771148
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1670771148
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1670771148
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1670771148
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1670771148
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_89
timestamp 1670771148
transform 1 0 9292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1670771148
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1670771148
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1670771148
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1670771148
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1670771148
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1670771148
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1670771148
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1670771148
transform 1 0 17664 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1670771148
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1670771148
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1670771148
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1670771148
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_239
timestamp 1670771148
transform 1 0 23092 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_247
timestamp 1670771148
transform 1 0 23828 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1670771148
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1670771148
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1670771148
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_264
timestamp 1670771148
transform 1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_270
timestamp 1670771148
transform 1 0 25944 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_273
timestamp 1670771148
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_282
timestamp 1670771148
transform 1 0 27048 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_290
timestamp 1670771148
transform 1 0 27784 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_300
timestamp 1670771148
transform 1 0 28704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1670771148
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1670771148
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_327
timestamp 1670771148
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_331
timestamp 1670771148
transform 1 0 31556 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_348
timestamp 1670771148
transform 1 0 33120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_355
timestamp 1670771148
transform 1 0 33764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1670771148
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1670771148
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1670771148
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_392
timestamp 1670771148
transform 1 0 37168 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_396
timestamp 1670771148
transform 1 0 37536 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1670771148
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_405
timestamp 1670771148
transform 1 0 38364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_411
timestamp 1670771148
transform 1 0 38916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1670771148
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1670771148
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_425
timestamp 1670771148
transform 1 0 40204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_433
timestamp 1670771148
transform 1 0 40940 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_441
timestamp 1670771148
transform 1 0 41676 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_446
timestamp 1670771148
transform 1 0 42136 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_454
timestamp 1670771148
transform 1 0 42872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1670771148
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_477
timestamp 1670771148
transform 1 0 44988 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_486
timestamp 1670771148
transform 1 0 45816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_506
timestamp 1670771148
transform 1 0 47656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_518
timestamp 1670771148
transform 1 0 48760 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_524
timestamp 1670771148
transform 1 0 49312 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_530
timestamp 1670771148
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_533
timestamp 1670771148
transform 1 0 50140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_539
timestamp 1670771148
transform 1 0 50692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_545
timestamp 1670771148
transform 1 0 51244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_549
timestamp 1670771148
transform 1 0 51612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_566
timestamp 1670771148
transform 1 0 53176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_586
timestamp 1670771148
transform 1 0 55016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_589
timestamp 1670771148
transform 1 0 55292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_607
timestamp 1670771148
transform 1 0 56948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_619
timestamp 1670771148
transform 1 0 58052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_628
timestamp 1670771148
transform 1 0 58880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_634
timestamp 1670771148
transform 1 0 59432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_642
timestamp 1670771148
transform 1 0 60168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_645
timestamp 1670771148
transform 1 0 60444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_663
timestamp 1670771148
transform 1 0 62100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_671
timestamp 1670771148
transform 1 0 62836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_675
timestamp 1670771148
transform 1 0 63204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_678
timestamp 1670771148
transform 1 0 63480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_698
timestamp 1670771148
transform 1 0 65320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_701
timestamp 1670771148
transform 1 0 65596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_705
timestamp 1670771148
transform 1 0 65964 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_711
timestamp 1670771148
transform 1 0 66516 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_715
timestamp 1670771148
transform 1 0 66884 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_721
timestamp 1670771148
transform 1 0 67436 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_742
timestamp 1670771148
transform 1 0 69368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_751
timestamp 1670771148
transform 1 0 70196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1670771148
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_757
timestamp 1670771148
transform 1 0 70748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_765
timestamp 1670771148
transform 1 0 71484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_785
timestamp 1670771148
transform 1 0 73324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_791
timestamp 1670771148
transform 1 0 73876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_794
timestamp 1670771148
transform 1 0 74152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_798
timestamp 1670771148
transform 1 0 74520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_801
timestamp 1670771148
transform 1 0 74796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_805
timestamp 1670771148
transform 1 0 75164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_809
timestamp 1670771148
transform 1 0 75532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_813
timestamp 1670771148
transform 1 0 75900 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_819
timestamp 1670771148
transform 1 0 76452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_836
timestamp 1670771148
transform 1 0 78016 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_846
timestamp 1670771148
transform 1 0 78936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_866
timestamp 1670771148
transform 1 0 80776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_869
timestamp 1670771148
transform 1 0 81052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_873
timestamp 1670771148
transform 1 0 81420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_877
timestamp 1670771148
transform 1 0 81788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_880
timestamp 1670771148
transform 1 0 82064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_900
timestamp 1670771148
transform 1 0 83904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_912
timestamp 1670771148
transform 1 0 85008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_922
timestamp 1670771148
transform 1 0 85928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_925
timestamp 1670771148
transform 1 0 86204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_929
timestamp 1670771148
transform 1 0 86572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_951
timestamp 1670771148
transform 1 0 88596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_971
timestamp 1670771148
transform 1 0 90436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_977
timestamp 1670771148
transform 1 0 90988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_981
timestamp 1670771148
transform 1 0 91356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_985
timestamp 1670771148
transform 1 0 91724 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_991
timestamp 1670771148
transform 1 0 92276 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1009
timestamp 1670771148
transform 1 0 93932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1015
timestamp 1670771148
transform 1 0 94484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1021
timestamp 1670771148
transform 1 0 95036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1027
timestamp 1670771148
transform 1 0 95588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1033
timestamp 1670771148
transform 1 0 96140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1037
timestamp 1670771148
transform 1 0 96508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1056
timestamp 1670771148
transform 1 0 98256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1063
timestamp 1670771148
transform 1 0 98900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1069
timestamp 1670771148
transform 1 0 99452 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1075
timestamp 1670771148
transform 1 0 100004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1087
timestamp 1670771148
transform 1 0 101108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1670771148
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1093
timestamp 1670771148
transform 1 0 101660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1112
timestamp 1670771148
transform 1 0 103408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1132
timestamp 1670771148
transform 1 0 105248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1138
timestamp 1670771148
transform 1 0 105800 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1144
timestamp 1670771148
transform 1 0 106352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1149
timestamp 1670771148
transform 1 0 106812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1153
timestamp 1670771148
transform 1 0 107180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1159
timestamp 1670771148
transform 1 0 107732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1163
timestamp 1670771148
transform 1 0 108100 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1166
timestamp 1670771148
transform 1 0 108376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1175
timestamp 1670771148
transform 1 0 109204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1195
timestamp 1670771148
transform 1 0 111044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1202
timestamp 1670771148
transform 1 0 111688 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1205
timestamp 1670771148
transform 1 0 111964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1209
timestamp 1670771148
transform 1 0 112332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1215
timestamp 1670771148
transform 1 0 112884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1221
timestamp 1670771148
transform 1 0 113436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1241
timestamp 1670771148
transform 1 0 115276 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1247
timestamp 1670771148
transform 1 0 115828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1253
timestamp 1670771148
transform 1 0 116380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1259
timestamp 1670771148
transform 1 0 116932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1261
timestamp 1670771148
transform 1 0 117116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1266
timestamp 1670771148
transform 1 0 117576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1284
timestamp 1670771148
transform 1 0 119232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1290
timestamp 1670771148
transform 1 0 119784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1296
timestamp 1670771148
transform 1 0 120336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1305
timestamp 1670771148
transform 1 0 121164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1313
timestamp 1670771148
transform 1 0 121900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1317
timestamp 1670771148
transform 1 0 122268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1321
timestamp 1670771148
transform 1 0 122636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1327
timestamp 1670771148
transform 1 0 123188 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1335
timestamp 1670771148
transform 1 0 123924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1352
timestamp 1670771148
transform 1 0 125488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1356
timestamp 1670771148
transform 1 0 125856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1362
timestamp 1670771148
transform 1 0 126408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1368
timestamp 1670771148
transform 1 0 126960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1373
timestamp 1670771148
transform 1 0 127420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1387
timestamp 1670771148
transform 1 0 128708 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1407
timestamp 1670771148
transform 1 0 130548 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1417
timestamp 1670771148
transform 1 0 131468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1426
timestamp 1670771148
transform 1 0 132296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1429
timestamp 1670771148
transform 1 0 132572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1451
timestamp 1670771148
transform 1 0 134596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1457
timestamp 1670771148
transform 1 0 135148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1463
timestamp 1670771148
transform 1 0 135700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1469
timestamp 1670771148
transform 1 0 136252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1473
timestamp 1670771148
transform 1 0 136620 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1476
timestamp 1670771148
transform 1 0 136896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1482
timestamp 1670771148
transform 1 0 137448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1485
timestamp 1670771148
transform 1 0 137724 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1491
timestamp 1670771148
transform 1 0 138276 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1494
timestamp 1670771148
transform 1 0 138552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1502
timestamp 1670771148
transform 1 0 139288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1509
timestamp 1670771148
transform 1 0 139932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1515
timestamp 1670771148
transform 1 0 140484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1526
timestamp 1670771148
transform 1 0 141496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1530
timestamp 1670771148
transform 1 0 141864 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1536
timestamp 1670771148
transform 1 0 142416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1541
timestamp 1670771148
transform 1 0 142876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1545
timestamp 1670771148
transform 1 0 143244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1563
timestamp 1670771148
transform 1 0 144900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1583
timestamp 1670771148
transform 1 0 146740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1591
timestamp 1670771148
transform 1 0 147476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1595
timestamp 1670771148
transform 1 0 147844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1597
timestamp 1670771148
transform 1 0 148028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1604
timestamp 1670771148
transform 1 0 148672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1608
timestamp 1670771148
transform 1 0 149040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1626
timestamp 1670771148
transform 1 0 150696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1646
timestamp 1670771148
transform 1 0 152536 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1653
timestamp 1670771148
transform 1 0 153180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1671
timestamp 1670771148
transform 1 0 154836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1680
timestamp 1670771148
transform 1 0 155664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1689
timestamp 1670771148
transform 1 0 156492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1696
timestamp 1670771148
transform 1 0 157136 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1703
timestamp 1670771148
transform 1 0 157780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1707
timestamp 1670771148
transform 1 0 158148 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1709
timestamp 1670771148
transform 1 0 158332 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1670771148
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1670771148
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1670771148
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1670771148
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1670771148
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1670771148
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1670771148
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1670771148
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1670771148
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_82
timestamp 1670771148
transform 1 0 8648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1670771148
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1670771148
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_97
timestamp 1670771148
transform 1 0 10028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1670771148
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1670771148
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1670771148
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 1670771148
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1670771148
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1670771148
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1670771148
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1670771148
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1670771148
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1670771148
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_190
timestamp 1670771148
transform 1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_194
timestamp 1670771148
transform 1 0 18952 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1670771148
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1670771148
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1670771148
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1670771148
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1670771148
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1670771148
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_231
timestamp 1670771148
transform 1 0 22356 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_240
timestamp 1670771148
transform 1 0 23184 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1670771148
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_257
timestamp 1670771148
transform 1 0 24748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1670771148
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 1670771148
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1670771148
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1670771148
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_326
timestamp 1670771148
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1670771148
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1670771148
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_341
timestamp 1670771148
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_347
timestamp 1670771148
transform 1 0 33028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_351
timestamp 1670771148
transform 1 0 33396 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_354
timestamp 1670771148
transform 1 0 33672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_358
timestamp 1670771148
transform 1 0 34040 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_361
timestamp 1670771148
transform 1 0 34316 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_367
timestamp 1670771148
transform 1 0 34868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_379
timestamp 1670771148
transform 1 0 35972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_384
timestamp 1670771148
transform 1 0 36432 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1670771148
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1670771148
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_397
timestamp 1670771148
transform 1 0 37628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_400
timestamp 1670771148
transform 1 0 37904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_420
timestamp 1670771148
transform 1 0 39744 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_433
timestamp 1670771148
transform 1 0 40940 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_441
timestamp 1670771148
transform 1 0 41676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1670771148
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_449
timestamp 1670771148
transform 1 0 42412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_456
timestamp 1670771148
transform 1 0 43056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_464
timestamp 1670771148
transform 1 0 43792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_472
timestamp 1670771148
transform 1 0 44528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_480
timestamp 1670771148
transform 1 0 45264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1670771148
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_505
timestamp 1670771148
transform 1 0 47564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_509
timestamp 1670771148
transform 1 0 47932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_517
timestamp 1670771148
transform 1 0 48668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_525
timestamp 1670771148
transform 1 0 49404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_545
timestamp 1670771148
transform 1 0 51244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_549
timestamp 1670771148
transform 1 0 51612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_555
timestamp 1670771148
transform 1 0 52164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1670771148
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_561
timestamp 1670771148
transform 1 0 52716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_566
timestamp 1670771148
transform 1 0 53176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_574
timestamp 1670771148
transform 1 0 53912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_594
timestamp 1670771148
transform 1 0 55752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1670771148
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_617
timestamp 1670771148
transform 1 0 57868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_635
timestamp 1670771148
transform 1 0 59524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_641
timestamp 1670771148
transform 1 0 60076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_650
timestamp 1670771148
transform 1 0 60904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_670
timestamp 1670771148
transform 1 0 62744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_673
timestamp 1670771148
transform 1 0 63020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_679
timestamp 1670771148
transform 1 0 63572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_687
timestamp 1670771148
transform 1 0 64308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_697
timestamp 1670771148
transform 1 0 65228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_717
timestamp 1670771148
transform 1 0 67068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_726
timestamp 1670771148
transform 1 0 67896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_729
timestamp 1670771148
transform 1 0 68172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_736
timestamp 1670771148
transform 1 0 68816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_756
timestamp 1670771148
transform 1 0 70656 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_762
timestamp 1670771148
transform 1 0 71208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_776
timestamp 1670771148
transform 1 0 72496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_782
timestamp 1670771148
transform 1 0 73048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_785
timestamp 1670771148
transform 1 0 73324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_789
timestamp 1670771148
transform 1 0 73692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_792
timestamp 1670771148
transform 1 0 73968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_798
timestamp 1670771148
transform 1 0 74520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_806
timestamp 1670771148
transform 1 0 75256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_814
timestamp 1670771148
transform 1 0 75992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_831
timestamp 1670771148
transform 1 0 77556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_835
timestamp 1670771148
transform 1 0 77924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_838
timestamp 1670771148
transform 1 0 78200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_841
timestamp 1670771148
transform 1 0 78476 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_847
timestamp 1670771148
transform 1 0 79028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_864
timestamp 1670771148
transform 1 0 80592 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_870
timestamp 1670771148
transform 1 0 81144 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_882
timestamp 1670771148
transform 1 0 82248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_891
timestamp 1670771148
transform 1 0 83076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1670771148
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_897
timestamp 1670771148
transform 1 0 83628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_904
timestamp 1670771148
transform 1 0 84272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_912
timestamp 1670771148
transform 1 0 85008 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_932
timestamp 1670771148
transform 1 0 86848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_940
timestamp 1670771148
transform 1 0 87584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_946
timestamp 1670771148
transform 1 0 88136 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_953
timestamp 1670771148
transform 1 0 88780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_971
timestamp 1670771148
transform 1 0 90436 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_995
timestamp 1670771148
transform 1 0 92644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1670771148
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1670771148
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1009
timestamp 1670771148
transform 1 0 93932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1015
timestamp 1670771148
transform 1 0 94484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1023
timestamp 1670771148
transform 1 0 95220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1029
timestamp 1670771148
transform 1 0 95772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1035
timestamp 1670771148
transform 1 0 96324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1041
timestamp 1670771148
transform 1 0 96876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1047
timestamp 1670771148
transform 1 0 97428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1053
timestamp 1670771148
transform 1 0 97980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1059
timestamp 1670771148
transform 1 0 98532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1670771148
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1065
timestamp 1670771148
transform 1 0 99084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1069
timestamp 1670771148
transform 1 0 99452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1075
timestamp 1670771148
transform 1 0 100004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1098
timestamp 1670771148
transform 1 0 102120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1104
timestamp 1670771148
transform 1 0 102672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1114
timestamp 1670771148
transform 1 0 103592 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1121
timestamp 1670771148
transform 1 0 104236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1140
timestamp 1670771148
transform 1 0 105984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1146
timestamp 1670771148
transform 1 0 106536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1152
timestamp 1670771148
transform 1 0 107088 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1160
timestamp 1670771148
transform 1 0 107824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1164
timestamp 1670771148
transform 1 0 108192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1170
timestamp 1670771148
transform 1 0 108744 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1177
timestamp 1670771148
transform 1 0 109388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1181
timestamp 1670771148
transform 1 0 109756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1187
timestamp 1670771148
transform 1 0 110308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1191
timestamp 1670771148
transform 1 0 110676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1212
timestamp 1670771148
transform 1 0 112608 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1218
timestamp 1670771148
transform 1 0 113160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1222
timestamp 1670771148
transform 1 0 113528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1228
timestamp 1670771148
transform 1 0 114080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1233
timestamp 1670771148
transform 1 0 114540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1237
timestamp 1670771148
transform 1 0 114908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1248
timestamp 1670771148
transform 1 0 115920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1268
timestamp 1670771148
transform 1 0 117760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1277
timestamp 1670771148
transform 1 0 118588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1283
timestamp 1670771148
transform 1 0 119140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1287
timestamp 1670771148
transform 1 0 119508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1289
timestamp 1670771148
transform 1 0 119692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1293
timestamp 1670771148
transform 1 0 120060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1299
timestamp 1670771148
transform 1 0 120612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1308
timestamp 1670771148
transform 1 0 121440 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1316
timestamp 1670771148
transform 1 0 122176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1322
timestamp 1670771148
transform 1 0 122728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1328
timestamp 1670771148
transform 1 0 123280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1334
timestamp 1670771148
transform 1 0 123832 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1340
timestamp 1670771148
transform 1 0 124384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1345
timestamp 1670771148
transform 1 0 124844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1349
timestamp 1670771148
transform 1 0 125212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1355
timestamp 1670771148
transform 1 0 125764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1364
timestamp 1670771148
transform 1 0 126592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1373
timestamp 1670771148
transform 1 0 127420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1380
timestamp 1670771148
transform 1 0 128064 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1389
timestamp 1670771148
transform 1 0 128892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1395
timestamp 1670771148
transform 1 0 129444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1399
timestamp 1670771148
transform 1 0 129812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1401
timestamp 1670771148
transform 1 0 129996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1405
timestamp 1670771148
transform 1 0 130364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1411
timestamp 1670771148
transform 1 0 130916 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1417
timestamp 1670771148
transform 1 0 131468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1423
timestamp 1670771148
transform 1 0 132020 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1429
timestamp 1670771148
transform 1 0 132572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1433
timestamp 1670771148
transform 1 0 132940 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1450
timestamp 1670771148
transform 1 0 134504 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1457
timestamp 1670771148
transform 1 0 135148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1475
timestamp 1670771148
transform 1 0 136804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1481
timestamp 1670771148
transform 1 0 137356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1487
timestamp 1670771148
transform 1 0 137908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1490
timestamp 1670771148
transform 1 0 138184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1510
timestamp 1670771148
transform 1 0 140024 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1513
timestamp 1670771148
transform 1 0 140300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1520
timestamp 1670771148
transform 1 0 140944 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1542
timestamp 1670771148
transform 1 0 142968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1562
timestamp 1670771148
transform 1 0 144808 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1569
timestamp 1670771148
transform 1 0 145452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1587
timestamp 1670771148
transform 1 0 147108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1607
timestamp 1670771148
transform 1 0 148948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1615
timestamp 1670771148
transform 1 0 149684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1622
timestamp 1670771148
transform 1 0 150328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1625
timestamp 1670771148
transform 1 0 150604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1643
timestamp 1670771148
transform 1 0 152260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1663
timestamp 1670771148
transform 1 0 154100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1672
timestamp 1670771148
transform 1 0 154928 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1678
timestamp 1670771148
transform 1 0 155480 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1681
timestamp 1670771148
transform 1 0 155756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1688
timestamp 1670771148
transform 1 0 156400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1697
timestamp 1670771148
transform 1 0 157228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1704
timestamp 1670771148
transform 1 0 157872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1710
timestamp 1670771148
transform 1 0 158424 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1670771148
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1670771148
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1670771148
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1670771148
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_35
timestamp 1670771148
transform 1 0 4324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_39
timestamp 1670771148
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_51
timestamp 1670771148
transform 1 0 5796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_73
timestamp 1670771148
transform 1 0 7820 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1670771148
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1670771148
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1670771148
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1670771148
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1670771148
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_104
timestamp 1670771148
transform 1 0 10672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1670771148
transform 1 0 12512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1670771148
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1670771148
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1670771148
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_145
timestamp 1670771148
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1670771148
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_173
timestamp 1670771148
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1670771148
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1670771148
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_203
timestamp 1670771148
transform 1 0 19780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1670771148
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_229
timestamp 1670771148
transform 1 0 22172 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1670771148
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_245
timestamp 1670771148
transform 1 0 23644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1670771148
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1670771148
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1670771148
transform 1 0 26036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1670771148
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_287
timestamp 1670771148
transform 1 0 27508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_295
timestamp 1670771148
transform 1 0 28244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_303
timestamp 1670771148
transform 1 0 28980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1670771148
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1670771148
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_315
timestamp 1670771148
transform 1 0 30084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1670771148
transform 1 0 32108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_345
timestamp 1670771148
transform 1 0 32844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1670771148
transform 1 0 33580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1670771148
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_365
timestamp 1670771148
transform 1 0 34684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_373
timestamp 1670771148
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_385
timestamp 1670771148
transform 1 0 36524 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_397
timestamp 1670771148
transform 1 0 37628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1670771148
transform 1 0 38732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_413
timestamp 1670771148
transform 1 0 39100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1670771148
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1670771148
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_441
timestamp 1670771148
transform 1 0 41676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_448
timestamp 1670771148
transform 1 0 42320 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_457
timestamp 1670771148
transform 1 0 43148 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_461
timestamp 1670771148
transform 1 0 43516 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_466
timestamp 1670771148
transform 1 0 43976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1670771148
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_477
timestamp 1670771148
transform 1 0 44988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_483
timestamp 1670771148
transform 1 0 45540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_503
timestamp 1670771148
transform 1 0 47380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_523
timestamp 1670771148
transform 1 0 49220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_527
timestamp 1670771148
transform 1 0 49588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_530
timestamp 1670771148
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_533
timestamp 1670771148
transform 1 0 50140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_537
timestamp 1670771148
transform 1 0 50508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_542
timestamp 1670771148
transform 1 0 50968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_550
timestamp 1670771148
transform 1 0 51704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_570
timestamp 1670771148
transform 1 0 53544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_578
timestamp 1670771148
transform 1 0 54280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_586
timestamp 1670771148
transform 1 0 55016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_589
timestamp 1670771148
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_596
timestamp 1670771148
transform 1 0 55936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_600
timestamp 1670771148
transform 1 0 56304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_606
timestamp 1670771148
transform 1 0 56856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_626
timestamp 1670771148
transform 1 0 58696 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1670771148
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1670771148
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_645
timestamp 1670771148
transform 1 0 60444 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_667
timestamp 1670771148
transform 1 0 62468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_677
timestamp 1670771148
transform 1 0 63388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_685
timestamp 1670771148
transform 1 0 64124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_697
timestamp 1670771148
transform 1 0 65228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_701
timestamp 1670771148
transform 1 0 65596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_707
timestamp 1670771148
transform 1 0 66148 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_713
timestamp 1670771148
transform 1 0 66700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_719
timestamp 1670771148
transform 1 0 67252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_725
timestamp 1670771148
transform 1 0 67804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_731
timestamp 1670771148
transform 1 0 68356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_739
timestamp 1670771148
transform 1 0 69092 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_751
timestamp 1670771148
transform 1 0 70196 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1670771148
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_757
timestamp 1670771148
transform 1 0 70748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_761
timestamp 1670771148
transform 1 0 71116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_765
timestamp 1670771148
transform 1 0 71484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_768
timestamp 1670771148
transform 1 0 71760 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_776
timestamp 1670771148
transform 1 0 72496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_782
timestamp 1670771148
transform 1 0 73048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_788
timestamp 1670771148
transform 1 0 73600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_808
timestamp 1670771148
transform 1 0 75440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_813
timestamp 1670771148
transform 1 0 75900 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_819
timestamp 1670771148
transform 1 0 76452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_822
timestamp 1670771148
transform 1 0 76728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_826
timestamp 1670771148
transform 1 0 77096 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_829
timestamp 1670771148
transform 1 0 77372 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_849
timestamp 1670771148
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1670771148
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1670771148
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_869
timestamp 1670771148
transform 1 0 81052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_876
timestamp 1670771148
transform 1 0 81696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_882
timestamp 1670771148
transform 1 0 82248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_888
timestamp 1670771148
transform 1 0 82800 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_894
timestamp 1670771148
transform 1 0 83352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_900
timestamp 1670771148
transform 1 0 83904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_906
timestamp 1670771148
transform 1 0 84456 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_914
timestamp 1670771148
transform 1 0 85192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_919
timestamp 1670771148
transform 1 0 85652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1670771148
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_925
timestamp 1670771148
transform 1 0 86204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_931
timestamp 1670771148
transform 1 0 86756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_937
timestamp 1670771148
transform 1 0 87308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_941
timestamp 1670771148
transform 1 0 87676 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_958
timestamp 1670771148
transform 1 0 89240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_966
timestamp 1670771148
transform 1 0 89976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_974
timestamp 1670771148
transform 1 0 90712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_981
timestamp 1670771148
transform 1 0 91356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_999
timestamp 1670771148
transform 1 0 93012 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1007
timestamp 1670771148
transform 1 0 93748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1013
timestamp 1670771148
transform 1 0 94300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1034
timestamp 1670771148
transform 1 0 96232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1037
timestamp 1670771148
transform 1 0 96508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1043
timestamp 1670771148
transform 1 0 97060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1047
timestamp 1670771148
transform 1 0 97428 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1051
timestamp 1670771148
transform 1 0 97796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1057
timestamp 1670771148
transform 1 0 98348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1063
timestamp 1670771148
transform 1 0 98900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1069
timestamp 1670771148
transform 1 0 99452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1075
timestamp 1670771148
transform 1 0 100004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1081
timestamp 1670771148
transform 1 0 100556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1087
timestamp 1670771148
transform 1 0 101108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1090
timestamp 1670771148
transform 1 0 101384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1093
timestamp 1670771148
transform 1 0 101660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1097
timestamp 1670771148
transform 1 0 102028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1108
timestamp 1670771148
transform 1 0 103040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1114
timestamp 1670771148
transform 1 0 103592 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1127
timestamp 1670771148
transform 1 0 104788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1135
timestamp 1670771148
transform 1 0 105524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1143
timestamp 1670771148
transform 1 0 106260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1147
timestamp 1670771148
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1149
timestamp 1670771148
transform 1 0 106812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1155
timestamp 1670771148
transform 1 0 107364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1161
timestamp 1670771148
transform 1 0 107916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1181
timestamp 1670771148
transform 1 0 109756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1189
timestamp 1670771148
transform 1 0 110492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1198
timestamp 1670771148
transform 1 0 111320 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1205
timestamp 1670771148
transform 1 0 111964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1211
timestamp 1670771148
transform 1 0 112516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1217
timestamp 1670771148
transform 1 0 113068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1223
timestamp 1670771148
transform 1 0 113620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1229
timestamp 1670771148
transform 1 0 114172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1235
timestamp 1670771148
transform 1 0 114724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1243
timestamp 1670771148
transform 1 0 115460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1255
timestamp 1670771148
transform 1 0 116564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1670771148
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1261
timestamp 1670771148
transform 1 0 117116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1265
timestamp 1670771148
transform 1 0 117484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1271
timestamp 1670771148
transform 1 0 118036 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1296
timestamp 1670771148
transform 1 0 120336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1302
timestamp 1670771148
transform 1 0 120888 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1314
timestamp 1670771148
transform 1 0 121992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1317
timestamp 1670771148
transform 1 0 122268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1335
timestamp 1670771148
transform 1 0 123924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1343
timestamp 1670771148
transform 1 0 124660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1349
timestamp 1670771148
transform 1 0 125212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1355
timestamp 1670771148
transform 1 0 125764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1361
timestamp 1670771148
transform 1 0 126316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1367
timestamp 1670771148
transform 1 0 126868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1371
timestamp 1670771148
transform 1 0 127236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1373
timestamp 1670771148
transform 1 0 127420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1379
timestamp 1670771148
transform 1 0 127972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1385
timestamp 1670771148
transform 1 0 128524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1391
timestamp 1670771148
transform 1 0 129076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1397
timestamp 1670771148
transform 1 0 129628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1403
timestamp 1670771148
transform 1 0 130180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1409
timestamp 1670771148
transform 1 0 130732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1415
timestamp 1670771148
transform 1 0 131284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1421
timestamp 1670771148
transform 1 0 131836 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1427
timestamp 1670771148
transform 1 0 132388 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1429
timestamp 1670771148
transform 1 0 132572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1433
timestamp 1670771148
transform 1 0 132940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1439
timestamp 1670771148
transform 1 0 133492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1445
timestamp 1670771148
transform 1 0 134044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1462
timestamp 1670771148
transform 1 0 135608 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1473
timestamp 1670771148
transform 1 0 136620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1479
timestamp 1670771148
transform 1 0 137172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1483
timestamp 1670771148
transform 1 0 137540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1485
timestamp 1670771148
transform 1 0 137724 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1489
timestamp 1670771148
transform 1 0 138092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1495
timestamp 1670771148
transform 1 0 138644 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1499
timestamp 1670771148
transform 1 0 139012 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1516
timestamp 1670771148
transform 1 0 140576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1526
timestamp 1670771148
transform 1 0 141496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1534
timestamp 1670771148
transform 1 0 142232 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1541
timestamp 1670771148
transform 1 0 142876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1560
timestamp 1670771148
transform 1 0 144624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1580
timestamp 1670771148
transform 1 0 146464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1588
timestamp 1670771148
transform 1 0 147200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1594
timestamp 1670771148
transform 1 0 147752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1597
timestamp 1670771148
transform 1 0 148028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1603
timestamp 1670771148
transform 1 0 148580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1611
timestamp 1670771148
transform 1 0 149316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1634
timestamp 1670771148
transform 1 0 151432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1641
timestamp 1670771148
transform 1 0 152076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1650
timestamp 1670771148
transform 1 0 152904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1653
timestamp 1670771148
transform 1 0 153180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1671
timestamp 1670771148
transform 1 0 154836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1680
timestamp 1670771148
transform 1 0 155664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1688
timestamp 1670771148
transform 1 0 156400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1696
timestamp 1670771148
transform 1 0 157136 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1703
timestamp 1670771148
transform 1 0 157780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1707
timestamp 1670771148
transform 1 0 158148 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1709
timestamp 1670771148
transform 1 0 158332 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1670771148
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1670771148
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1670771148
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1670771148
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1670771148
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1670771148
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1670771148
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1670771148
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1670771148
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1670771148
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 1670771148
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1670771148
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_94
timestamp 1670771148
transform 1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_102
timestamp 1670771148
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1670771148
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1670771148
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_120
timestamp 1670771148
transform 1 0 12144 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_126
timestamp 1670771148
transform 1 0 12696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1670771148
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1670771148
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_158
timestamp 1670771148
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1670771148
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1670771148
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1670771148
transform 1 0 17020 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1670771148
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1670771148
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1670771148
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1670771148
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1670771148
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1670771148
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_229
timestamp 1670771148
transform 1 0 22172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1670771148
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1670771148
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_265
timestamp 1670771148
transform 1 0 25484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_273
timestamp 1670771148
transform 1 0 26220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1670771148
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1670771148
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_303
timestamp 1670771148
transform 1 0 28980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_309
timestamp 1670771148
transform 1 0 29532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_314
timestamp 1670771148
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1670771148
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1670771148
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_343
timestamp 1670771148
transform 1 0 32660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_355
timestamp 1670771148
transform 1 0 33764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1670771148
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_379
timestamp 1670771148
transform 1 0 35972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_382
timestamp 1670771148
transform 1 0 36248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1670771148
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1670771148
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_397
timestamp 1670771148
transform 1 0 37628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_402
timestamp 1670771148
transform 1 0 38088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_410
timestamp 1670771148
transform 1 0 38824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1670771148
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_426
timestamp 1670771148
transform 1 0 40296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1670771148
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1670771148
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_467
timestamp 1670771148
transform 1 0 44068 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_479
timestamp 1670771148
transform 1 0 45172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_499
timestamp 1670771148
transform 1 0 47012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1670771148
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1670771148
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_523
timestamp 1670771148
transform 1 0 49220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_527
timestamp 1670771148
transform 1 0 49588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_530
timestamp 1670771148
transform 1 0 49864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_538
timestamp 1670771148
transform 1 0 50600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_558
timestamp 1670771148
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_561
timestamp 1670771148
transform 1 0 52716 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_571
timestamp 1670771148
transform 1 0 53636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_591
timestamp 1670771148
transform 1 0 55476 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_597
timestamp 1670771148
transform 1 0 56028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_614
timestamp 1670771148
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1670771148
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_622
timestamp 1670771148
transform 1 0 58328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_630
timestamp 1670771148
transform 1 0 59064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_650
timestamp 1670771148
transform 1 0 60904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_670
timestamp 1670771148
transform 1 0 62744 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_673
timestamp 1670771148
transform 1 0 63020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_677
timestamp 1670771148
transform 1 0 63388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_685
timestamp 1670771148
transform 1 0 64124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_693
timestamp 1670771148
transform 1 0 64860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_701
timestamp 1670771148
transform 1 0 65596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_709
timestamp 1670771148
transform 1 0 66332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_713
timestamp 1670771148
transform 1 0 66700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_718
timestamp 1670771148
transform 1 0 67160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_726
timestamp 1670771148
transform 1 0 67896 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_729
timestamp 1670771148
transform 1 0 68172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_747
timestamp 1670771148
transform 1 0 69828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_751
timestamp 1670771148
transform 1 0 70196 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_754
timestamp 1670771148
transform 1 0 70472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_774
timestamp 1670771148
transform 1 0 72312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_782
timestamp 1670771148
transform 1 0 73048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_785
timestamp 1670771148
transform 1 0 73324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_789
timestamp 1670771148
transform 1 0 73692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_794
timestamp 1670771148
transform 1 0 74152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_802
timestamp 1670771148
transform 1 0 74888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_806
timestamp 1670771148
transform 1 0 75256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_811
timestamp 1670771148
transform 1 0 75716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_823
timestamp 1670771148
transform 1 0 76820 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_835
timestamp 1670771148
transform 1 0 77924 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1670771148
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_841
timestamp 1670771148
transform 1 0 78476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_847
timestamp 1670771148
transform 1 0 79028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_853
timestamp 1670771148
transform 1 0 79580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_859
timestamp 1670771148
transform 1 0 80132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_865
timestamp 1670771148
transform 1 0 80684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_885
timestamp 1670771148
transform 1 0 82524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_893
timestamp 1670771148
transform 1 0 83260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_897
timestamp 1670771148
transform 1 0 83628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_903
timestamp 1670771148
transform 1 0 84180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_909
timestamp 1670771148
transform 1 0 84732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_918
timestamp 1670771148
transform 1 0 85560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_922
timestamp 1670771148
transform 1 0 85928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_939
timestamp 1670771148
transform 1 0 87492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_947
timestamp 1670771148
transform 1 0 88228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1670771148
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_953
timestamp 1670771148
transform 1 0 88780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_959
timestamp 1670771148
transform 1 0 89332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_967
timestamp 1670771148
transform 1 0 90068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_976
timestamp 1670771148
transform 1 0 90896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_996
timestamp 1670771148
transform 1 0 92736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1004
timestamp 1670771148
transform 1 0 93472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1009
timestamp 1670771148
transform 1 0 93932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1015
timestamp 1670771148
transform 1 0 94484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1021
timestamp 1670771148
transform 1 0 95036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1041
timestamp 1670771148
transform 1 0 96876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1049
timestamp 1670771148
transform 1 0 97612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1057
timestamp 1670771148
transform 1 0 98348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1063
timestamp 1670771148
transform 1 0 98900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1065
timestamp 1670771148
transform 1 0 99084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1072
timestamp 1670771148
transform 1 0 99728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1080
timestamp 1670771148
transform 1 0 100464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1088
timestamp 1670771148
transform 1 0 101200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1096
timestamp 1670771148
transform 1 0 101936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1104
timestamp 1670771148
transform 1 0 102672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1112
timestamp 1670771148
transform 1 0 103408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1118
timestamp 1670771148
transform 1 0 103960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1121
timestamp 1670771148
transform 1 0 104236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1127
timestamp 1670771148
transform 1 0 104788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1135
timestamp 1670771148
transform 1 0 105524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1152
timestamp 1670771148
transform 1 0 107088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1160
timestamp 1670771148
transform 1 0 107824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1168
timestamp 1670771148
transform 1 0 108560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1174
timestamp 1670771148
transform 1 0 109112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1177
timestamp 1670771148
transform 1 0 109388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1183
timestamp 1670771148
transform 1 0 109940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1189
timestamp 1670771148
transform 1 0 110492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1193
timestamp 1670771148
transform 1 0 110860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1210
timestamp 1670771148
transform 1 0 112424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1218
timestamp 1670771148
transform 1 0 113160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1226
timestamp 1670771148
transform 1 0 113896 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1233
timestamp 1670771148
transform 1 0 114540 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1251
timestamp 1670771148
transform 1 0 116196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1271
timestamp 1670771148
transform 1 0 118036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1279
timestamp 1670771148
transform 1 0 118772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1285
timestamp 1670771148
transform 1 0 119324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1289
timestamp 1670771148
transform 1 0 119692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1295
timestamp 1670771148
transform 1 0 120244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1303
timestamp 1670771148
transform 1 0 120980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1311
timestamp 1670771148
transform 1 0 121716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1315
timestamp 1670771148
transform 1 0 122084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1332
timestamp 1670771148
transform 1 0 123648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1340
timestamp 1670771148
transform 1 0 124384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1345
timestamp 1670771148
transform 1 0 124844 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1351
timestamp 1670771148
transform 1 0 125396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1359
timestamp 1670771148
transform 1 0 126132 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1383
timestamp 1670771148
transform 1 0 128340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1391
timestamp 1670771148
transform 1 0 129076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1397
timestamp 1670771148
transform 1 0 129628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1401
timestamp 1670771148
transform 1 0 129996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1407
timestamp 1670771148
transform 1 0 130548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1415
timestamp 1670771148
transform 1 0 131284 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1423
timestamp 1670771148
transform 1 0 132020 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1441
timestamp 1670771148
transform 1 0 133676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1449
timestamp 1670771148
transform 1 0 134412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1455
timestamp 1670771148
transform 1 0 134964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1457
timestamp 1670771148
transform 1 0 135148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1463
timestamp 1670771148
transform 1 0 135700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1469
timestamp 1670771148
transform 1 0 136252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1477
timestamp 1670771148
transform 1 0 136988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1489
timestamp 1670771148
transform 1 0 138092 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1499
timestamp 1670771148
transform 1 0 139012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1507
timestamp 1670771148
transform 1 0 139748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1511
timestamp 1670771148
transform 1 0 140116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1513
timestamp 1670771148
transform 1 0 140300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1535
timestamp 1670771148
transform 1 0 142324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1543
timestamp 1670771148
transform 1 0 143060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1549
timestamp 1670771148
transform 1 0 143612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1566
timestamp 1670771148
transform 1 0 145176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1569
timestamp 1670771148
transform 1 0 145452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1587
timestamp 1670771148
transform 1 0 147108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1607
timestamp 1670771148
transform 1 0 148948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1615
timestamp 1670771148
transform 1 0 149684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1622
timestamp 1670771148
transform 1 0 150328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1625
timestamp 1670771148
transform 1 0 150604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1643
timestamp 1670771148
transform 1 0 152260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1663
timestamp 1670771148
transform 1 0 154100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1672
timestamp 1670771148
transform 1 0 154928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1678
timestamp 1670771148
transform 1 0 155480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1681
timestamp 1670771148
transform 1 0 155756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1687
timestamp 1670771148
transform 1 0 156308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1695
timestamp 1670771148
transform 1 0 157044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1702
timestamp 1670771148
transform 1 0 157688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1709
timestamp 1670771148
transform 1 0 158332 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1670771148
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1670771148
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1670771148
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1670771148
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1670771148
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1670771148
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_57
timestamp 1670771148
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1670771148
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1670771148
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1670771148
transform 1 0 7912 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1670771148
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1670771148
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1670771148
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1670771148
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1670771148
transform 1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1670771148
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1670771148
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1670771148
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1670771148
transform 1 0 12328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1670771148
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1670771148
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1670771148
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1670771148
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_163
timestamp 1670771148
transform 1 0 16100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1670771148
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp 1670771148
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1670771148
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1670771148
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1670771148
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1670771148
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1670771148
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1670771148
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1670771148
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_214
timestamp 1670771148
transform 1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_222
timestamp 1670771148
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1670771148
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_229
timestamp 1670771148
transform 1 0 22172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1670771148
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1670771148
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1670771148
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1670771148
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1670771148
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_278
timestamp 1670771148
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_281
timestamp 1670771148
transform 1 0 26956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_285
timestamp 1670771148
transform 1 0 27324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_290
timestamp 1670771148
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_298
timestamp 1670771148
transform 1 0 28520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1670771148
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_309
timestamp 1670771148
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_315
timestamp 1670771148
transform 1 0 30084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1670771148
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_337
timestamp 1670771148
transform 1 0 32108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_341
timestamp 1670771148
transform 1 0 32476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1670771148
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_354
timestamp 1670771148
transform 1 0 33672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1670771148
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1670771148
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_383
timestamp 1670771148
transform 1 0 36340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_387
timestamp 1670771148
transform 1 0 36708 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_390
timestamp 1670771148
transform 1 0 36984 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_393
timestamp 1670771148
transform 1 0 37260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_397
timestamp 1670771148
transform 1 0 37628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_402
timestamp 1670771148
transform 1 0 38088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_410
timestamp 1670771148
transform 1 0 38824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1670771148
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1670771148
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_428
timestamp 1670771148
transform 1 0 40480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_432
timestamp 1670771148
transform 1 0 40848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_437
timestamp 1670771148
transform 1 0 41308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_446
timestamp 1670771148
transform 1 0 42136 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_449
timestamp 1670771148
transform 1 0 42412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_454
timestamp 1670771148
transform 1 0 42872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1670771148
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1670771148
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_495
timestamp 1670771148
transform 1 0 46644 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_499
timestamp 1670771148
transform 1 0 47012 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_502
timestamp 1670771148
transform 1 0 47288 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_505
timestamp 1670771148
transform 1 0 47564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_510
timestamp 1670771148
transform 1 0 48024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_530
timestamp 1670771148
transform 1 0 49864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_533
timestamp 1670771148
transform 1 0 50140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_538
timestamp 1670771148
transform 1 0 50600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_558
timestamp 1670771148
transform 1 0 52440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_561
timestamp 1670771148
transform 1 0 52716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_566
timestamp 1670771148
transform 1 0 53176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_586
timestamp 1670771148
transform 1 0 55016 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_589
timestamp 1670771148
transform 1 0 55292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_594
timestamp 1670771148
transform 1 0 55752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_614
timestamp 1670771148
transform 1 0 57592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_617
timestamp 1670771148
transform 1 0 57868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_622
timestamp 1670771148
transform 1 0 58328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_642
timestamp 1670771148
transform 1 0 60168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_645
timestamp 1670771148
transform 1 0 60444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_665
timestamp 1670771148
transform 1 0 62284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_671
timestamp 1670771148
transform 1 0 62836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_673
timestamp 1670771148
transform 1 0 63020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_681
timestamp 1670771148
transform 1 0 63756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_685
timestamp 1670771148
transform 1 0 64124 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_688
timestamp 1670771148
transform 1 0 64400 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_698
timestamp 1670771148
transform 1 0 65320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_701
timestamp 1670771148
transform 1 0 65596 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_707
timestamp 1670771148
transform 1 0 66148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_717
timestamp 1670771148
transform 1 0 67068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_721
timestamp 1670771148
transform 1 0 67436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_726
timestamp 1670771148
transform 1 0 67896 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_729
timestamp 1670771148
transform 1 0 68172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_733
timestamp 1670771148
transform 1 0 68540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_738
timestamp 1670771148
transform 1 0 69000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_746
timestamp 1670771148
transform 1 0 69736 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_754
timestamp 1670771148
transform 1 0 70472 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_757
timestamp 1670771148
transform 1 0 70748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_761
timestamp 1670771148
transform 1 0 71116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_766
timestamp 1670771148
transform 1 0 71576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_774
timestamp 1670771148
transform 1 0 72312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_782
timestamp 1670771148
transform 1 0 73048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_785
timestamp 1670771148
transform 1 0 73324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_789
timestamp 1670771148
transform 1 0 73692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_794
timestamp 1670771148
transform 1 0 74152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_802
timestamp 1670771148
transform 1 0 74888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_810
timestamp 1670771148
transform 1 0 75624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_813
timestamp 1670771148
transform 1 0 75900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_819
timestamp 1670771148
transform 1 0 76452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_829
timestamp 1670771148
transform 1 0 77372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_833
timestamp 1670771148
transform 1 0 77740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_838
timestamp 1670771148
transform 1 0 78200 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_841
timestamp 1670771148
transform 1 0 78476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_849
timestamp 1670771148
transform 1 0 79212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_857
timestamp 1670771148
transform 1 0 79948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_865
timestamp 1670771148
transform 1 0 80684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_869
timestamp 1670771148
transform 1 0 81052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_875
timestamp 1670771148
transform 1 0 81604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_883
timestamp 1670771148
transform 1 0 82340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_891
timestamp 1670771148
transform 1 0 83076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_895
timestamp 1670771148
transform 1 0 83444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_897
timestamp 1670771148
transform 1 0 83628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_903
timestamp 1670771148
transform 1 0 84180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_911
timestamp 1670771148
transform 1 0 84916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_919
timestamp 1670771148
transform 1 0 85652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1670771148
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_925
timestamp 1670771148
transform 1 0 86204 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_929
timestamp 1670771148
transform 1 0 86572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_933
timestamp 1670771148
transform 1 0 86940 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_950
timestamp 1670771148
transform 1 0 88504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_953
timestamp 1670771148
transform 1 0 88780 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_957
timestamp 1670771148
transform 1 0 89148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_961
timestamp 1670771148
transform 1 0 89516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_968
timestamp 1670771148
transform 1 0 90160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_976
timestamp 1670771148
transform 1 0 90896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_981
timestamp 1670771148
transform 1 0 91356 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1001
timestamp 1670771148
transform 1 0 93196 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1007
timestamp 1670771148
transform 1 0 93748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1009
timestamp 1670771148
transform 1 0 93932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1015
timestamp 1670771148
transform 1 0 94484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1023
timestamp 1670771148
transform 1 0 95220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1031
timestamp 1670771148
transform 1 0 95956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1035
timestamp 1670771148
transform 1 0 96324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1037
timestamp 1670771148
transform 1 0 96508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1043
timestamp 1670771148
transform 1 0 97060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1051
timestamp 1670771148
transform 1 0 97796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1059
timestamp 1670771148
transform 1 0 98532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1063
timestamp 1670771148
transform 1 0 98900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1065
timestamp 1670771148
transform 1 0 99084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1071
timestamp 1670771148
transform 1 0 99636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1079
timestamp 1670771148
transform 1 0 100372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1087
timestamp 1670771148
transform 1 0 101108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1091
timestamp 1670771148
transform 1 0 101476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1093
timestamp 1670771148
transform 1 0 101660 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1104
timestamp 1670771148
transform 1 0 102672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1112
timestamp 1670771148
transform 1 0 103408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1118
timestamp 1670771148
transform 1 0 103960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1121
timestamp 1670771148
transform 1 0 104236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1127
timestamp 1670771148
transform 1 0 104788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1135
timestamp 1670771148
transform 1 0 105524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1143
timestamp 1670771148
transform 1 0 106260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1670771148
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1149
timestamp 1670771148
transform 1 0 106812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1153
timestamp 1670771148
transform 1 0 107180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1157
timestamp 1670771148
transform 1 0 107548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1174
timestamp 1670771148
transform 1 0 109112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1177
timestamp 1670771148
transform 1 0 109388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1183
timestamp 1670771148
transform 1 0 109940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1191
timestamp 1670771148
transform 1 0 110676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1199
timestamp 1670771148
transform 1 0 111412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1203
timestamp 1670771148
transform 1 0 111780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1205
timestamp 1670771148
transform 1 0 111964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1211
timestamp 1670771148
transform 1 0 112516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1219
timestamp 1670771148
transform 1 0 113252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1227
timestamp 1670771148
transform 1 0 113988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1231
timestamp 1670771148
transform 1 0 114356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1233
timestamp 1670771148
transform 1 0 114540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1239
timestamp 1670771148
transform 1 0 115092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1247
timestamp 1670771148
transform 1 0 115828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1255
timestamp 1670771148
transform 1 0 116564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1259
timestamp 1670771148
transform 1 0 116932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1261
timestamp 1670771148
transform 1 0 117116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1267
timestamp 1670771148
transform 1 0 117668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1275
timestamp 1670771148
transform 1 0 118404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1283
timestamp 1670771148
transform 1 0 119140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1287
timestamp 1670771148
transform 1 0 119508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1289
timestamp 1670771148
transform 1 0 119692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1295
timestamp 1670771148
transform 1 0 120244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1303
timestamp 1670771148
transform 1 0 120980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1311
timestamp 1670771148
transform 1 0 121716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1315
timestamp 1670771148
transform 1 0 122084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1317
timestamp 1670771148
transform 1 0 122268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1335
timestamp 1670771148
transform 1 0 123924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1341
timestamp 1670771148
transform 1 0 124476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1345
timestamp 1670771148
transform 1 0 124844 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1351
timestamp 1670771148
transform 1 0 125396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1359
timestamp 1670771148
transform 1 0 126132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1367
timestamp 1670771148
transform 1 0 126868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1371
timestamp 1670771148
transform 1 0 127236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1373
timestamp 1670771148
transform 1 0 127420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1379
timestamp 1670771148
transform 1 0 127972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1387
timestamp 1670771148
transform 1 0 128708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1395
timestamp 1670771148
transform 1 0 129444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1399
timestamp 1670771148
transform 1 0 129812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1401
timestamp 1670771148
transform 1 0 129996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1407
timestamp 1670771148
transform 1 0 130548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1415
timestamp 1670771148
transform 1 0 131284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1423
timestamp 1670771148
transform 1 0 132020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1427
timestamp 1670771148
transform 1 0 132388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1429
timestamp 1670771148
transform 1 0 132572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1435
timestamp 1670771148
transform 1 0 133124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1443
timestamp 1670771148
transform 1 0 133860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1451
timestamp 1670771148
transform 1 0 134596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1455
timestamp 1670771148
transform 1 0 134964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1457
timestamp 1670771148
transform 1 0 135148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1463
timestamp 1670771148
transform 1 0 135700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1471
timestamp 1670771148
transform 1 0 136436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1479
timestamp 1670771148
transform 1 0 137172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1483
timestamp 1670771148
transform 1 0 137540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1485
timestamp 1670771148
transform 1 0 137724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1491
timestamp 1670771148
transform 1 0 138276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1499
timestamp 1670771148
transform 1 0 139012 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1507
timestamp 1670771148
transform 1 0 139748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1511
timestamp 1670771148
transform 1 0 140116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1513
timestamp 1670771148
transform 1 0 140300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1519
timestamp 1670771148
transform 1 0 140852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1527
timestamp 1670771148
transform 1 0 141588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1535
timestamp 1670771148
transform 1 0 142324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1539
timestamp 1670771148
transform 1 0 142692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1541
timestamp 1670771148
transform 1 0 142876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1545
timestamp 1670771148
transform 1 0 143244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1549
timestamp 1670771148
transform 1 0 143612 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1566
timestamp 1670771148
transform 1 0 145176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1569
timestamp 1670771148
transform 1 0 145452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1573
timestamp 1670771148
transform 1 0 145820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1590
timestamp 1670771148
transform 1 0 147384 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1597
timestamp 1670771148
transform 1 0 148028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1615
timestamp 1670771148
transform 1 0 149684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1622
timestamp 1670771148
transform 1 0 150328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1625
timestamp 1670771148
transform 1 0 150604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1643
timestamp 1670771148
transform 1 0 152260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1650
timestamp 1670771148
transform 1 0 152904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1653
timestamp 1670771148
transform 1 0 153180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1659
timestamp 1670771148
transform 1 0 153732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1667
timestamp 1670771148
transform 1 0 154468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1675
timestamp 1670771148
transform 1 0 155204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1679
timestamp 1670771148
transform 1 0 155572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1681
timestamp 1670771148
transform 1 0 155756 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1687
timestamp 1670771148
transform 1 0 156308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1695
timestamp 1670771148
transform 1 0 157044 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1703
timestamp 1670771148
transform 1 0 157780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1707
timestamp 1670771148
transform 1 0 158148 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1709
timestamp 1670771148
transform 1 0 158332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1670771148
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1670771148
transform -1 0 158884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1670771148
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1670771148
transform -1 0 158884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1670771148
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1670771148
transform -1 0 158884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1670771148
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1670771148
transform -1 0 158884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1670771148
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1670771148
transform -1 0 158884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1670771148
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1670771148
transform -1 0 158884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1670771148
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1670771148
transform -1 0 158884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1670771148
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1670771148
transform -1 0 158884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1670771148
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1670771148
transform -1 0 158884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1670771148
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1670771148
transform -1 0 158884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1670771148
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1670771148
transform -1 0 158884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1670771148
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1670771148
transform -1 0 158884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1670771148
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1670771148
transform -1 0 158884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1670771148
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1670771148
transform -1 0 158884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1670771148
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1670771148
transform -1 0 158884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1670771148
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1670771148
transform -1 0 158884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1670771148
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1670771148
transform -1 0 158884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1670771148
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1670771148
transform -1 0 158884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1670771148
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1670771148
transform -1 0 158884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1670771148
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1670771148
transform -1 0 158884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1670771148
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1670771148
transform -1 0 158884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1670771148
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1670771148
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1670771148
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1670771148
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1670771148
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1670771148
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1670771148
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1670771148
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1670771148
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1670771148
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1670771148
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1670771148
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1670771148
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1670771148
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1670771148
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1670771148
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1670771148
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1670771148
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1670771148
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1670771148
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1670771148
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1670771148
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1670771148
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1670771148
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1670771148
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1670771148
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1670771148
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1670771148
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1670771148
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1670771148
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1670771148
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1670771148
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1670771148
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1670771148
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1670771148
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1670771148
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1670771148
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1670771148
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1670771148
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1670771148
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1670771148
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1670771148
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1670771148
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1670771148
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1670771148
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1670771148
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1670771148
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1670771148
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1670771148
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1670771148
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1670771148
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1670771148
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1670771148
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1670771148
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1670771148
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1670771148
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1670771148
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1670771148
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1670771148
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1670771148
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1670771148
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1670771148
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1670771148
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1670771148
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1670771148
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1670771148
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1670771148
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1670771148
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1670771148
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1670771148
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1670771148
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1670771148
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1670771148
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1670771148
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1670771148
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1670771148
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1670771148
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1670771148
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1670771148
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1670771148
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1670771148
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1670771148
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1670771148
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1670771148
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1670771148
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1670771148
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1670771148
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1670771148
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1670771148
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1670771148
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1670771148
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1670771148
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1670771148
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1670771148
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1670771148
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1670771148
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1670771148
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1670771148
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1670771148
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1670771148
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1670771148
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1670771148
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1670771148
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1670771148
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1670771148
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1670771148
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1670771148
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1670771148
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1670771148
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1670771148
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1670771148
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1670771148
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1670771148
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1670771148
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1670771148
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1670771148
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1670771148
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1670771148
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1670771148
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1670771148
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1670771148
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1670771148
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1670771148
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1670771148
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1670771148
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1670771148
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1670771148
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1670771148
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1670771148
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1670771148
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1670771148
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1670771148
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1670771148
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1670771148
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1670771148
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1670771148
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1670771148
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1670771148
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1670771148
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1670771148
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1670771148
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1670771148
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1670771148
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1670771148
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1670771148
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1670771148
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1670771148
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1670771148
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1670771148
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1670771148
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1670771148
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1670771148
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1670771148
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1670771148
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1670771148
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1670771148
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1670771148
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1670771148
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1670771148
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1670771148
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1670771148
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1670771148
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1670771148
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1670771148
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1670771148
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1670771148
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1670771148
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1670771148
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1670771148
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1670771148
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1670771148
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1670771148
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1670771148
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1670771148
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1670771148
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1670771148
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1670771148
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1670771148
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1670771148
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1670771148
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1670771148
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1670771148
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1670771148
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1670771148
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1670771148
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1670771148
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1670771148
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1670771148
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1670771148
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1670771148
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1670771148
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1670771148
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1670771148
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1670771148
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1670771148
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1670771148
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1670771148
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1670771148
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1670771148
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1670771148
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1670771148
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1670771148
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1670771148
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1670771148
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1670771148
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1670771148
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1670771148
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1670771148
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1670771148
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1670771148
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1670771148
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1670771148
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1670771148
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1670771148
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1670771148
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1670771148
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1670771148
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1670771148
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1670771148
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1670771148
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1670771148
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1670771148
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1670771148
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1670771148
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1670771148
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1670771148
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1670771148
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1670771148
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1670771148
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1670771148
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1670771148
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1670771148
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1670771148
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1670771148
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1670771148
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1670771148
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1670771148
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1670771148
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1670771148
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1670771148
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1670771148
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1670771148
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1670771148
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1670771148
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1670771148
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1670771148
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1670771148
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1670771148
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1670771148
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1670771148
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1670771148
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1670771148
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1670771148
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1670771148
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1670771148
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1670771148
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1670771148
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1670771148
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1670771148
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1670771148
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1670771148
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1670771148
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1670771148
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1670771148
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1670771148
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1670771148
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1670771148
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1670771148
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1670771148
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1670771148
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1670771148
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1670771148
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1670771148
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1670771148
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1670771148
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1670771148
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1670771148
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1670771148
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1670771148
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1670771148
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1670771148
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1670771148
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1670771148
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1670771148
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1670771148
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1670771148
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1670771148
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1670771148
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1670771148
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1670771148
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1670771148
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1670771148
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1670771148
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1670771148
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1670771148
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1670771148
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1670771148
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1670771148
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1670771148
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1670771148
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1670771148
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1670771148
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1670771148
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1670771148
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1670771148
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1670771148
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1670771148
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1670771148
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1670771148
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1670771148
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1670771148
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1670771148
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1670771148
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1670771148
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1670771148
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1670771148
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1670771148
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1670771148
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1670771148
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1670771148
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1670771148
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1670771148
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1670771148
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1670771148
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1670771148
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1670771148
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1670771148
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1670771148
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1670771148
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1670771148
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1670771148
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1670771148
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1670771148
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1670771148
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1670771148
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1670771148
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1670771148
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1670771148
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1670771148
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1670771148
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1670771148
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1670771148
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1670771148
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1670771148
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1670771148
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1670771148
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1670771148
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1670771148
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1670771148
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1670771148
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1670771148
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1670771148
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1670771148
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1670771148
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1670771148
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1670771148
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1670771148
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1670771148
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1670771148
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1670771148
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1670771148
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1670771148
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1670771148
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1670771148
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1670771148
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1670771148
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1670771148
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1670771148
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1670771148
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1670771148
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1670771148
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1670771148
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1670771148
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1670771148
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1670771148
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1670771148
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1670771148
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1670771148
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1670771148
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1670771148
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1670771148
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1670771148
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1670771148
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1670771148
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1670771148
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1670771148
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1670771148
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1670771148
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1670771148
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1670771148
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1670771148
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1670771148
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1670771148
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1670771148
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1670771148
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1670771148
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1670771148
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1670771148
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1670771148
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1670771148
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1670771148
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1670771148
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1670771148
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1670771148
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1670771148
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1670771148
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1670771148
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1670771148
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1670771148
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1670771148
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1670771148
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1670771148
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1670771148
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1670771148
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1670771148
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1670771148
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1670771148
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1670771148
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1670771148
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1670771148
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1670771148
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1670771148
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1670771148
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1670771148
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1670771148
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1670771148
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1670771148
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1670771148
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1670771148
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1670771148
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1670771148
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1670771148
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1670771148
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1670771148
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1670771148
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1670771148
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1670771148
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1670771148
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1670771148
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1670771148
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1670771148
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1670771148
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1670771148
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1670771148
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1670771148
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1670771148
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1670771148
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1670771148
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1670771148
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1670771148
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1670771148
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1670771148
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1670771148
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1670771148
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1670771148
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1670771148
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1670771148
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1670771148
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1670771148
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1670771148
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1670771148
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1670771148
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1670771148
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1670771148
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1670771148
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1670771148
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1670771148
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1670771148
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1670771148
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1670771148
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1670771148
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1670771148
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1670771148
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1670771148
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1670771148
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1670771148
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1670771148
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1670771148
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1670771148
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1670771148
transform 1 0 122176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1670771148
transform 1 0 127328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1670771148
transform 1 0 132480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1670771148
transform 1 0 137632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1670771148
transform 1 0 142784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1670771148
transform 1 0 147936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1670771148
transform 1 0 153088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1670771148
transform 1 0 158240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1670771148
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1670771148
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1670771148
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1670771148
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1670771148
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1670771148
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1670771148
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1670771148
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1670771148
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1670771148
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1670771148
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1670771148
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1670771148
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1670771148
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1670771148
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1670771148
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1670771148
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1670771148
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1670771148
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1670771148
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1670771148
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1670771148
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1670771148
transform 1 0 119600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1670771148
transform 1 0 124752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1670771148
transform 1 0 129904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1670771148
transform 1 0 135056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1670771148
transform 1 0 140208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1670771148
transform 1 0 145360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1670771148
transform 1 0 150512 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1670771148
transform 1 0 155664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1670771148
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1670771148
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1670771148
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1670771148
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1670771148
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1670771148
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1670771148
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1670771148
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1670771148
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1670771148
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1670771148
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1670771148
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1670771148
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1670771148
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1670771148
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1670771148
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1670771148
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1670771148
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1670771148
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1670771148
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1670771148
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1670771148
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1670771148
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1670771148
transform 1 0 122176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1670771148
transform 1 0 127328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1670771148
transform 1 0 132480 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1670771148
transform 1 0 137632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1670771148
transform 1 0 142784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1670771148
transform 1 0 147936 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1670771148
transform 1 0 153088 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1670771148
transform 1 0 158240 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1670771148
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1670771148
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1670771148
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1670771148
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1670771148
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1670771148
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1670771148
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1670771148
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1670771148
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1670771148
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1670771148
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1670771148
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1670771148
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1670771148
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1670771148
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1670771148
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1670771148
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1670771148
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1670771148
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1670771148
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1670771148
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1670771148
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1670771148
transform 1 0 119600 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1670771148
transform 1 0 124752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1670771148
transform 1 0 129904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1670771148
transform 1 0 135056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1670771148
transform 1 0 140208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1670771148
transform 1 0 145360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1670771148
transform 1 0 150512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1670771148
transform 1 0 155664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1670771148
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1670771148
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1670771148
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1670771148
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1670771148
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1670771148
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1670771148
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1670771148
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1670771148
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1670771148
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1670771148
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1670771148
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1670771148
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1670771148
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1670771148
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1670771148
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1670771148
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1670771148
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1670771148
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1670771148
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1670771148
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1670771148
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1670771148
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1670771148
transform 1 0 122176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1670771148
transform 1 0 127328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1670771148
transform 1 0 132480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1670771148
transform 1 0 137632 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1670771148
transform 1 0 142784 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1670771148
transform 1 0 147936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1670771148
transform 1 0 153088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1670771148
transform 1 0 158240 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1670771148
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1670771148
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1670771148
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1670771148
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1670771148
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1670771148
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1670771148
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1670771148
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1670771148
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1670771148
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1670771148
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1670771148
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1670771148
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1670771148
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1670771148
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1670771148
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1670771148
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1670771148
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1670771148
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1670771148
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1670771148
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1670771148
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1670771148
transform 1 0 119600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1670771148
transform 1 0 124752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1670771148
transform 1 0 129904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1670771148
transform 1 0 135056 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1670771148
transform 1 0 140208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1670771148
transform 1 0 145360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1670771148
transform 1 0 150512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1670771148
transform 1 0 155664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1670771148
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1670771148
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1670771148
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1670771148
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1670771148
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1670771148
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1670771148
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1670771148
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1670771148
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1670771148
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1670771148
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1670771148
transform 1 0 32016 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1670771148
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1670771148
transform 1 0 37168 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1670771148
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1670771148
transform 1 0 42320 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1670771148
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1670771148
transform 1 0 47472 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1670771148
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1670771148
transform 1 0 52624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1670771148
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1670771148
transform 1 0 57776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1670771148
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1670771148
transform 1 0 62928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1670771148
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1670771148
transform 1 0 68080 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1670771148
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1670771148
transform 1 0 73232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1670771148
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1670771148
transform 1 0 78384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1670771148
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1670771148
transform 1 0 83536 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1670771148
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1670771148
transform 1 0 88688 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1670771148
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1670771148
transform 1 0 93840 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1670771148
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1670771148
transform 1 0 98992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1670771148
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1670771148
transform 1 0 104144 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1670771148
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1670771148
transform 1 0 109296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1670771148
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1670771148
transform 1 0 114448 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1670771148
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1670771148
transform 1 0 119600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1670771148
transform 1 0 122176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1670771148
transform 1 0 124752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1670771148
transform 1 0 127328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1670771148
transform 1 0 129904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1670771148
transform 1 0 132480 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1670771148
transform 1 0 135056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1670771148
transform 1 0 137632 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1670771148
transform 1 0 140208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1670771148
transform 1 0 142784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1670771148
transform 1 0 145360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1670771148
transform 1 0 147936 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1670771148
transform 1 0 150512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1670771148
transform 1 0 153088 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1670771148
transform 1 0 155664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1670771148
transform 1 0 158240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0540_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 12788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0541_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 16836 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0542_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0543_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 5980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0544_
timestamp 1670771148
transform -1 0 15272 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1670771148
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0546_
timestamp 1670771148
transform 1 0 14904 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0547_
timestamp 1670771148
transform 1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0548_
timestamp 1670771148
transform 1 0 17020 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1670771148
transform -1 0 18952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0550_
timestamp 1670771148
transform -1 0 18768 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1670771148
transform -1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0552_
timestamp 1670771148
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1670771148
transform -1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0554_
timestamp 1670771148
transform 1 0 25300 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1670771148
transform -1 0 26128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0556_
timestamp 1670771148
transform -1 0 24380 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1670771148
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0558_
timestamp 1670771148
transform 1 0 21988 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1670771148
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0560_
timestamp 1670771148
transform 1 0 25760 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1670771148
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0562_
timestamp 1670771148
transform -1 0 20148 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1670771148
transform 1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0564_
timestamp 1670771148
transform -1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0565_
timestamp 1670771148
transform -1 0 5704 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1670771148
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0567_
timestamp 1670771148
transform -1 0 6992 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1670771148
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0569_
timestamp 1670771148
transform -1 0 5244 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1670771148
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0571_
timestamp 1670771148
transform -1 0 4876 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1670771148
transform 1 0 4416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0573_
timestamp 1670771148
transform 1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1670771148
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0575_
timestamp 1670771148
transform -1 0 12328 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1670771148
transform -1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0577_
timestamp 1670771148
transform -1 0 8648 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1670771148
transform 1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0579_
timestamp 1670771148
transform -1 0 9568 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1670771148
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0581_
timestamp 1670771148
transform 1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1670771148
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0583_
timestamp 1670771148
transform 1 0 11408 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1670771148
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0585_
timestamp 1670771148
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0586_
timestamp 1670771148
transform -1 0 14720 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1670771148
transform -1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0588_
timestamp 1670771148
transform -1 0 13800 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1670771148
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0590_
timestamp 1670771148
transform -1 0 15824 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1670771148
transform -1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0592_
timestamp 1670771148
transform -1 0 16652 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1670771148
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0594_
timestamp 1670771148
transform 1 0 11224 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1670771148
transform -1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0596_
timestamp 1670771148
transform 1 0 17756 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1670771148
transform -1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0598_
timestamp 1670771148
transform -1 0 17388 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1670771148
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0600_
timestamp 1670771148
transform -1 0 13708 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0601_
timestamp 1670771148
transform -1 0 11224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0602_
timestamp 1670771148
transform -1 0 17112 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1670771148
transform -1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0604_
timestamp 1670771148
transform 1 0 18032 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0605_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 25668 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0606_
timestamp 1670771148
transform 1 0 32936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1670771148
transform -1 0 54372 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1670771148
transform 1 0 53544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0609_
timestamp 1670771148
transform -1 0 52072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1670771148
transform 1 0 48760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0611_
timestamp 1670771148
transform 1 0 45816 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1670771148
transform 1 0 46460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0613_
timestamp 1670771148
transform 1 0 49404 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1670771148
transform 1 0 50232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0615_
timestamp 1670771148
transform -1 0 45908 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1670771148
transform -1 0 41032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0617_
timestamp 1670771148
transform 1 0 40480 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1670771148
transform -1 0 45264 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0619_
timestamp 1670771148
transform -1 0 37444 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1670771148
transform 1 0 36708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0621_
timestamp 1670771148
transform -1 0 45816 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1670771148
transform 1 0 41124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1670771148
transform -1 0 40480 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1670771148
transform 1 0 38364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0625_
timestamp 1670771148
transform 1 0 37812 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1670771148
transform 1 0 39100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0627_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 101936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0628_
timestamp 1670771148
transform -1 0 67068 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 1670771148
transform 1 0 29256 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1670771148
transform 1 0 33304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0631_
timestamp 1670771148
transform 1 0 33488 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1670771148
transform -1 0 38088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0633_
timestamp 1670771148
transform 1 0 33304 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1670771148
transform -1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1670771148
transform -1 0 37168 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1670771148
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0637_
timestamp 1670771148
transform -1 0 34040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1670771148
transform 1 0 31556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0639_
timestamp 1670771148
transform 1 0 29900 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1670771148
transform 1 0 30728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 1670771148
transform 1 0 32292 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1670771148
transform 1 0 32568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0643_
timestamp 1670771148
transform 1 0 30636 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1670771148
transform 1 0 33488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 1670771148
transform 1 0 26588 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0646_
timestamp 1670771148
transform -1 0 27416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0647_
timestamp 1670771148
transform 1 0 33672 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1670771148
transform -1 0 36800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0649_
timestamp 1670771148
transform -1 0 77372 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0650_
timestamp 1670771148
transform -1 0 40480 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1670771148
transform -1 0 39560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1670771148
transform 1 0 42688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1670771148
transform 1 0 44436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1670771148
transform 1 0 43516 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0655_
timestamp 1670771148
transform 1 0 46092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1670771148
transform 1 0 47196 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1670771148
transform 1 0 47748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0658_
timestamp 1670771148
transform -1 0 47196 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1670771148
transform -1 0 45448 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1670771148
transform -1 0 36800 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1670771148
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1670771148
transform 1 0 40204 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1670771148
transform -1 0 41492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0664_
timestamp 1670771148
transform 1 0 46828 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1670771148
transform -1 0 48024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0666_
timestamp 1670771148
transform 1 0 51428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1670771148
transform 1 0 54004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0668_
timestamp 1670771148
transform -1 0 45816 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1670771148
transform -1 0 42320 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0670_
timestamp 1670771148
transform -1 0 65320 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1670771148
transform 1 0 48208 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1670771148
transform 1 0 48484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0673_
timestamp 1670771148
transform -1 0 58880 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1670771148
transform 1 0 57040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0675_
timestamp 1670771148
transform -1 0 41676 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1670771148
transform -1 0 40756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0677_
timestamp 1670771148
transform 1 0 41676 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1670771148
transform -1 0 42872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0679_
timestamp 1670771148
transform 1 0 50784 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1670771148
transform -1 0 56488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0681_
timestamp 1670771148
transform 1 0 51704 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0682_
timestamp 1670771148
transform -1 0 53084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1670771148
transform -1 0 66240 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1670771148
transform 1 0 64860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0685_
timestamp 1670771148
transform -1 0 59708 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0686_
timestamp 1670771148
transform 1 0 58420 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0687_
timestamp 1670771148
transform -1 0 52440 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1670771148
transform 1 0 50692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0689_
timestamp 1670771148
transform 1 0 54464 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1670771148
transform -1 0 56764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0691_
timestamp 1670771148
transform -1 0 64860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1670771148
transform -1 0 56856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1670771148
transform -1 0 55752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0694_
timestamp 1670771148
transform -1 0 58880 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1670771148
transform 1 0 55936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1670771148
transform 1 0 51796 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1670771148
transform 1 0 52900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1670771148
transform -1 0 59708 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1670771148
transform 1 0 58052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0700_
timestamp 1670771148
transform -1 0 60904 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1670771148
transform 1 0 58052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1670771148
transform 1 0 63296 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1670771148
transform -1 0 64768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1670771148
transform 1 0 63664 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0705_
timestamp 1670771148
transform -1 0 64860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0706_
timestamp 1670771148
transform -1 0 54096 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1670771148
transform 1 0 53176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0708_
timestamp 1670771148
transform 1 0 54280 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1670771148
transform 1 0 54740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0710_
timestamp 1670771148
transform -1 0 57592 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1670771148
transform 1 0 56488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0712_
timestamp 1670771148
transform -1 0 66148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1670771148
transform -1 0 55936 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 1670771148
transform -1 0 55384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1670771148
transform -1 0 65136 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1670771148
transform -1 0 63848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1670771148
transform -1 0 67896 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0718_
timestamp 1670771148
transform 1 0 67436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1670771148
transform 1 0 56764 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1670771148
transform 1 0 57316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0721_
timestamp 1670771148
transform -1 0 60904 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1670771148
transform -1 0 60812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0723_
timestamp 1670771148
transform 1 0 63020 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0724_
timestamp 1670771148
transform 1 0 63204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 1670771148
transform -1 0 70196 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0726_
timestamp 1670771148
transform -1 0 67160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0727_
timestamp 1670771148
transform 1 0 72312 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0728_
timestamp 1670771148
transform -1 0 77280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0729_
timestamp 1670771148
transform -1 0 73968 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0730_
timestamp 1670771148
transform -1 0 73416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 1670771148
transform -1 0 68816 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0732_
timestamp 1670771148
transform 1 0 66608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1670771148
transform -1 0 74152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1670771148
transform 1 0 73508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1670771148
transform -1 0 79672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1670771148
transform -1 0 73140 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1670771148
transform 1 0 67620 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0738_
timestamp 1670771148
transform -1 0 76544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1670771148
transform 1 0 74888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0740_
timestamp 1670771148
transform 1 0 82340 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 1670771148
transform -1 0 84548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0742_
timestamp 1670771148
transform -1 0 87860 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1670771148
transform -1 0 87032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0744_
timestamp 1670771148
transform -1 0 82432 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0745_
timestamp 1670771148
transform 1 0 78844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0746_
timestamp 1670771148
transform -1 0 76544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 1670771148
transform 1 0 76084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1670771148
transform 1 0 74428 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 1670771148
transform -1 0 75532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0750_
timestamp 1670771148
transform 1 0 82524 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1670771148
transform -1 0 84088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0752_
timestamp 1670771148
transform -1 0 84272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1670771148
transform 1 0 81880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0754_
timestamp 1670771148
transform -1 0 90160 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0755_
timestamp 1670771148
transform -1 0 85560 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0756_
timestamp 1670771148
transform 1 0 84456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp 1670771148
transform 1 0 107364 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0758_
timestamp 1670771148
transform 1 0 108192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1670771148
transform 1 0 98348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0760_
timestamp 1670771148
transform 1 0 98624 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1670771148
transform 1 0 81236 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1670771148
transform 1 0 82800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1670771148
transform 1 0 104328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1670771148
transform 1 0 105432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1670771148
transform -1 0 111504 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0766_
timestamp 1670771148
transform 1 0 110952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1670771148
transform -1 0 99728 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 1670771148
transform 1 0 97520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1670771148
transform 1 0 90436 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 1670771148
transform -1 0 98072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1670771148
transform 1 0 91908 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1670771148
transform -1 0 93380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1670771148
transform 1 0 94116 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1670771148
transform 1 0 95128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0775_
timestamp 1670771148
transform 1 0 112332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0776_
timestamp 1670771148
transform -1 0 121164 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0777_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 119784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0778_
timestamp 1670771148
transform -1 0 118588 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0779_
timestamp 1670771148
transform 1 0 117944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1670771148
transform 1 0 116104 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0781_
timestamp 1670771148
transform 1 0 117668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0782_
timestamp 1670771148
transform 1 0 118588 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0783_
timestamp 1670771148
transform 1 0 123924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0784_
timestamp 1670771148
transform 1 0 121072 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0785_
timestamp 1670771148
transform -1 0 123188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0786_
timestamp 1670771148
transform 1 0 107732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 1670771148
transform 1 0 108744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0788_
timestamp 1670771148
transform 1 0 117944 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0789_
timestamp 1670771148
transform 1 0 118496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0790_
timestamp 1670771148
transform 1 0 114724 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0791_
timestamp 1670771148
transform -1 0 115736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0792_
timestamp 1670771148
transform 1 0 115460 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0793_
timestamp 1670771148
transform 1 0 118312 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0794_
timestamp 1670771148
transform 1 0 113252 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0795_
timestamp 1670771148
transform 1 0 117300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1670771148
transform 1 0 117208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0797_
timestamp 1670771148
transform -1 0 125488 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0798_
timestamp 1670771148
transform 1 0 125028 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0799_
timestamp 1670771148
transform -1 0 128892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0800_
timestamp 1670771148
transform 1 0 128524 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0801_
timestamp 1670771148
transform -1 0 114632 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0802_
timestamp 1670771148
transform 1 0 113896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0803_
timestamp 1670771148
transform 1 0 126132 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1670771148
transform 1 0 127788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0805_
timestamp 1670771148
transform -1 0 130640 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0806_
timestamp 1670771148
transform -1 0 130088 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0807_
timestamp 1670771148
transform -1 0 114264 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 1670771148
transform 1 0 112148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1670771148
transform -1 0 133216 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0810_
timestamp 1670771148
transform 1 0 132756 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 1670771148
transform 1 0 129720 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0812_
timestamp 1670771148
transform -1 0 130548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0813_
timestamp 1670771148
transform 1 0 131836 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0814_
timestamp 1670771148
transform 1 0 132756 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1670771148
transform -1 0 133216 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0816_
timestamp 1670771148
transform -1 0 133124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0817_
timestamp 1670771148
transform 1 0 119140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1670771148
transform 1 0 126960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0819_
timestamp 1670771148
transform 1 0 128524 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0820_
timestamp 1670771148
transform -1 0 128156 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0821_
timestamp 1670771148
transform -1 0 126868 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1670771148
transform 1 0 130732 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0823_
timestamp 1670771148
transform -1 0 132112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0824_
timestamp 1670771148
transform -1 0 121440 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1670771148
transform -1 0 120612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0826_
timestamp 1670771148
transform 1 0 118772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0827_
timestamp 1670771148
transform -1 0 119416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 1670771148
transform 1 0 126592 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0829_
timestamp 1670771148
transform -1 0 128156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1670771148
transform -1 0 128156 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0831_
timestamp 1670771148
transform 1 0 127788 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0832_
timestamp 1670771148
transform -1 0 122912 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0833_
timestamp 1670771148
transform -1 0 122820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0834_
timestamp 1670771148
transform -1 0 119232 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0835_
timestamp 1670771148
transform 1 0 118036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0836_
timestamp 1670771148
transform 1 0 125856 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0837_
timestamp 1670771148
transform -1 0 130640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0838_
timestamp 1670771148
transform 1 0 137448 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0839_
timestamp 1670771148
transform 1 0 150052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0840_
timestamp 1670771148
transform 1 0 154100 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 1670771148
transform 1 0 157596 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0842_
timestamp 1670771148
transform 1 0 149408 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0843_
timestamp 1670771148
transform 1 0 156584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0844_
timestamp 1670771148
transform 1 0 154560 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0845_
timestamp 1670771148
transform 1 0 157504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0846_
timestamp 1670771148
transform 1 0 155296 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1670771148
transform 1 0 157412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1670771148
transform -1 0 155756 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1670771148
transform 1 0 136344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1670771148
transform 1 0 156768 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1670771148
transform 1 0 156952 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0852_
timestamp 1670771148
transform 1 0 154468 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1670771148
transform 1 0 157596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0854_
timestamp 1670771148
transform 1 0 155940 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1670771148
transform 1 0 157412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1670771148
transform 1 0 154468 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1670771148
transform 1 0 158056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1670771148
transform -1 0 154376 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1670771148
transform 1 0 140392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1670771148
transform 1 0 147108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0861_
timestamp 1670771148
transform 1 0 156768 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0862_
timestamp 1670771148
transform 1 0 157228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0863_
timestamp 1670771148
transform -1 0 154928 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0864_
timestamp 1670771148
transform 1 0 153456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1670771148
transform -1 0 156400 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1670771148
transform 1 0 130180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0867_
timestamp 1670771148
transform -1 0 148672 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 1670771148
transform 1 0 141128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0869_
timestamp 1670771148
transform -1 0 156860 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1670771148
transform 1 0 155940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1670771148
transform -1 0 152536 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0872_
timestamp 1670771148
transform -1 0 152352 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0873_
timestamp 1670771148
transform 1 0 146740 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1670771148
transform 1 0 147476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1670771148
transform 1 0 151892 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0876_
timestamp 1670771148
transform -1 0 152352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1670771148
transform -1 0 142416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0878_
timestamp 1670771148
transform 1 0 141680 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0879_
timestamp 1670771148
transform 1 0 138552 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0880_
timestamp 1670771148
transform -1 0 142232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0881_
timestamp 1670771148
transform 1 0 152720 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1670771148
transform 1 0 113804 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0883_
timestamp 1670771148
transform 1 0 125948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1670771148
transform 1 0 118220 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0885_
timestamp 1670771148
transform 1 0 118312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1670771148
transform -1 0 121256 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1670771148
transform -1 0 119784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1670771148
transform -1 0 122912 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1670771148
transform 1 0 122452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0890_
timestamp 1670771148
transform 1 0 155020 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1670771148
transform 1 0 156768 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1670771148
transform 1 0 155940 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1670771148
transform 1 0 156768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1670771148
transform 1 0 156032 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1670771148
transform 1 0 156768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0896_
timestamp 1670771148
transform -1 0 155664 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1670771148
transform 1 0 152260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1670771148
transform 1 0 156768 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1670771148
transform 1 0 157596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1670771148
transform 1 0 156492 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1670771148
transform 1 0 157596 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0902_
timestamp 1670771148
transform 1 0 142048 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1670771148
transform -1 0 154928 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1670771148
transform 1 0 150052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0905_
timestamp 1670771148
transform 1 0 149316 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0906_
timestamp 1670771148
transform 1 0 150788 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1670771148
transform -1 0 125764 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1670771148
transform -1 0 108652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1670771148
transform -1 0 126408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1670771148
transform 1 0 125580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1670771148
transform 1 0 130548 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1670771148
transform -1 0 135608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1670771148
transform -1 0 141128 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1670771148
transform -1 0 140392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1670771148
transform 1 0 154744 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1670771148
transform 1 0 157596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1670771148
transform 1 0 154100 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1670771148
transform 1 0 156400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0919_
timestamp 1670771148
transform 1 0 154192 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0920_
timestamp 1670771148
transform 1 0 158056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1670771148
transform 1 0 153548 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0922_
timestamp 1670771148
transform 1 0 155112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1670771148
transform 1 0 135608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0924_
timestamp 1670771148
transform 1 0 155940 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 1670771148
transform 1 0 156768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1670771148
transform 1 0 156676 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1670771148
transform 1 0 156584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0928_
timestamp 1670771148
transform 1 0 147108 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1670771148
transform 1 0 150788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1670771148
transform 1 0 156124 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1670771148
transform 1 0 157504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1670771148
transform 1 0 154928 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 1670771148
transform 1 0 158056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0934_
timestamp 1670771148
transform 1 0 155940 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1670771148
transform -1 0 157320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1670771148
transform 1 0 154468 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1670771148
transform 1 0 158056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0938_
timestamp 1670771148
transform -1 0 145084 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1670771148
transform 1 0 141404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0940_
timestamp 1670771148
transform 1 0 140484 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1670771148
transform 1 0 140944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1670771148
transform -1 0 152720 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1670771148
transform 1 0 151432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1670771148
transform 1 0 140944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1670771148
transform 1 0 149316 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1670771148
transform 1 0 150052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1670771148
transform 1 0 155940 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1670771148
transform 1 0 156952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0949_
timestamp 1670771148
transform -1 0 155664 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1670771148
transform 1 0 151800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0951_
timestamp 1670771148
transform 1 0 155664 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1670771148
transform 1 0 157504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1670771148
transform -1 0 157228 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1670771148
transform 1 0 150052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0955_
timestamp 1670771148
transform -1 0 151248 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1670771148
transform 1 0 150052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1670771148
transform -1 0 141220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0958_
timestamp 1670771148
transform -1 0 139748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1670771148
transform -1 0 144440 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1670771148
transform -1 0 139840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1670771148
transform -1 0 156400 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1670771148
transform 1 0 150880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1670771148
transform 1 0 154192 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1670771148
transform 1 0 154376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0965_
timestamp 1670771148
transform 1 0 149316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0966_
timestamp 1670771148
transform 1 0 155940 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1670771148
transform 1 0 158056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1670771148
transform 1 0 155112 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 1670771148
transform 1 0 157412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1670771148
transform 1 0 155020 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1670771148
transform 1 0 157596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1670771148
transform 1 0 150052 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1670771148
transform 1 0 157412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1670771148
transform 1 0 151892 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 1670771148
transform 1 0 157320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0976_
timestamp 1670771148
transform -1 0 155204 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1670771148
transform 1 0 153456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1670771148
transform -1 0 156584 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1670771148
transform 1 0 122360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0980_
timestamp 1670771148
transform -1 0 141496 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1670771148
transform 1 0 137908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1670771148
transform -1 0 143520 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1670771148
transform 1 0 127236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0984_
timestamp 1670771148
transform 1 0 156768 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1670771148
transform 1 0 157412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0986_
timestamp 1670771148
transform 1 0 153548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0987_
timestamp 1670771148
transform 1 0 150604 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1670771148
transform 1 0 150788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0989_
timestamp 1670771148
transform -1 0 153824 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1670771148
transform 1 0 152628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1670771148
transform -1 0 152904 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1670771148
transform 1 0 151616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1670771148
transform 1 0 153364 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1670771148
transform 1 0 156860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1670771148
transform 1 0 152628 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1670771148
transform 1 0 155940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0997_
timestamp 1670771148
transform 1 0 152444 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1670771148
transform 1 0 152628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0999_
timestamp 1670771148
transform 1 0 151432 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1670771148
transform 1 0 152076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1670771148
transform -1 0 153548 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1670771148
transform 1 0 150788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1003_
timestamp 1670771148
transform 1 0 153640 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1670771148
transform 1 0 157228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1670771148
transform -1 0 156032 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1670771148
transform 1 0 151616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1007_
timestamp 1670771148
transform 1 0 149684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1670771148
transform -1 0 156308 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1670771148
transform -1 0 143796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1010_
timestamp 1670771148
transform -1 0 155388 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1670771148
transform 1 0 150052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1012_
timestamp 1670771148
transform -1 0 146096 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1670771148
transform -1 0 140576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1014_
timestamp 1670771148
transform -1 0 138644 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1670771148
transform -1 0 137080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1670771148
transform -1 0 141036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1670771148
transform -1 0 140024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1018_
timestamp 1670771148
transform 1 0 139012 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1670771148
transform 1 0 140300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1020_
timestamp 1670771148
transform -1 0 140668 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1670771148
transform 1 0 138368 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1022_
timestamp 1670771148
transform -1 0 147660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1670771148
transform -1 0 140760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1024_
timestamp 1670771148
transform -1 0 151248 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1670771148
transform 1 0 142968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1026_
timestamp 1670771148
transform -1 0 154100 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1027_
timestamp 1670771148
transform -1 0 153548 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1028_
timestamp 1670771148
transform -1 0 139932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1029_
timestamp 1670771148
transform -1 0 127144 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1670771148
transform 1 0 126684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1031_
timestamp 1670771148
transform 1 0 110400 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1670771148
transform 1 0 111320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1670771148
transform 1 0 110492 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1670771148
transform 1 0 115460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1670771148
transform -1 0 115000 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1670771148
transform 1 0 113620 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1037_
timestamp 1670771148
transform -1 0 114080 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1670771148
transform 1 0 113252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1039_
timestamp 1670771148
transform -1 0 111688 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1670771148
transform 1 0 110860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1041_
timestamp 1670771148
transform 1 0 104420 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1670771148
transform -1 0 105984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1043_
timestamp 1670771148
transform 1 0 110860 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 1670771148
transform 1 0 111412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1045_
timestamp 1670771148
transform -1 0 109204 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1670771148
transform 1 0 107916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1047_
timestamp 1670771148
transform 1 0 102212 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1670771148
transform 1 0 102764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1049_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 62560 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1050_
timestamp 1670771148
transform -1 0 97244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1670771148
transform 1 0 83996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1052_
timestamp 1670771148
transform -1 0 113068 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1670771148
transform 1 0 108100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1054_
timestamp 1670771148
transform 1 0 9108 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1670771148
transform -1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1056_
timestamp 1670771148
transform -1 0 30452 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1670771148
transform -1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1670771148
transform -1 0 23184 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1670771148
transform 1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 1670771148
transform 1 0 16928 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1670771148
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1062_
timestamp 1670771148
transform -1 0 16560 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1063_
timestamp 1670771148
transform 1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1064_
timestamp 1670771148
transform 1 0 14260 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1670771148
transform -1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1066_
timestamp 1670771148
transform 1 0 12788 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1067_
timestamp 1670771148
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1068_
timestamp 1670771148
transform 1 0 11684 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1069_
timestamp 1670771148
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1070_
timestamp 1670771148
transform 1 0 14996 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1071_
timestamp 1670771148
transform -1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1072_
timestamp 1670771148
transform 1 0 17756 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1073_
timestamp 1670771148
transform -1 0 20976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1670771148
transform 1 0 14996 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1670771148
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1076_
timestamp 1670771148
transform -1 0 16100 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1670771148
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1078_
timestamp 1670771148
transform 1 0 16836 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1670771148
transform 1 0 19596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1080_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1670771148
transform 1 0 12236 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1670771148
transform 1 0 16192 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1670771148
transform 1 0 21896 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1670771148
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1670771148
transform 1 0 22724 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1670771148
transform 1 0 27140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1670771148
transform 1 0 20148 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1670771148
transform 1 0 24564 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1670771148
transform -1 0 26404 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1670771148
transform -1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1670771148
transform 1 0 3772 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1670771148
transform 1 0 3956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1670771148
transform 1 0 3956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1670771148
transform 1 0 3772 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1670771148
transform -1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1670771148
transform 1 0 14352 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1097_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 3772 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1670771148
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1670771148
transform 1 0 13524 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1670771148
transform 1 0 3772 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1670771148
transform 1 0 13800 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1670771148
transform 1 0 11040 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1670771148
transform 1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1670771148
transform -1 0 13156 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1670771148
transform 1 0 12328 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1670771148
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1670771148
transform -1 0 15732 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1670771148
transform 1 0 14260 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1670771148
transform 1 0 17388 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1670771148
transform 1 0 50692 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1670771148
transform 1 0 46184 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1670771148
transform -1 0 44068 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1670771148
transform 1 0 37168 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1670771148
transform -1 0 49864 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1670771148
transform -1 0 41860 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1670771148
transform -1 0 55752 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1670771148
transform 1 0 36248 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1670771148
transform -1 0 39008 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1670771148
transform -1 0 36800 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1670771148
transform -1 0 36800 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1670771148
transform 1 0 32660 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1670771148
transform 1 0 38364 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1670771148
transform 1 0 38640 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1670771148
transform -1 0 34408 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1670771148
transform -1 0 31280 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1670771148
transform 1 0 29072 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1670771148
transform 1 0 27784 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1670771148
transform -1 0 29256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1670771148
transform 1 0 29716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1670771148
transform 1 0 39100 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1670771148
transform 1 0 42596 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1670771148
transform 1 0 42780 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1670771148
transform -1 0 44068 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1670771148
transform 1 0 45632 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1670771148
transform -1 0 46736 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1670771148
transform -1 0 33856 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1670771148
transform 1 0 45816 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1670771148
transform 1 0 47748 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1670771148
transform -1 0 53636 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1670771148
transform 1 0 43240 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1670771148
transform 1 0 43240 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1670771148
transform -1 0 52440 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1670771148
transform 1 0 40664 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1670771148
transform 1 0 43148 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1670771148
transform 1 0 56120 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1670771148
transform 1 0 63480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1670771148
transform -1 0 61824 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1670771148
transform -1 0 58604 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1670771148
transform 1 0 43240 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1670771148
transform -1 0 65320 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1670771148
transform -1 0 64768 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1670771148
transform -1 0 49220 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1670771148
transform 1 0 45908 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1670771148
transform 1 0 57684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1670771148
transform 1 0 50232 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1670771148
transform -1 0 76636 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1670771148
transform -1 0 65320 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1670771148
transform 1 0 52624 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1670771148
transform -1 0 52440 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1670771148
transform 1 0 54280 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1670771148
transform 1 0 58696 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1670771148
transform 1 0 63848 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1670771148
transform -1 0 62652 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1670771148
transform 1 0 56120 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1670771148
transform 1 0 60996 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1670771148
transform 1 0 60628 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1670771148
transform 1 0 67528 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1670771148
transform -1 0 78016 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1670771148
transform -1 0 73784 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1670771148
transform -1 0 65136 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1670771148
transform -1 0 93012 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1670771148
transform 1 0 65780 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1670771148
transform 1 0 72588 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1670771148
transform -1 0 89332 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1670771148
transform -1 0 93380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1670771148
transform -1 0 75532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1670771148
transform -1 0 75624 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp 1670771148
transform 1 0 89056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1670771148
transform 1 0 88780 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1670771148
transform 1 0 81236 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1670771148
transform 1 0 76728 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1670771148
transform -1 0 95956 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1670771148
transform -1 0 82892 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1670771148
transform 1 0 79304 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1670771148
transform -1 0 87860 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1670771148
transform -1 0 92276 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1670771148
transform -1 0 96876 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1670771148
transform -1 0 100832 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1670771148
transform -1 0 95404 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1670771148
transform 1 0 78292 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1191_
timestamp 1670771148
transform -1 0 75532 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1670771148
transform -1 0 115276 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1670771148
transform -1 0 108468 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1194_
timestamp 1670771148
transform -1 0 96232 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1670771148
transform 1 0 76084 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1196_
timestamp 1670771148
transform -1 0 90896 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1670771148
transform -1 0 109756 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1198_
timestamp 1670771148
transform -1 0 117392 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1670771148
transform -1 0 92736 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1200_
timestamp 1670771148
transform -1 0 116932 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1670771148
transform -1 0 103316 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1670771148
transform -1 0 100280 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1203_
timestamp 1670771148
transform -1 0 100188 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1204_
timestamp 1670771148
transform -1 0 121440 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1670771148
transform 1 0 104604 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1206_
timestamp 1670771148
transform -1 0 102120 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1207_
timestamp 1670771148
transform -1 0 105984 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1208_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 76268 0 -1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1209_
timestamp 1670771148
transform -1 0 103408 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1210_
timestamp 1670771148
transform -1 0 98256 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1211_
timestamp 1670771148
transform -1 0 101384 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1212_
timestamp 1670771148
transform -1 0 93932 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1213_
timestamp 1670771148
transform -1 0 94300 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1214_
timestamp 1670771148
transform 1 0 62100 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1670771148
transform 1 0 87124 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1216_
timestamp 1670771148
transform -1 0 86756 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1217_
timestamp 1670771148
transform -1 0 95864 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1218_
timestamp 1670771148
transform -1 0 73048 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp 1670771148
transform 1 0 96692 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1220_
timestamp 1670771148
transform 1 0 133400 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1221_
timestamp 1670771148
transform 1 0 145360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp 1670771148
transform 1 0 147476 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp 1670771148
transform 1 0 143336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1224_
timestamp 1670771148
transform -1 0 147752 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1225_
timestamp 1670771148
transform -1 0 120336 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1226_
timestamp 1670771148
transform -1 0 136620 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1227_
timestamp 1670771148
transform -1 0 138736 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1228_
timestamp 1670771148
transform -1 0 140208 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1229_
timestamp 1670771148
transform -1 0 145176 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1230_
timestamp 1670771148
transform -1 0 135608 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 1670771148
transform -1 0 145084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 1670771148
transform 1 0 147476 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1670771148
transform -1 0 129720 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1670771148
transform -1 0 134504 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1670771148
transform -1 0 148948 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1236_
timestamp 1670771148
transform -1 0 116840 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1670771148
transform 1 0 122912 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1238_
timestamp 1670771148
transform -1 0 109756 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1239_
timestamp 1670771148
transform -1 0 118864 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1670771148
transform -1 0 109112 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1670771148
transform -1 0 117760 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1670771148
transform 1 0 106996 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1670771148
transform 1 0 119876 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1244_
timestamp 1670771148
transform -1 0 121716 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1670771148
transform 1 0 143704 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1670771148
transform 1 0 145636 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1670771148
transform -1 0 144532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1670771148
transform -1 0 146464 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1670771148
transform -1 0 143336 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1670771148
transform -1 0 143244 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1670771148
transform -1 0 146372 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1670771148
transform -1 0 129076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1670771148
transform 1 0 108376 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1670771148
transform 1 0 117760 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1670771148
transform 1 0 135332 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1670771148
transform 1 0 147476 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1257_
timestamp 1670771148
transform -1 0 142600 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1670771148
transform 1 0 143060 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1259_
timestamp 1670771148
transform -1 0 142048 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1670771148
transform 1 0 145912 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1670771148
transform 1 0 144900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1670771148
transform 1 0 144256 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1670771148
transform 1 0 147476 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1670771148
transform 1 0 145636 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1670771148
transform 1 0 145176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1670771148
transform -1 0 147108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1670771148
transform -1 0 143888 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1670771148
transform -1 0 140576 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1670771148
transform 1 0 131284 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1670771148
transform 1 0 147568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1670771148
transform -1 0 142968 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1670771148
transform 1 0 148212 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1670771148
transform 1 0 147476 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1670771148
transform 1 0 148212 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1670771148
transform 1 0 148212 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1670771148
transform -1 0 147108 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1670771148
transform 1 0 143060 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1670771148
transform 1 0 140944 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1670771148
transform -1 0 147108 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1670771148
transform -1 0 135884 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1670771148
transform 1 0 145636 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1670771148
transform -1 0 148948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1670771148
transform -1 0 148120 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1670771148
transform 1 0 143704 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1670771148
transform 1 0 143612 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1670771148
transform -1 0 147568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1670771148
transform 1 0 120428 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1670771148
transform -1 0 129352 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1670771148
transform -1 0 123924 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1670771148
transform 1 0 148212 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1670771148
transform -1 0 142508 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1670771148
transform -1 0 144808 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1670771148
transform -1 0 147108 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1670771148
transform 1 0 148212 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1295_
timestamp 1670771148
transform -1 0 147660 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1670771148
transform -1 0 146740 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1670771148
transform -1 0 147200 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1298_
timestamp 1670771148
transform -1 0 144900 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1670771148
transform -1 0 145176 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1670771148
transform -1 0 145176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1670771148
transform 1 0 144164 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1670771148
transform -1 0 143336 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1670771148
transform 1 0 148212 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1670771148
transform 1 0 137264 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1670771148
transform -1 0 143244 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1670771148
transform -1 0 139932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1670771148
transform -1 0 137448 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1670771148
transform 1 0 145636 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1670771148
transform -1 0 139932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1670771148
transform -1 0 130916 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1670771148
transform 1 0 105064 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1670771148
transform -1 0 109020 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1670771148
transform 1 0 113712 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1670771148
transform 1 0 111320 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1670771148
transform -1 0 112424 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1670771148
transform 1 0 94760 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1670771148
transform 1 0 107364 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1670771148
transform -1 0 111044 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1319_
timestamp 1670771148
transform 1 0 97060 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1670771148
transform -1 0 102304 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1321_
timestamp 1670771148
transform 1 0 79028 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1322_
timestamp 1670771148
transform 1 0 99268 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1670771148
transform -1 0 25484 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1670771148
transform -1 0 21528 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1670771148
transform -1 0 30820 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1670771148
transform -1 0 21252 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1670771148
transform -1 0 20976 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1670771148
transform -1 0 18216 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1670771148
transform -1 0 15088 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1670771148
transform -1 0 33856 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1670771148
transform -1 0 34408 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1670771148
transform 1 0 30268 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1670771148
transform -1 0 31832 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1670771148
transform -1 0 31832 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1670771148
transform -1 0 29992 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1670771148
transform -1 0 26404 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1670771148
transform -1 0 34316 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1670771148
transform -1 0 28980 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1670771148
transform -1 0 25300 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1670771148
transform 1 0 21344 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1670771148
transform 1 0 29624 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1670771148
transform -1 0 32108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1670771148
transform -1 0 28704 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1670771148
transform -1 0 37444 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1670771148
transform -1 0 44068 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1670771148
transform -1 0 26312 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1670771148
transform -1 0 35420 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1670771148
transform 1 0 38088 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1670771148
transform 1 0 30176 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1670771148
transform 1 0 29992 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1670771148
transform 1 0 20700 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1670771148
transform -1 0 36156 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1670771148
transform -1 0 51060 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1670771148
transform 1 0 35512 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1670771148
transform -1 0 52440 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1670771148
transform -1 0 42136 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1670771148
transform -1 0 46644 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1670771148
transform 1 0 17112 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1670771148
transform 1 0 17388 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1670771148
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1670771148
transform 1 0 17480 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1670771148
transform 1 0 27784 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1670771148
transform 1 0 21620 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1670771148
transform 1 0 24840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1670771148
transform 1 0 31096 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1670771148
transform -1 0 55568 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1670771148
transform -1 0 49864 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1670771148
transform -1 0 36340 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1670771148
transform -1 0 42136 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1670771148
transform -1 0 55384 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1670771148
transform 1 0 31648 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1670771148
transform 1 0 29716 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1670771148
transform 1 0 47840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1670771148
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1670771148
transform 1 0 34132 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1670771148
transform -1 0 44712 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1670771148
transform -1 0 44712 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1670771148
transform -1 0 58880 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1670771148
transform -1 0 42872 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1670771148
transform -1 0 46460 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1670771148
transform 1 0 25208 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1670771148
transform -1 0 46092 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1670771148
transform 1 0 38272 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1670771148
transform -1 0 46644 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1670771148
transform -1 0 50876 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1670771148
transform 1 0 40204 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1670771148
transform 1 0 56120 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1670771148
transform -1 0 47288 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1670771148
transform 1 0 41400 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1670771148
transform -1 0 60904 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1670771148
transform 1 0 27784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1670771148
transform 1 0 31740 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1670771148
transform 1 0 55384 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1670771148
transform -1 0 64676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1670771148
transform -1 0 60812 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1670771148
transform -1 0 55016 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1670771148
transform -1 0 74612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1670771148
transform 1 0 47748 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1670771148
transform 1 0 42504 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1670771148
transform -1 0 52440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1670771148
transform 1 0 48392 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1670771148
transform -1 0 76268 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1670771148
transform -1 0 70380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1670771148
transform -1 0 67712 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1670771148
transform -1 0 52440 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1670771148
transform 1 0 48392 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1670771148
transform 1 0 52900 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1670771148
transform 1 0 45540 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1670771148
transform -1 0 55752 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1670771148
transform 1 0 60628 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1670771148
transform 1 0 53544 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1670771148
transform 1 0 51704 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1670771148
transform 1 0 56120 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1670771148
transform 1 0 52072 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1670771148
transform 1 0 49772 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1670771148
transform 1 0 55476 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1670771148
transform 1 0 52900 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1670771148
transform 1 0 61272 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1670771148
transform 1 0 54004 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1670771148
transform 1 0 61088 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1670771148
transform 1 0 57224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1670771148
transform -1 0 67252 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1670771148
transform -1 0 67252 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1670771148
transform -1 0 65596 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1670771148
transform -1 0 76360 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1670771148
transform 1 0 58696 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1670771148
transform -1 0 77556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1670771148
transform -1 0 69828 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1670771148
transform -1 0 75624 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1670771148
transform -1 0 88228 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1670771148
transform -1 0 93012 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1670771148
transform 1 0 66516 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1670771148
transform -1 0 79212 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1670771148
transform -1 0 92368 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1670771148
transform 1 0 93380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1670771148
transform -1 0 87492 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1670771148
transform -1 0 80500 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1670771148
transform -1 0 82708 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1670771148
transform -1 0 90436 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1670771148
transform -1 0 83904 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1670771148
transform -1 0 85928 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1670771148
transform -1 0 76452 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1670771148
transform 1 0 73968 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1670771148
transform -1 0 90436 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1670771148
transform -1 0 92092 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1670771148
transform -1 0 89240 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1670771148
transform 1 0 73692 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1670771148
transform -1 0 80592 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1670771148
transform -1 0 87676 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1670771148
transform 1 0 70840 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1670771148
transform 1 0 79672 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1670771148
transform 1 0 69828 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1670771148
transform -1 0 85284 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1670771148
transform 1 0 56120 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1670771148
transform -1 0 88504 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1670771148
transform 1 0 68356 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1670771148
transform -1 0 93012 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1670771148
transform -1 0 90436 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1670771148
transform -1 0 93196 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1670771148
transform 1 0 60812 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1670771148
transform -1 0 86848 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1670771148
transform 1 0 71852 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1670771148
transform 1 0 69644 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1670771148
transform 1 0 59248 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1670771148
transform -1 0 90436 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1670771148
transform 1 0 61272 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1670771148
transform 1 0 81052 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1670771148
transform 1 0 86388 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1670771148
transform 1 0 60996 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1670771148
transform 1 0 65596 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1670771148
transform -1 0 111044 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1670771148
transform 1 0 69184 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1670771148
transform 1 0 58052 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1670771148
transform 1 0 58052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1670771148
transform -1 0 98164 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1476_
timestamp 1670771148
transform -1 0 142048 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1477_
timestamp 1670771148
transform -1 0 150696 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1478_
timestamp 1670771148
transform -1 0 154928 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1479_
timestamp 1670771148
transform -1 0 144624 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1670771148
transform -1 0 107088 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1670771148
transform 1 0 95404 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1670771148
transform 1 0 91172 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1670771148
transform 1 0 76728 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1670771148
transform 1 0 91540 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1485_
timestamp 1670771148
transform -1 0 123924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1486_
timestamp 1670771148
transform 1 0 98348 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1670771148
transform -1 0 124936 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1488_
timestamp 1670771148
transform -1 0 151432 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1489_
timestamp 1670771148
transform -1 0 119416 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1490_
timestamp 1670771148
transform -1 0 123188 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1491_
timestamp 1670771148
transform -1 0 121348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1492_
timestamp 1670771148
transform 1 0 89516 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1670771148
transform -1 0 125488 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1670771148
transform 1 0 81144 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1670771148
transform 1 0 91264 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1670771148
transform -1 0 103316 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1670771148
transform -1 0 123280 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1670771148
transform -1 0 109756 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1670771148
transform -1 0 117760 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1670771148
transform -1 0 116840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1501_
timestamp 1670771148
transform 1 0 154468 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1502_
timestamp 1670771148
transform -1 0 155296 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1503_
timestamp 1670771148
transform -1 0 129812 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1504_
timestamp 1670771148
transform -1 0 152352 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1505_
timestamp 1670771148
transform -1 0 151892 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1506_
timestamp 1670771148
transform -1 0 150236 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1507_
timestamp 1670771148
transform 1 0 109112 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1508_
timestamp 1670771148
transform 1 0 127604 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1670771148
transform -1 0 119232 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1670771148
transform -1 0 121072 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1670771148
transform -1 0 131652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1670771148
transform -1 0 116196 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1513_
timestamp 1670771148
transform 1 0 109572 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1670771148
transform -1 0 152260 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1670771148
transform 1 0 107640 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1670771148
transform -1 0 154100 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1670771148
transform -1 0 154100 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1670771148
transform -1 0 152260 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1670771148
transform -1 0 154100 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1670771148
transform -1 0 149960 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1670771148
transform -1 0 151524 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1670771148
transform -1 0 136804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1670771148
transform -1 0 133492 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1670771148
transform -1 0 133032 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1670771148
transform -1 0 147108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1670771148
transform -1 0 152260 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1670771148
transform -1 0 155204 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1670771148
transform -1 0 154836 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1670771148
transform -1 0 152260 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1670771148
transform -1 0 152536 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1670771148
transform -1 0 144532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1670771148
transform -1 0 129076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1670771148
transform -1 0 149684 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1670771148
transform -1 0 144900 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1670771148
transform -1 0 145084 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1670771148
transform 1 0 126040 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1670771148
transform -1 0 152720 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1670771148
transform -1 0 142324 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1670771148
transform -1 0 142232 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1670771148
transform -1 0 149684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1670771148
transform -1 0 154744 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1670771148
transform -1 0 136896 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1543_
timestamp 1670771148
transform -1 0 134872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1670771148
transform 1 0 124108 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1670771148
transform 1 0 122452 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1670771148
transform 1 0 122176 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1547_
timestamp 1670771148
transform 1 0 123004 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1548_
timestamp 1670771148
transform 1 0 117300 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1670771148
transform 1 0 118956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1550_
timestamp 1670771148
transform 1 0 126868 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1551_
timestamp 1670771148
transform 1 0 104604 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1552_
timestamp 1670771148
transform 1 0 125488 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1670771148
transform 1 0 121808 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1554_
timestamp 1670771148
transform -1 0 115000 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1555_
timestamp 1670771148
transform 1 0 135976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1556_
timestamp 1670771148
transform 1 0 114724 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1557_
timestamp 1670771148
transform 1 0 138000 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1670771148
transform 1 0 125120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1670771148
transform -1 0 151524 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1670771148
transform -1 0 122452 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1670771148
transform 1 0 133216 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1562_
timestamp 1670771148
transform 1 0 116564 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1670771148
transform 1 0 134136 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1670771148
transform -1 0 152260 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1565_
timestamp 1670771148
transform -1 0 154836 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1670771148
transform 1 0 131192 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1670771148
transform 1 0 133676 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1670771148
transform 1 0 103776 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1670771148
transform 1 0 121716 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1670771148
transform 1 0 148488 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1670771148
transform 1 0 133124 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1670771148
transform 1 0 137908 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1670771148
transform 1 0 129168 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1670771148
transform -1 0 130548 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1670771148
transform 1 0 150788 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1576_
timestamp 1670771148
transform 1 0 105064 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1670771148
transform 1 0 133400 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1670771148
transform 1 0 138552 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1670771148
transform 1 0 25944 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1670771148
transform 1 0 11776 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1670771148
transform 1 0 16192 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1670771148
transform 1 0 19412 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1670771148
transform 1 0 14628 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1670771148
transform 1 0 14444 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1670771148
transform -1 0 13800 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1670771148
transform 1 0 14260 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1670771148
transform 1 0 20056 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1670771148
transform 1 0 22540 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1670771148
transform 1 0 18492 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1670771148
transform 1 0 15088 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1670771148
transform -1 0 19320 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_sclk pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 81236 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_sclk
timestamp 1670771148
transform -1 0 77280 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_sclk
timestamp 1670771148
transform 1 0 81236 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_sclk
timestamp 1670771148
transform 1 0 34500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_sclk
timestamp 1670771148
transform -1 0 21252 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_sclk
timestamp 1670771148
transform -1 0 69368 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_sclk
timestamp 1670771148
transform -1 0 112608 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_sclk
timestamp 1670771148
transform 1 0 141772 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_sclk
timestamp 1670771148
transform 1 0 119416 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_sclk
timestamp 1670771148
transform 1 0 141220 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_sclk
timestamp 1670771148
transform 1 0 131560 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_sclk
timestamp 1670771148
transform 1 0 76728 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_sclk
timestamp 1670771148
transform 1 0 24564 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_sclk
timestamp 1670771148
transform 1 0 64216 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout261
timestamp 1670771148
transform -1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout262
timestamp 1670771148
transform -1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout263
timestamp 1670771148
transform 1 0 25024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout264
timestamp 1670771148
transform 1 0 31464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout265
timestamp 1670771148
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout266
timestamp 1670771148
transform 1 0 41768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout267
timestamp 1670771148
transform 1 0 41768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout268
timestamp 1670771148
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout269
timestamp 1670771148
transform -1 0 48760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout270
timestamp 1670771148
transform 1 0 52900 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout271
timestamp 1670771148
transform 1 0 47656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout272
timestamp 1670771148
transform 1 0 54648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout273
timestamp 1670771148
transform 1 0 57592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout274
timestamp 1670771148
transform -1 0 66884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout275
timestamp 1670771148
transform 1 0 74888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout276
timestamp 1670771148
transform 1 0 68080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout277
timestamp 1670771148
transform 1 0 49036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout278
timestamp 1670771148
transform 1 0 88964 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout279
timestamp 1670771148
transform 1 0 85376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout280
timestamp 1670771148
transform 1 0 84640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout281
timestamp 1670771148
transform -1 0 115828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout282
timestamp 1670771148
transform 1 0 103316 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout283
timestamp 1670771148
transform 1 0 121532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout284
timestamp 1670771148
transform -1 0 122176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout285
timestamp 1670771148
transform 1 0 128524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout286
timestamp 1670771148
transform 1 0 130456 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout287
timestamp 1670771148
transform 1 0 137908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout288
timestamp 1670771148
transform 1 0 150052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout289
timestamp 1670771148
transform 1 0 149316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout290
timestamp 1670771148
transform 1 0 149316 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout291
timestamp 1670771148
transform 1 0 138000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout292
timestamp 1670771148
transform 1 0 85376 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1670771148
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1670771148
transform 1 0 1564 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1670771148
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1670771148
transform -1 0 8648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1670771148
transform -1 0 65228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1670771148
transform 1 0 65228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1670771148
transform -1 0 66332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1670771148
transform 1 0 65780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1670771148
transform 1 0 66792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1670771148
transform -1 0 67896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1670771148
transform -1 0 67896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1670771148
transform -1 0 69092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1670771148
transform 1 0 68632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1670771148
transform 1 0 69828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1670771148
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1670771148
transform -1 0 69736 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1670771148
transform -1 0 70472 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1670771148
transform -1 0 71576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1670771148
transform -1 0 72312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1670771148
transform -1 0 73048 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1670771148
transform -1 0 73048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1670771148
transform -1 0 74888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1670771148
transform -1 0 74152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1670771148
transform -1 0 74888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1670771148
transform 1 0 75348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1670771148
transform -1 0 13800 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1670771148
transform 1 0 75256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1670771148
transform -1 0 76820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1670771148
transform -1 0 76452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1670771148
transform -1 0 77924 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1670771148
transform 1 0 77832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1670771148
transform -1 0 79028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1670771148
transform -1 0 79212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1670771148
transform 1 0 79580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1670771148
transform -1 0 80684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1670771148
transform 1 0 81236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1670771148
transform 1 0 14812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1670771148
transform -1 0 82340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1670771148
transform -1 0 83076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1670771148
transform -1 0 83260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1670771148
transform -1 0 84180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1670771148
transform -1 0 84180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1670771148
transform -1 0 84916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1670771148
transform -1 0 85652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1670771148
transform -1 0 85652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1670771148
transform 1 0 86388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1670771148
transform 1 0 87860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1670771148
transform -1 0 16376 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1670771148
transform 1 0 87216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1670771148
transform -1 0 89332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1670771148
transform 1 0 89700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1670771148
transform -1 0 90896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1670771148
transform 1 0 89608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1670771148
transform 1 0 90344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1670771148
transform -1 0 93472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1670771148
transform -1 0 94484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1670771148
transform -1 0 95220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1670771148
transform -1 0 93748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1670771148
transform -1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1670771148
transform -1 0 94484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1670771148
transform -1 0 95956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1670771148
transform -1 0 94484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1670771148
transform -1 0 97060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1670771148
transform -1 0 95220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1670771148
transform -1 0 97796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1670771148
transform -1 0 97612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1670771148
transform -1 0 97060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1670771148
transform 1 0 98164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1670771148
transform 1 0 97980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1670771148
transform -1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1670771148
transform -1 0 99636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1670771148
transform 1 0 100004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1670771148
transform -1 0 101108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1670771148
transform 1 0 100096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1670771148
transform -1 0 101200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1670771148
transform -1 0 101936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1670771148
transform -1 0 103408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1670771148
transform -1 0 102672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1670771148
transform -1 0 103408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1670771148
transform -1 0 104788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1670771148
transform -1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1670771148
transform -1 0 105524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1670771148
transform -1 0 104788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1670771148
transform 1 0 105892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1670771148
transform 1 0 105156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1670771148
transform -1 0 106260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1670771148
transform -1 0 107824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1670771148
transform -1 0 107364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1670771148
transform -1 0 108560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1670771148
transform -1 0 109940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1670771148
transform -1 0 109940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1670771148
transform -1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1670771148
transform -1 0 110676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1670771148
transform -1 0 111412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1670771148
transform -1 0 110492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1670771148
transform -1 0 112516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1670771148
transform 1 0 112884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1670771148
transform -1 0 112516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1670771148
transform -1 0 113160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1670771148
transform -1 0 113988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1670771148
transform -1 0 113896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1670771148
transform 1 0 114724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1670771148
transform -1 0 18952 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1670771148
transform 1 0 116196 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1670771148
transform -1 0 115460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1670771148
transform 1 0 117300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1670771148
transform -1 0 116564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1670771148
transform -1 0 118404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1670771148
transform -1 0 119140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1670771148
transform -1 0 118772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1670771148
transform -1 0 120244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1670771148
transform -1 0 120980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1670771148
transform -1 0 120244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1670771148
transform -1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1670771148
transform -1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1670771148
transform -1 0 120980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1670771148
transform -1 0 121716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1670771148
transform -1 0 121716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1670771148
transform -1 0 121992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1670771148
transform -1 0 124384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1670771148
transform -1 0 125396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1670771148
transform -1 0 125396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1670771148
transform -1 0 124660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1670771148
transform -1 0 126132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1670771148
transform -1 0 126132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1670771148
transform -1 0 21068 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1670771148
transform -1 0 126868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1670771148
transform -1 0 127972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1670771148
transform -1 0 128708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1670771148
transform 1 0 127604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1670771148
transform -1 0 129444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1670771148
transform -1 0 129076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1670771148
transform -1 0 130548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1670771148
transform -1 0 130548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1670771148
transform -1 0 131284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1670771148
transform -1 0 131284 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1670771148
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1670771148
transform -1 0 132020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1670771148
transform 1 0 131652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1670771148
transform 1 0 132756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1670771148
transform 1 0 133492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1670771148
transform 1 0 134228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1670771148
transform -1 0 134412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1670771148
transform -1 0 135700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1670771148
transform 1 0 135332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1670771148
transform 1 0 136068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1670771148
transform 1 0 136804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1670771148
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1670771148
transform 1 0 136620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1670771148
transform -1 0 138276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1670771148
transform 1 0 137724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1670771148
transform -1 0 139012 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1670771148
transform 1 0 139380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1670771148
transform 1 0 139380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1670771148
transform -1 0 140852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1670771148
transform 1 0 141220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1670771148
transform 1 0 141956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1670771148
transform 1 0 141128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1670771148
transform -1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1670771148
transform 1 0 142692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1670771148
transform -1 0 139012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1670771148
transform -1 0 147200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1670771148
transform -1 0 148580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1670771148
transform -1 0 149684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1670771148
transform 1 0 148948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1670771148
transform 1 0 153364 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1670771148
transform 1 0 154100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1670771148
transform 1 0 154836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1670771148
transform 1 0 155940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1670771148
transform -1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1670771148
transform 1 0 156676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1670771148
transform 1 0 155940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1670771148
transform 1 0 156032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1670771148
transform 1 0 157412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1670771148
transform 1 0 156676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1670771148
transform 1 0 156768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1670771148
transform -1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1670771148
transform -1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1670771148
transform -1 0 24104 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1670771148
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1670771148
transform -1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1670771148
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1670771148
transform 1 0 23736 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1670771148
transform -1 0 26680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1670771148
transform -1 0 27508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1670771148
transform -1 0 28244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1670771148
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1670771148
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1670771148
transform 1 0 29716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1670771148
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1670771148
transform 1 0 28888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1670771148
transform 1 0 31464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1670771148
transform 1 0 9384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1670771148
transform 1 0 32476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1670771148
transform 1 0 32292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1670771148
transform 1 0 32568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1670771148
transform -1 0 33764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1670771148
transform -1 0 34316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1670771148
transform -1 0 33672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1670771148
transform -1 0 35420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1670771148
transform -1 0 34408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1670771148
transform 1 0 36156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1670771148
transform 1 0 36616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1670771148
transform -1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1670771148
transform -1 0 37628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1670771148
transform 1 0 37720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1670771148
transform 1 0 38364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1670771148
transform -1 0 38824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1670771148
transform -1 0 38088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1670771148
transform 1 0 39192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1670771148
transform -1 0 40940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1670771148
transform -1 0 38824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1670771148
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1670771148
transform -1 0 40296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1670771148
transform -1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1670771148
transform -1 0 39560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1670771148
transform -1 0 42136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1670771148
transform -1 0 42872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1670771148
transform 1 0 42688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1670771148
transform -1 0 45356 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1670771148
transform -1 0 41308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1670771148
transform 1 0 43424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1670771148
transform -1 0 46368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1670771148
transform 1 0 43608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1670771148
transform 1 0 44160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1670771148
transform -1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1670771148
transform 1 0 44896 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1670771148
transform 1 0 44344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1670771148
transform -1 0 45540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1670771148
transform -1 0 45172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1670771148
transform -1 0 50692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1670771148
transform -1 0 48668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1670771148
transform 1 0 51060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1670771148
transform -1 0 49404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1670771148
transform 1 0 50876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1670771148
transform -1 0 53636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1670771148
transform 1 0 10856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1670771148
transform 1 0 50600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1670771148
transform -1 0 50600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1670771148
transform -1 0 51704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1670771148
transform 1 0 53544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1670771148
transform 1 0 56028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1670771148
transform 1 0 56580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1670771148
transform -1 0 54280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1670771148
transform -1 0 53636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1670771148
transform 1 0 58236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1670771148
transform 1 0 58788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1670771148
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1670771148
transform 1 0 57684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1670771148
transform 1 0 59800 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1670771148
transform 1 0 63940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1670771148
transform 1 0 59800 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1670771148
transform 1 0 58696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1670771148
transform -1 0 62836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1670771148
transform 1 0 63204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1670771148
transform 1 0 63020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1670771148
transform 1 0 63756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1670771148
transform -1 0 64124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1670771148
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1670771148
transform 1 0 158056 0 -1 8704
box -38 -48 406 592
<< labels >>
flabel metal2 s 9586 15200 9642 16000 0 FreeSans 224 90 0 0 dq[0]
port 0 nsew signal tristate
flabel metal2 s 64786 15200 64842 16000 0 FreeSans 224 90 0 0 dq[100]
port 1 nsew signal tristate
flabel metal2 s 65338 15200 65394 16000 0 FreeSans 224 90 0 0 dq[101]
port 2 nsew signal tristate
flabel metal2 s 65890 15200 65946 16000 0 FreeSans 224 90 0 0 dq[102]
port 3 nsew signal tristate
flabel metal2 s 66442 15200 66498 16000 0 FreeSans 224 90 0 0 dq[103]
port 4 nsew signal tristate
flabel metal2 s 66994 15200 67050 16000 0 FreeSans 224 90 0 0 dq[104]
port 5 nsew signal tristate
flabel metal2 s 67546 15200 67602 16000 0 FreeSans 224 90 0 0 dq[105]
port 6 nsew signal tristate
flabel metal2 s 68098 15200 68154 16000 0 FreeSans 224 90 0 0 dq[106]
port 7 nsew signal tristate
flabel metal2 s 68650 15200 68706 16000 0 FreeSans 224 90 0 0 dq[107]
port 8 nsew signal tristate
flabel metal2 s 69202 15200 69258 16000 0 FreeSans 224 90 0 0 dq[108]
port 9 nsew signal tristate
flabel metal2 s 69754 15200 69810 16000 0 FreeSans 224 90 0 0 dq[109]
port 10 nsew signal tristate
flabel metal2 s 15106 15200 15162 16000 0 FreeSans 224 90 0 0 dq[10]
port 11 nsew signal tristate
flabel metal2 s 70306 15200 70362 16000 0 FreeSans 224 90 0 0 dq[110]
port 12 nsew signal tristate
flabel metal2 s 70858 15200 70914 16000 0 FreeSans 224 90 0 0 dq[111]
port 13 nsew signal tristate
flabel metal2 s 71410 15200 71466 16000 0 FreeSans 224 90 0 0 dq[112]
port 14 nsew signal tristate
flabel metal2 s 71962 15200 72018 16000 0 FreeSans 224 90 0 0 dq[113]
port 15 nsew signal tristate
flabel metal2 s 72514 15200 72570 16000 0 FreeSans 224 90 0 0 dq[114]
port 16 nsew signal tristate
flabel metal2 s 73066 15200 73122 16000 0 FreeSans 224 90 0 0 dq[115]
port 17 nsew signal tristate
flabel metal2 s 73618 15200 73674 16000 0 FreeSans 224 90 0 0 dq[116]
port 18 nsew signal tristate
flabel metal2 s 74170 15200 74226 16000 0 FreeSans 224 90 0 0 dq[117]
port 19 nsew signal tristate
flabel metal2 s 74722 15200 74778 16000 0 FreeSans 224 90 0 0 dq[118]
port 20 nsew signal tristate
flabel metal2 s 75274 15200 75330 16000 0 FreeSans 224 90 0 0 dq[119]
port 21 nsew signal tristate
flabel metal2 s 15658 15200 15714 16000 0 FreeSans 224 90 0 0 dq[11]
port 22 nsew signal tristate
flabel metal2 s 75826 15200 75882 16000 0 FreeSans 224 90 0 0 dq[120]
port 23 nsew signal tristate
flabel metal2 s 76378 15200 76434 16000 0 FreeSans 224 90 0 0 dq[121]
port 24 nsew signal tristate
flabel metal2 s 76930 15200 76986 16000 0 FreeSans 224 90 0 0 dq[122]
port 25 nsew signal tristate
flabel metal2 s 77482 15200 77538 16000 0 FreeSans 224 90 0 0 dq[123]
port 26 nsew signal tristate
flabel metal2 s 78034 15200 78090 16000 0 FreeSans 224 90 0 0 dq[124]
port 27 nsew signal tristate
flabel metal2 s 78586 15200 78642 16000 0 FreeSans 224 90 0 0 dq[125]
port 28 nsew signal tristate
flabel metal2 s 79138 15200 79194 16000 0 FreeSans 224 90 0 0 dq[126]
port 29 nsew signal tristate
flabel metal2 s 79690 15200 79746 16000 0 FreeSans 224 90 0 0 dq[127]
port 30 nsew signal tristate
flabel metal2 s 80242 15200 80298 16000 0 FreeSans 224 90 0 0 dq[128]
port 31 nsew signal tristate
flabel metal2 s 80794 15200 80850 16000 0 FreeSans 224 90 0 0 dq[129]
port 32 nsew signal tristate
flabel metal2 s 16210 15200 16266 16000 0 FreeSans 224 90 0 0 dq[12]
port 33 nsew signal tristate
flabel metal2 s 81346 15200 81402 16000 0 FreeSans 224 90 0 0 dq[130]
port 34 nsew signal tristate
flabel metal2 s 81898 15200 81954 16000 0 FreeSans 224 90 0 0 dq[131]
port 35 nsew signal tristate
flabel metal2 s 82450 15200 82506 16000 0 FreeSans 224 90 0 0 dq[132]
port 36 nsew signal tristate
flabel metal2 s 83002 15200 83058 16000 0 FreeSans 224 90 0 0 dq[133]
port 37 nsew signal tristate
flabel metal2 s 83554 15200 83610 16000 0 FreeSans 224 90 0 0 dq[134]
port 38 nsew signal tristate
flabel metal2 s 84106 15200 84162 16000 0 FreeSans 224 90 0 0 dq[135]
port 39 nsew signal tristate
flabel metal2 s 84658 15200 84714 16000 0 FreeSans 224 90 0 0 dq[136]
port 40 nsew signal tristate
flabel metal2 s 85210 15200 85266 16000 0 FreeSans 224 90 0 0 dq[137]
port 41 nsew signal tristate
flabel metal2 s 85762 15200 85818 16000 0 FreeSans 224 90 0 0 dq[138]
port 42 nsew signal tristate
flabel metal2 s 86314 15200 86370 16000 0 FreeSans 224 90 0 0 dq[139]
port 43 nsew signal tristate
flabel metal2 s 16762 15200 16818 16000 0 FreeSans 224 90 0 0 dq[13]
port 44 nsew signal tristate
flabel metal2 s 86866 15200 86922 16000 0 FreeSans 224 90 0 0 dq[140]
port 45 nsew signal tristate
flabel metal2 s 87418 15200 87474 16000 0 FreeSans 224 90 0 0 dq[141]
port 46 nsew signal tristate
flabel metal2 s 87970 15200 88026 16000 0 FreeSans 224 90 0 0 dq[142]
port 47 nsew signal tristate
flabel metal2 s 88522 15200 88578 16000 0 FreeSans 224 90 0 0 dq[143]
port 48 nsew signal tristate
flabel metal2 s 89074 15200 89130 16000 0 FreeSans 224 90 0 0 dq[144]
port 49 nsew signal tristate
flabel metal2 s 89626 15200 89682 16000 0 FreeSans 224 90 0 0 dq[145]
port 50 nsew signal tristate
flabel metal2 s 90178 15200 90234 16000 0 FreeSans 224 90 0 0 dq[146]
port 51 nsew signal tristate
flabel metal2 s 90730 15200 90786 16000 0 FreeSans 224 90 0 0 dq[147]
port 52 nsew signal tristate
flabel metal2 s 91282 15200 91338 16000 0 FreeSans 224 90 0 0 dq[148]
port 53 nsew signal tristate
flabel metal2 s 91834 15200 91890 16000 0 FreeSans 224 90 0 0 dq[149]
port 54 nsew signal tristate
flabel metal2 s 17314 15200 17370 16000 0 FreeSans 224 90 0 0 dq[14]
port 55 nsew signal tristate
flabel metal2 s 92386 15200 92442 16000 0 FreeSans 224 90 0 0 dq[150]
port 56 nsew signal tristate
flabel metal2 s 92938 15200 92994 16000 0 FreeSans 224 90 0 0 dq[151]
port 57 nsew signal tristate
flabel metal2 s 93490 15200 93546 16000 0 FreeSans 224 90 0 0 dq[152]
port 58 nsew signal tristate
flabel metal2 s 94042 15200 94098 16000 0 FreeSans 224 90 0 0 dq[153]
port 59 nsew signal tristate
flabel metal2 s 94594 15200 94650 16000 0 FreeSans 224 90 0 0 dq[154]
port 60 nsew signal tristate
flabel metal2 s 95146 15200 95202 16000 0 FreeSans 224 90 0 0 dq[155]
port 61 nsew signal tristate
flabel metal2 s 95698 15200 95754 16000 0 FreeSans 224 90 0 0 dq[156]
port 62 nsew signal tristate
flabel metal2 s 96250 15200 96306 16000 0 FreeSans 224 90 0 0 dq[157]
port 63 nsew signal tristate
flabel metal2 s 96802 15200 96858 16000 0 FreeSans 224 90 0 0 dq[158]
port 64 nsew signal tristate
flabel metal2 s 97354 15200 97410 16000 0 FreeSans 224 90 0 0 dq[159]
port 65 nsew signal tristate
flabel metal2 s 17866 15200 17922 16000 0 FreeSans 224 90 0 0 dq[15]
port 66 nsew signal tristate
flabel metal2 s 97906 15200 97962 16000 0 FreeSans 224 90 0 0 dq[160]
port 67 nsew signal tristate
flabel metal2 s 98458 15200 98514 16000 0 FreeSans 224 90 0 0 dq[161]
port 68 nsew signal tristate
flabel metal2 s 99010 15200 99066 16000 0 FreeSans 224 90 0 0 dq[162]
port 69 nsew signal tristate
flabel metal2 s 99562 15200 99618 16000 0 FreeSans 224 90 0 0 dq[163]
port 70 nsew signal tristate
flabel metal2 s 100114 15200 100170 16000 0 FreeSans 224 90 0 0 dq[164]
port 71 nsew signal tristate
flabel metal2 s 100666 15200 100722 16000 0 FreeSans 224 90 0 0 dq[165]
port 72 nsew signal tristate
flabel metal2 s 101218 15200 101274 16000 0 FreeSans 224 90 0 0 dq[166]
port 73 nsew signal tristate
flabel metal2 s 101770 15200 101826 16000 0 FreeSans 224 90 0 0 dq[167]
port 74 nsew signal tristate
flabel metal2 s 102322 15200 102378 16000 0 FreeSans 224 90 0 0 dq[168]
port 75 nsew signal tristate
flabel metal2 s 102874 15200 102930 16000 0 FreeSans 224 90 0 0 dq[169]
port 76 nsew signal tristate
flabel metal2 s 18418 15200 18474 16000 0 FreeSans 224 90 0 0 dq[16]
port 77 nsew signal tristate
flabel metal2 s 103426 15200 103482 16000 0 FreeSans 224 90 0 0 dq[170]
port 78 nsew signal tristate
flabel metal2 s 103978 15200 104034 16000 0 FreeSans 224 90 0 0 dq[171]
port 79 nsew signal tristate
flabel metal2 s 104530 15200 104586 16000 0 FreeSans 224 90 0 0 dq[172]
port 80 nsew signal tristate
flabel metal2 s 105082 15200 105138 16000 0 FreeSans 224 90 0 0 dq[173]
port 81 nsew signal tristate
flabel metal2 s 105634 15200 105690 16000 0 FreeSans 224 90 0 0 dq[174]
port 82 nsew signal tristate
flabel metal2 s 106186 15200 106242 16000 0 FreeSans 224 90 0 0 dq[175]
port 83 nsew signal tristate
flabel metal2 s 106738 15200 106794 16000 0 FreeSans 224 90 0 0 dq[176]
port 84 nsew signal tristate
flabel metal2 s 107290 15200 107346 16000 0 FreeSans 224 90 0 0 dq[177]
port 85 nsew signal tristate
flabel metal2 s 107842 15200 107898 16000 0 FreeSans 224 90 0 0 dq[178]
port 86 nsew signal tristate
flabel metal2 s 108394 15200 108450 16000 0 FreeSans 224 90 0 0 dq[179]
port 87 nsew signal tristate
flabel metal2 s 18970 15200 19026 16000 0 FreeSans 224 90 0 0 dq[17]
port 88 nsew signal tristate
flabel metal2 s 108946 15200 109002 16000 0 FreeSans 224 90 0 0 dq[180]
port 89 nsew signal tristate
flabel metal2 s 109498 15200 109554 16000 0 FreeSans 224 90 0 0 dq[181]
port 90 nsew signal tristate
flabel metal2 s 110050 15200 110106 16000 0 FreeSans 224 90 0 0 dq[182]
port 91 nsew signal tristate
flabel metal2 s 110602 15200 110658 16000 0 FreeSans 224 90 0 0 dq[183]
port 92 nsew signal tristate
flabel metal2 s 111154 15200 111210 16000 0 FreeSans 224 90 0 0 dq[184]
port 93 nsew signal tristate
flabel metal2 s 111706 15200 111762 16000 0 FreeSans 224 90 0 0 dq[185]
port 94 nsew signal tristate
flabel metal2 s 112258 15200 112314 16000 0 FreeSans 224 90 0 0 dq[186]
port 95 nsew signal tristate
flabel metal2 s 112810 15200 112866 16000 0 FreeSans 224 90 0 0 dq[187]
port 96 nsew signal tristate
flabel metal2 s 113362 15200 113418 16000 0 FreeSans 224 90 0 0 dq[188]
port 97 nsew signal tristate
flabel metal2 s 113914 15200 113970 16000 0 FreeSans 224 90 0 0 dq[189]
port 98 nsew signal tristate
flabel metal2 s 19522 15200 19578 16000 0 FreeSans 224 90 0 0 dq[18]
port 99 nsew signal tristate
flabel metal2 s 114466 15200 114522 16000 0 FreeSans 224 90 0 0 dq[190]
port 100 nsew signal tristate
flabel metal2 s 115018 15200 115074 16000 0 FreeSans 224 90 0 0 dq[191]
port 101 nsew signal tristate
flabel metal2 s 115570 15200 115626 16000 0 FreeSans 224 90 0 0 dq[192]
port 102 nsew signal tristate
flabel metal2 s 116122 15200 116178 16000 0 FreeSans 224 90 0 0 dq[193]
port 103 nsew signal tristate
flabel metal2 s 116674 15200 116730 16000 0 FreeSans 224 90 0 0 dq[194]
port 104 nsew signal tristate
flabel metal2 s 117226 15200 117282 16000 0 FreeSans 224 90 0 0 dq[195]
port 105 nsew signal tristate
flabel metal2 s 117778 15200 117834 16000 0 FreeSans 224 90 0 0 dq[196]
port 106 nsew signal tristate
flabel metal2 s 118330 15200 118386 16000 0 FreeSans 224 90 0 0 dq[197]
port 107 nsew signal tristate
flabel metal2 s 118882 15200 118938 16000 0 FreeSans 224 90 0 0 dq[198]
port 108 nsew signal tristate
flabel metal2 s 119434 15200 119490 16000 0 FreeSans 224 90 0 0 dq[199]
port 109 nsew signal tristate
flabel metal2 s 20074 15200 20130 16000 0 FreeSans 224 90 0 0 dq[19]
port 110 nsew signal tristate
flabel metal2 s 10138 15200 10194 16000 0 FreeSans 224 90 0 0 dq[1]
port 111 nsew signal tristate
flabel metal2 s 119986 15200 120042 16000 0 FreeSans 224 90 0 0 dq[200]
port 112 nsew signal tristate
flabel metal2 s 120538 15200 120594 16000 0 FreeSans 224 90 0 0 dq[201]
port 113 nsew signal tristate
flabel metal2 s 121090 15200 121146 16000 0 FreeSans 224 90 0 0 dq[202]
port 114 nsew signal tristate
flabel metal2 s 121642 15200 121698 16000 0 FreeSans 224 90 0 0 dq[203]
port 115 nsew signal tristate
flabel metal2 s 122194 15200 122250 16000 0 FreeSans 224 90 0 0 dq[204]
port 116 nsew signal tristate
flabel metal2 s 122746 15200 122802 16000 0 FreeSans 224 90 0 0 dq[205]
port 117 nsew signal tristate
flabel metal2 s 123298 15200 123354 16000 0 FreeSans 224 90 0 0 dq[206]
port 118 nsew signal tristate
flabel metal2 s 123850 15200 123906 16000 0 FreeSans 224 90 0 0 dq[207]
port 119 nsew signal tristate
flabel metal2 s 124402 15200 124458 16000 0 FreeSans 224 90 0 0 dq[208]
port 120 nsew signal tristate
flabel metal2 s 124954 15200 125010 16000 0 FreeSans 224 90 0 0 dq[209]
port 121 nsew signal tristate
flabel metal2 s 20626 15200 20682 16000 0 FreeSans 224 90 0 0 dq[20]
port 122 nsew signal tristate
flabel metal2 s 125506 15200 125562 16000 0 FreeSans 224 90 0 0 dq[210]
port 123 nsew signal tristate
flabel metal2 s 126058 15200 126114 16000 0 FreeSans 224 90 0 0 dq[211]
port 124 nsew signal tristate
flabel metal2 s 126610 15200 126666 16000 0 FreeSans 224 90 0 0 dq[212]
port 125 nsew signal tristate
flabel metal2 s 127162 15200 127218 16000 0 FreeSans 224 90 0 0 dq[213]
port 126 nsew signal tristate
flabel metal2 s 127714 15200 127770 16000 0 FreeSans 224 90 0 0 dq[214]
port 127 nsew signal tristate
flabel metal2 s 128266 15200 128322 16000 0 FreeSans 224 90 0 0 dq[215]
port 128 nsew signal tristate
flabel metal2 s 128818 15200 128874 16000 0 FreeSans 224 90 0 0 dq[216]
port 129 nsew signal tristate
flabel metal2 s 129370 15200 129426 16000 0 FreeSans 224 90 0 0 dq[217]
port 130 nsew signal tristate
flabel metal2 s 129922 15200 129978 16000 0 FreeSans 224 90 0 0 dq[218]
port 131 nsew signal tristate
flabel metal2 s 130474 15200 130530 16000 0 FreeSans 224 90 0 0 dq[219]
port 132 nsew signal tristate
flabel metal2 s 21178 15200 21234 16000 0 FreeSans 224 90 0 0 dq[21]
port 133 nsew signal tristate
flabel metal2 s 131026 15200 131082 16000 0 FreeSans 224 90 0 0 dq[220]
port 134 nsew signal tristate
flabel metal2 s 131578 15200 131634 16000 0 FreeSans 224 90 0 0 dq[221]
port 135 nsew signal tristate
flabel metal2 s 132130 15200 132186 16000 0 FreeSans 224 90 0 0 dq[222]
port 136 nsew signal tristate
flabel metal2 s 132682 15200 132738 16000 0 FreeSans 224 90 0 0 dq[223]
port 137 nsew signal tristate
flabel metal2 s 133234 15200 133290 16000 0 FreeSans 224 90 0 0 dq[224]
port 138 nsew signal tristate
flabel metal2 s 133786 15200 133842 16000 0 FreeSans 224 90 0 0 dq[225]
port 139 nsew signal tristate
flabel metal2 s 134338 15200 134394 16000 0 FreeSans 224 90 0 0 dq[226]
port 140 nsew signal tristate
flabel metal2 s 134890 15200 134946 16000 0 FreeSans 224 90 0 0 dq[227]
port 141 nsew signal tristate
flabel metal2 s 135442 15200 135498 16000 0 FreeSans 224 90 0 0 dq[228]
port 142 nsew signal tristate
flabel metal2 s 135994 15200 136050 16000 0 FreeSans 224 90 0 0 dq[229]
port 143 nsew signal tristate
flabel metal2 s 21730 15200 21786 16000 0 FreeSans 224 90 0 0 dq[22]
port 144 nsew signal tristate
flabel metal2 s 136546 15200 136602 16000 0 FreeSans 224 90 0 0 dq[230]
port 145 nsew signal tristate
flabel metal2 s 137098 15200 137154 16000 0 FreeSans 224 90 0 0 dq[231]
port 146 nsew signal tristate
flabel metal2 s 137650 15200 137706 16000 0 FreeSans 224 90 0 0 dq[232]
port 147 nsew signal tristate
flabel metal2 s 138202 15200 138258 16000 0 FreeSans 224 90 0 0 dq[233]
port 148 nsew signal tristate
flabel metal2 s 138754 15200 138810 16000 0 FreeSans 224 90 0 0 dq[234]
port 149 nsew signal tristate
flabel metal2 s 139306 15200 139362 16000 0 FreeSans 224 90 0 0 dq[235]
port 150 nsew signal tristate
flabel metal2 s 139858 15200 139914 16000 0 FreeSans 224 90 0 0 dq[236]
port 151 nsew signal tristate
flabel metal2 s 140410 15200 140466 16000 0 FreeSans 224 90 0 0 dq[237]
port 152 nsew signal tristate
flabel metal2 s 140962 15200 141018 16000 0 FreeSans 224 90 0 0 dq[238]
port 153 nsew signal tristate
flabel metal2 s 141514 15200 141570 16000 0 FreeSans 224 90 0 0 dq[239]
port 154 nsew signal tristate
flabel metal2 s 22282 15200 22338 16000 0 FreeSans 224 90 0 0 dq[23]
port 155 nsew signal tristate
flabel metal2 s 142066 15200 142122 16000 0 FreeSans 224 90 0 0 dq[240]
port 156 nsew signal tristate
flabel metal2 s 142618 15200 142674 16000 0 FreeSans 224 90 0 0 dq[241]
port 157 nsew signal tristate
flabel metal2 s 143170 15200 143226 16000 0 FreeSans 224 90 0 0 dq[242]
port 158 nsew signal tristate
flabel metal2 s 143722 15200 143778 16000 0 FreeSans 224 90 0 0 dq[243]
port 159 nsew signal tristate
flabel metal2 s 144274 15200 144330 16000 0 FreeSans 224 90 0 0 dq[244]
port 160 nsew signal tristate
flabel metal2 s 144826 15200 144882 16000 0 FreeSans 224 90 0 0 dq[245]
port 161 nsew signal tristate
flabel metal2 s 145378 15200 145434 16000 0 FreeSans 224 90 0 0 dq[246]
port 162 nsew signal tristate
flabel metal2 s 145930 15200 145986 16000 0 FreeSans 224 90 0 0 dq[247]
port 163 nsew signal tristate
flabel metal2 s 146482 15200 146538 16000 0 FreeSans 224 90 0 0 dq[248]
port 164 nsew signal tristate
flabel metal2 s 147034 15200 147090 16000 0 FreeSans 224 90 0 0 dq[249]
port 165 nsew signal tristate
flabel metal2 s 22834 15200 22890 16000 0 FreeSans 224 90 0 0 dq[24]
port 166 nsew signal tristate
flabel metal2 s 147586 15200 147642 16000 0 FreeSans 224 90 0 0 dq[250]
port 167 nsew signal tristate
flabel metal2 s 148138 15200 148194 16000 0 FreeSans 224 90 0 0 dq[251]
port 168 nsew signal tristate
flabel metal2 s 148690 15200 148746 16000 0 FreeSans 224 90 0 0 dq[252]
port 169 nsew signal tristate
flabel metal2 s 149242 15200 149298 16000 0 FreeSans 224 90 0 0 dq[253]
port 170 nsew signal tristate
flabel metal2 s 149794 15200 149850 16000 0 FreeSans 224 90 0 0 dq[254]
port 171 nsew signal tristate
flabel metal2 s 150346 15200 150402 16000 0 FreeSans 224 90 0 0 dq[255]
port 172 nsew signal tristate
flabel metal2 s 23386 15200 23442 16000 0 FreeSans 224 90 0 0 dq[25]
port 173 nsew signal tristate
flabel metal2 s 23938 15200 23994 16000 0 FreeSans 224 90 0 0 dq[26]
port 174 nsew signal tristate
flabel metal2 s 24490 15200 24546 16000 0 FreeSans 224 90 0 0 dq[27]
port 175 nsew signal tristate
flabel metal2 s 25042 15200 25098 16000 0 FreeSans 224 90 0 0 dq[28]
port 176 nsew signal tristate
flabel metal2 s 25594 15200 25650 16000 0 FreeSans 224 90 0 0 dq[29]
port 177 nsew signal tristate
flabel metal2 s 10690 15200 10746 16000 0 FreeSans 224 90 0 0 dq[2]
port 178 nsew signal tristate
flabel metal2 s 26146 15200 26202 16000 0 FreeSans 224 90 0 0 dq[30]
port 179 nsew signal tristate
flabel metal2 s 26698 15200 26754 16000 0 FreeSans 224 90 0 0 dq[31]
port 180 nsew signal tristate
flabel metal2 s 27250 15200 27306 16000 0 FreeSans 224 90 0 0 dq[32]
port 181 nsew signal tristate
flabel metal2 s 27802 15200 27858 16000 0 FreeSans 224 90 0 0 dq[33]
port 182 nsew signal tristate
flabel metal2 s 28354 15200 28410 16000 0 FreeSans 224 90 0 0 dq[34]
port 183 nsew signal tristate
flabel metal2 s 28906 15200 28962 16000 0 FreeSans 224 90 0 0 dq[35]
port 184 nsew signal tristate
flabel metal2 s 29458 15200 29514 16000 0 FreeSans 224 90 0 0 dq[36]
port 185 nsew signal tristate
flabel metal2 s 30010 15200 30066 16000 0 FreeSans 224 90 0 0 dq[37]
port 186 nsew signal tristate
flabel metal2 s 30562 15200 30618 16000 0 FreeSans 224 90 0 0 dq[38]
port 187 nsew signal tristate
flabel metal2 s 31114 15200 31170 16000 0 FreeSans 224 90 0 0 dq[39]
port 188 nsew signal tristate
flabel metal2 s 11242 15200 11298 16000 0 FreeSans 224 90 0 0 dq[3]
port 189 nsew signal tristate
flabel metal2 s 31666 15200 31722 16000 0 FreeSans 224 90 0 0 dq[40]
port 190 nsew signal tristate
flabel metal2 s 32218 15200 32274 16000 0 FreeSans 224 90 0 0 dq[41]
port 191 nsew signal tristate
flabel metal2 s 32770 15200 32826 16000 0 FreeSans 224 90 0 0 dq[42]
port 192 nsew signal tristate
flabel metal2 s 33322 15200 33378 16000 0 FreeSans 224 90 0 0 dq[43]
port 193 nsew signal tristate
flabel metal2 s 33874 15200 33930 16000 0 FreeSans 224 90 0 0 dq[44]
port 194 nsew signal tristate
flabel metal2 s 34426 15200 34482 16000 0 FreeSans 224 90 0 0 dq[45]
port 195 nsew signal tristate
flabel metal2 s 34978 15200 35034 16000 0 FreeSans 224 90 0 0 dq[46]
port 196 nsew signal tristate
flabel metal2 s 35530 15200 35586 16000 0 FreeSans 224 90 0 0 dq[47]
port 197 nsew signal tristate
flabel metal2 s 36082 15200 36138 16000 0 FreeSans 224 90 0 0 dq[48]
port 198 nsew signal tristate
flabel metal2 s 36634 15200 36690 16000 0 FreeSans 224 90 0 0 dq[49]
port 199 nsew signal tristate
flabel metal2 s 11794 15200 11850 16000 0 FreeSans 224 90 0 0 dq[4]
port 200 nsew signal tristate
flabel metal2 s 37186 15200 37242 16000 0 FreeSans 224 90 0 0 dq[50]
port 201 nsew signal tristate
flabel metal2 s 37738 15200 37794 16000 0 FreeSans 224 90 0 0 dq[51]
port 202 nsew signal tristate
flabel metal2 s 38290 15200 38346 16000 0 FreeSans 224 90 0 0 dq[52]
port 203 nsew signal tristate
flabel metal2 s 38842 15200 38898 16000 0 FreeSans 224 90 0 0 dq[53]
port 204 nsew signal tristate
flabel metal2 s 39394 15200 39450 16000 0 FreeSans 224 90 0 0 dq[54]
port 205 nsew signal tristate
flabel metal2 s 39946 15200 40002 16000 0 FreeSans 224 90 0 0 dq[55]
port 206 nsew signal tristate
flabel metal2 s 40498 15200 40554 16000 0 FreeSans 224 90 0 0 dq[56]
port 207 nsew signal tristate
flabel metal2 s 41050 15200 41106 16000 0 FreeSans 224 90 0 0 dq[57]
port 208 nsew signal tristate
flabel metal2 s 41602 15200 41658 16000 0 FreeSans 224 90 0 0 dq[58]
port 209 nsew signal tristate
flabel metal2 s 42154 15200 42210 16000 0 FreeSans 224 90 0 0 dq[59]
port 210 nsew signal tristate
flabel metal2 s 12346 15200 12402 16000 0 FreeSans 224 90 0 0 dq[5]
port 211 nsew signal tristate
flabel metal2 s 42706 15200 42762 16000 0 FreeSans 224 90 0 0 dq[60]
port 212 nsew signal tristate
flabel metal2 s 43258 15200 43314 16000 0 FreeSans 224 90 0 0 dq[61]
port 213 nsew signal tristate
flabel metal2 s 43810 15200 43866 16000 0 FreeSans 224 90 0 0 dq[62]
port 214 nsew signal tristate
flabel metal2 s 44362 15200 44418 16000 0 FreeSans 224 90 0 0 dq[63]
port 215 nsew signal tristate
flabel metal2 s 44914 15200 44970 16000 0 FreeSans 224 90 0 0 dq[64]
port 216 nsew signal tristate
flabel metal2 s 45466 15200 45522 16000 0 FreeSans 224 90 0 0 dq[65]
port 217 nsew signal tristate
flabel metal2 s 46018 15200 46074 16000 0 FreeSans 224 90 0 0 dq[66]
port 218 nsew signal tristate
flabel metal2 s 46570 15200 46626 16000 0 FreeSans 224 90 0 0 dq[67]
port 219 nsew signal tristate
flabel metal2 s 47122 15200 47178 16000 0 FreeSans 224 90 0 0 dq[68]
port 220 nsew signal tristate
flabel metal2 s 47674 15200 47730 16000 0 FreeSans 224 90 0 0 dq[69]
port 221 nsew signal tristate
flabel metal2 s 12898 15200 12954 16000 0 FreeSans 224 90 0 0 dq[6]
port 222 nsew signal tristate
flabel metal2 s 48226 15200 48282 16000 0 FreeSans 224 90 0 0 dq[70]
port 223 nsew signal tristate
flabel metal2 s 48778 15200 48834 16000 0 FreeSans 224 90 0 0 dq[71]
port 224 nsew signal tristate
flabel metal2 s 49330 15200 49386 16000 0 FreeSans 224 90 0 0 dq[72]
port 225 nsew signal tristate
flabel metal2 s 49882 15200 49938 16000 0 FreeSans 224 90 0 0 dq[73]
port 226 nsew signal tristate
flabel metal2 s 50434 15200 50490 16000 0 FreeSans 224 90 0 0 dq[74]
port 227 nsew signal tristate
flabel metal2 s 50986 15200 51042 16000 0 FreeSans 224 90 0 0 dq[75]
port 228 nsew signal tristate
flabel metal2 s 51538 15200 51594 16000 0 FreeSans 224 90 0 0 dq[76]
port 229 nsew signal tristate
flabel metal2 s 52090 15200 52146 16000 0 FreeSans 224 90 0 0 dq[77]
port 230 nsew signal tristate
flabel metal2 s 52642 15200 52698 16000 0 FreeSans 224 90 0 0 dq[78]
port 231 nsew signal tristate
flabel metal2 s 53194 15200 53250 16000 0 FreeSans 224 90 0 0 dq[79]
port 232 nsew signal tristate
flabel metal2 s 13450 15200 13506 16000 0 FreeSans 224 90 0 0 dq[7]
port 233 nsew signal tristate
flabel metal2 s 53746 15200 53802 16000 0 FreeSans 224 90 0 0 dq[80]
port 234 nsew signal tristate
flabel metal2 s 54298 15200 54354 16000 0 FreeSans 224 90 0 0 dq[81]
port 235 nsew signal tristate
flabel metal2 s 54850 15200 54906 16000 0 FreeSans 224 90 0 0 dq[82]
port 236 nsew signal tristate
flabel metal2 s 55402 15200 55458 16000 0 FreeSans 224 90 0 0 dq[83]
port 237 nsew signal tristate
flabel metal2 s 55954 15200 56010 16000 0 FreeSans 224 90 0 0 dq[84]
port 238 nsew signal tristate
flabel metal2 s 56506 15200 56562 16000 0 FreeSans 224 90 0 0 dq[85]
port 239 nsew signal tristate
flabel metal2 s 57058 15200 57114 16000 0 FreeSans 224 90 0 0 dq[86]
port 240 nsew signal tristate
flabel metal2 s 57610 15200 57666 16000 0 FreeSans 224 90 0 0 dq[87]
port 241 nsew signal tristate
flabel metal2 s 58162 15200 58218 16000 0 FreeSans 224 90 0 0 dq[88]
port 242 nsew signal tristate
flabel metal2 s 58714 15200 58770 16000 0 FreeSans 224 90 0 0 dq[89]
port 243 nsew signal tristate
flabel metal2 s 14002 15200 14058 16000 0 FreeSans 224 90 0 0 dq[8]
port 244 nsew signal tristate
flabel metal2 s 59266 15200 59322 16000 0 FreeSans 224 90 0 0 dq[90]
port 245 nsew signal tristate
flabel metal2 s 59818 15200 59874 16000 0 FreeSans 224 90 0 0 dq[91]
port 246 nsew signal tristate
flabel metal2 s 60370 15200 60426 16000 0 FreeSans 224 90 0 0 dq[92]
port 247 nsew signal tristate
flabel metal2 s 60922 15200 60978 16000 0 FreeSans 224 90 0 0 dq[93]
port 248 nsew signal tristate
flabel metal2 s 61474 15200 61530 16000 0 FreeSans 224 90 0 0 dq[94]
port 249 nsew signal tristate
flabel metal2 s 62026 15200 62082 16000 0 FreeSans 224 90 0 0 dq[95]
port 250 nsew signal tristate
flabel metal2 s 62578 15200 62634 16000 0 FreeSans 224 90 0 0 dq[96]
port 251 nsew signal tristate
flabel metal2 s 63130 15200 63186 16000 0 FreeSans 224 90 0 0 dq[97]
port 252 nsew signal tristate
flabel metal2 s 63682 15200 63738 16000 0 FreeSans 224 90 0 0 dq[98]
port 253 nsew signal tristate
flabel metal2 s 64234 15200 64290 16000 0 FreeSans 224 90 0 0 dq[99]
port 254 nsew signal tristate
flabel metal2 s 14554 15200 14610 16000 0 FreeSans 224 90 0 0 dq[9]
port 255 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 latch
port 256 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 rst_n
port 257 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 sclk
port 258 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 sdi
port 259 nsew signal input
flabel metal3 s 159200 7896 160000 8016 0 FreeSans 480 0 0 0 sdo
port 260 nsew signal tristate
flabel metal4 s 20666 2128 20986 13648 0 FreeSans 1920 90 0 0 vccd1
port 261 nsew power bidirectional
flabel metal4 s 60111 2128 60431 13648 0 FreeSans 1920 90 0 0 vccd1
port 261 nsew power bidirectional
flabel metal4 s 99556 2128 99876 13648 0 FreeSans 1920 90 0 0 vccd1
port 261 nsew power bidirectional
flabel metal4 s 139001 2128 139321 13648 0 FreeSans 1920 90 0 0 vccd1
port 261 nsew power bidirectional
flabel metal4 s 40388 2128 40708 13648 0 FreeSans 1920 90 0 0 vssd1
port 262 nsew ground bidirectional
flabel metal4 s 79833 2128 80153 13648 0 FreeSans 1920 90 0 0 vssd1
port 262 nsew ground bidirectional
flabel metal4 s 119278 2128 119598 13648 0 FreeSans 1920 90 0 0 vssd1
port 262 nsew ground bidirectional
flabel metal4 s 158723 2128 159043 13648 0 FreeSans 1920 90 0 0 vssd1
port 262 nsew ground bidirectional
rlabel metal1 79994 13600 79994 13600 0 vccd1
rlabel via1 80073 13056 80073 13056 0 vssd1
rlabel metal1 150558 5542 150558 5542 0 _0000_
rlabel via2 136390 7803 136390 7803 0 _0001_
rlabel metal2 155986 2839 155986 2839 0 _0002_
rlabel metal1 151340 12614 151340 12614 0 _0003_
rlabel metal2 148810 3587 148810 3587 0 _0004_
rlabel metal2 155986 2074 155986 2074 0 _0005_
rlabel via1 143929 8466 143929 8466 0 _0006_
rlabel metal2 153502 3111 153502 3111 0 _0007_
rlabel metal1 121573 8534 121573 8534 0 _0008_
rlabel metal1 129459 4522 129459 4522 0 _0009_
rlabel metal1 126684 2822 126684 2822 0 _0010_
rlabel metal2 157274 4862 157274 4862 0 _0011_
rlabel metal1 147154 4556 147154 4556 0 _0012_
rlabel metal2 150466 6375 150466 6375 0 _0013_
rlabel metal1 151156 5814 151156 5814 0 _0014_
rlabel metal2 149178 2142 149178 2142 0 _0015_
rlabel metal1 155940 2278 155940 2278 0 _0016_
rlabel metal1 152536 13158 152536 13158 0 _0017_
rlabel metal1 151524 6630 151524 6630 0 _0018_
rlabel metal1 150650 6630 150650 6630 0 _0019_
rlabel metal1 156584 8058 156584 8058 0 _0020_
rlabel metal2 151662 7344 151662 7344 0 _0021_
rlabel metal1 144286 3434 144286 3434 0 _0022_
rlabel metal1 144118 9418 144118 9418 0 _0023_
rlabel metal1 146326 5644 146326 5644 0 _0024_
rlabel via1 137581 3094 137581 3094 0 _0025_
rlabel metal1 140760 5338 140760 5338 0 _0026_
rlabel metal1 139855 5610 139855 5610 0 _0027_
rlabel metal1 137586 4556 137586 4556 0 _0028_
rlabel metal2 140714 8704 140714 8704 0 _0029_
rlabel metal1 141864 2822 141864 2822 0 _0030_
rlabel metal1 147706 3604 147706 3604 0 _0031_
rlabel metal2 117898 10540 117898 10540 0 _0032_
rlabel metal1 109996 2414 109996 2414 0 _0033_
rlabel metal1 114765 7786 114765 7786 0 _0034_
rlabel metal1 112286 10030 112286 10030 0 _0035_
rlabel metal1 112715 12886 112715 12886 0 _0036_
rlabel metal1 96922 10132 96922 10132 0 _0037_
rlabel metal1 107440 6358 107440 6358 0 _0038_
rlabel metal1 110962 4114 110962 4114 0 _0039_
rlabel via1 97377 6290 97377 6290 0 _0040_
rlabel metal1 102181 10710 102181 10710 0 _0041_
rlabel metal2 83490 8670 83490 8670 0 _0042_
rlabel metal1 106214 8330 106214 8330 0 _0043_
rlabel metal1 19642 9928 19642 9928 0 _0044_
rlabel via1 12093 10710 12093 10710 0 _0045_
rlabel metal1 17475 11118 17475 11118 0 _0046_
rlabel metal1 19090 6154 19090 6154 0 _0047_
rlabel metal1 14996 6426 14996 6426 0 _0048_
rlabel metal2 14582 9180 14582 9180 0 _0049_
rlabel metal1 13390 8534 13390 8534 0 _0050_
rlabel viali 14577 5678 14577 5678 0 _0051_
rlabel metal2 19918 6018 19918 6018 0 _0052_
rlabel metal1 22662 3094 22662 3094 0 _0053_
rlabel metal1 17940 3162 17940 3162 0 _0054_
rlabel metal2 15686 7650 15686 7650 0 _0055_
rlabel metal1 19596 5882 19596 5882 0 _0056_
rlabel metal1 19074 3434 19074 3434 0 _0057_
rlabel metal1 12783 5202 12783 5202 0 _0058_
rlabel via1 16509 6766 16509 6766 0 _0059_
rlabel metal1 19412 2550 19412 2550 0 _0060_
rlabel metal1 18430 3094 18430 3094 0 _0061_
rlabel via1 23041 5270 23041 5270 0 _0062_
rlabel metal1 26680 8058 26680 8058 0 _0063_
rlabel metal2 21114 7650 21114 7650 0 _0064_
rlabel metal1 24840 5882 24840 5882 0 _0065_
rlabel metal2 26910 8092 26910 8092 0 _0066_
rlabel via1 17070 4590 17070 4590 0 _0067_
rlabel metal1 4324 6630 4324 6630 0 _0068_
rlabel metal2 5014 7378 5014 7378 0 _0069_
rlabel metal1 4457 5678 4457 5678 0 _0070_
rlabel metal1 4135 10710 4135 10710 0 _0071_
rlabel metal2 5290 8194 5290 8194 0 _0072_
rlabel metal1 12466 11152 12466 11152 0 _0073_
rlabel metal1 5796 5882 5796 5882 0 _0074_
rlabel metal1 7498 3978 7498 3978 0 _0075_
rlabel metal2 14122 8534 14122 8534 0 _0076_
rlabel metal1 4917 5202 4917 5202 0 _0077_
rlabel metal1 13846 3162 13846 3162 0 _0078_
rlabel metal2 11730 9384 11730 9384 0 _0079_
rlabel metal1 15272 10506 15272 10506 0 _0080_
rlabel metal1 13125 3094 13125 3094 0 _0081_
rlabel metal1 12519 8874 12519 8874 0 _0082_
rlabel metal1 24232 2414 24232 2414 0 _0083_
rlabel metal1 15368 13226 15368 13226 0 _0084_
rlabel metal1 13554 9962 13554 9962 0 _0085_
rlabel metal2 16330 9928 16330 9928 0 _0086_
rlabel metal2 37490 6120 37490 6120 0 _0087_
rlabel metal2 46874 7208 46874 7208 0 _0088_
rlabel metal1 43940 8466 43940 8466 0 _0089_
rlabel metal1 46506 6392 46506 6392 0 _0090_
rlabel via1 49546 9962 49546 9962 0 _0091_
rlabel metal1 41400 9894 41400 9894 0 _0092_
rlabel metal1 53249 4114 53249 4114 0 _0093_
rlabel metal1 36708 8058 36708 8058 0 _0094_
rlabel metal1 38788 9554 38788 9554 0 _0095_
rlabel metal1 37858 8058 37858 8058 0 _0096_
rlabel metal1 36580 5202 36580 5202 0 _0097_
rlabel metal2 33350 9078 33350 9078 0 _0098_
rlabel metal1 38364 5882 38364 5882 0 _0099_
rlabel metal1 37260 7990 37260 7990 0 _0100_
rlabel metal2 34086 6426 34086 6426 0 _0101_
rlabel metal2 31602 9010 31602 9010 0 _0102_
rlabel metal2 30774 7174 30774 7174 0 _0103_
rlabel metal1 32614 9928 32614 9928 0 _0104_
rlabel metal2 33534 10846 33534 10846 0 _0105_
rlabel metal1 29337 8874 29337 8874 0 _0106_
rlabel metal1 38072 7446 38072 7446 0 _0107_
rlabel metal1 42580 12886 42580 12886 0 _0108_
rlabel metal1 43557 4522 43557 4522 0 _0109_
rlabel metal1 45540 10030 45540 10030 0 _0110_
rlabel metal1 47702 3910 47702 3910 0 _0111_
rlabel via1 46418 8534 46418 8534 0 _0112_
rlabel metal1 34975 6358 34975 6358 0 _0113_
rlabel metal1 41446 7480 41446 7480 0 _0114_
rlabel via1 48065 3026 48065 3026 0 _0115_
rlabel metal1 53697 5610 53697 5610 0 _0116_
rlabel via1 43557 10030 43557 10030 0 _0117_
rlabel metal1 45954 5338 45954 5338 0 _0118_
rlabel metal1 56488 12886 56488 12886 0 _0119_
rlabel via1 40981 9622 40981 9622 0 _0120_
rlabel metal2 42872 11900 42872 11900 0 _0121_
rlabel via1 56437 3094 56437 3094 0 _0122_
rlabel metal1 61538 2414 61538 2414 0 _0123_
rlabel metal2 64906 3876 64906 3876 0 _0124_
rlabel metal1 58384 3502 58384 3502 0 _0125_
rlabel metal1 47012 12954 47012 12954 0 _0126_
rlabel metal2 63986 8058 63986 8058 0 _0127_
rlabel metal2 60674 13362 60674 13362 0 _0128_
rlabel metal1 54142 9622 54142 9622 0 _0129_
rlabel metal1 52900 11866 52900 11866 0 _0130_
rlabel metal1 58052 12614 58052 12614 0 _0131_
rlabel metal1 57960 7514 57960 7514 0 _0132_
rlabel metal1 75076 9554 75076 9554 0 _0133_
rlabel metal2 64814 9282 64814 9282 0 _0134_
rlabel metal2 53222 8194 53222 8194 0 _0135_
rlabel metal1 53467 7446 53467 7446 0 _0136_
rlabel metal1 56304 8330 56304 8330 0 _0137_
rlabel metal1 57812 2414 57812 2414 0 _0138_
rlabel metal1 63976 5678 63976 5678 0 _0139_
rlabel metal1 62432 7854 62432 7854 0 _0140_
rlabel metal1 56902 9350 56902 9350 0 _0141_
rlabel metal1 61216 5202 61216 5202 0 _0142_
rlabel metal2 63250 9282 63250 9282 0 _0143_
rlabel metal2 67114 7650 67114 7650 0 _0144_
rlabel metal1 77280 9418 77280 9418 0 _0145_
rlabel metal2 73370 5746 73370 5746 0 _0146_
rlabel metal1 64680 6766 64680 6766 0 _0147_
rlabel metal1 92935 12138 92935 12138 0 _0148_
rlabel metal1 66000 8942 66000 8942 0 _0149_
rlabel metal1 73089 7854 73089 7854 0 _0150_
rlabel metal1 86250 4794 86250 4794 0 _0151_
rlabel metal2 91402 7820 91402 7820 0 _0152_
rlabel metal1 78062 5066 78062 5066 0 _0153_
rlabel metal1 75685 6698 75685 6698 0 _0154_
rlabel metal2 79902 9333 79902 9333 0 _0155_
rlabel metal1 89000 4590 89000 4590 0 _0156_
rlabel metal1 81737 9962 81737 9962 0 _0157_
rlabel metal1 84088 7174 84088 7174 0 _0158_
rlabel metal1 95736 3502 95736 3502 0 _0159_
rlabel metal1 82815 2346 82815 2346 0 _0160_
rlabel metal2 82846 11288 82846 11288 0 _0161_
rlabel metal1 92322 6800 92322 6800 0 _0162_
rlabel metal2 97566 7718 97566 7718 0 _0163_
rlabel via1 96558 7378 96558 7378 0 _0164_
rlabel metal1 98026 9928 98026 9928 0 _0165_
rlabel metal1 93748 5066 93748 5066 0 _0166_
rlabel metal1 79115 9962 79115 9962 0 _0167_
rlabel metal1 75864 7378 75864 7378 0 _0168_
rlabel metal1 116932 9146 116932 9146 0 _0169_
rlabel metal2 116334 7310 116334 7310 0 _0170_
rlabel metal1 97075 12138 97075 12138 0 _0171_
rlabel via2 77326 12155 77326 12155 0 _0172_
rlabel metal2 108698 8398 108698 8398 0 _0173_
rlabel metal2 109526 5287 109526 5287 0 _0174_
rlabel metal2 115690 6868 115690 6868 0 _0175_
rlabel metal1 92516 5202 92516 5202 0 _0176_
rlabel via1 116614 9622 116614 9622 0 _0177_
rlabel metal1 113850 5848 113850 5848 0 _0178_
rlabel metal1 128892 10642 128892 10642 0 _0179_
rlabel metal1 110170 2890 110170 2890 0 _0180_
rlabel metal1 122738 7378 122738 7378 0 _0181_
rlabel metal2 129766 8041 129766 8041 0 _0182_
rlabel metal2 112194 4726 112194 4726 0 _0183_
rlabel metal1 133032 7922 133032 7922 0 _0184_
rlabel via2 76406 4539 76406 4539 0 _0185_
rlabel metal2 133078 13328 133078 13328 0 _0186_
rlabel metal2 98302 10234 98302 10234 0 _0187_
rlabel metal1 128662 8330 128662 8330 0 _0188_
rlabel metal2 94438 10914 94438 10914 0 _0189_
rlabel via1 93982 9962 93982 9962 0 _0190_
rlabel metal2 95358 9384 95358 9384 0 _0191_
rlabel metal1 117898 3944 117898 3944 0 _0192_
rlabel via2 87262 10523 87262 10523 0 _0193_
rlabel metal1 97244 9690 97244 9690 0 _0194_
rlabel metal1 72828 7378 72828 7378 0 _0195_
rlabel metal1 97791 4522 97791 4522 0 _0196_
rlabel metal1 132142 8534 132142 8534 0 _0197_
rlabel metal2 155710 9112 155710 9112 0 _0198_
rlabel metal2 156630 2176 156630 2176 0 _0199_
rlabel metal2 157090 11645 157090 11645 0 _0200_
rlabel metal1 147798 3128 147798 3128 0 _0201_
rlabel metal1 133446 12104 133446 12104 0 _0202_
rlabel metal1 136727 6698 136727 6698 0 _0203_
rlabel metal1 148212 13974 148212 13974 0 _0204_
rlabel via1 139890 7786 139890 7786 0 _0205_
rlabel metal2 147890 2040 147890 2040 0 _0206_
rlabel metal1 135485 9962 135485 9962 0 _0207_
rlabel metal2 157274 4352 157274 4352 0 _0208_
rlabel metal1 153272 4998 153272 4998 0 _0209_
rlabel metal2 130226 8500 130226 8500 0 _0210_
rlabel metal1 135746 8500 135746 8500 0 _0211_
rlabel metal1 155664 4454 155664 4454 0 _0212_
rlabel via2 117438 5899 117438 5899 0 _0213_
rlabel metal2 147522 2108 147522 2108 0 _0214_
rlabel metal2 110262 2043 110262 2043 0 _0215_
rlabel metal1 134458 2584 134458 2584 0 _0216_
rlabel metal1 109480 3162 109480 3162 0 _0217_
rlabel metal2 118082 4862 118082 4862 0 _0218_
rlabel metal1 118358 5746 118358 5746 0 _0219_
rlabel via1 120193 5270 120193 5270 0 _0220_
rlabel viali 121398 6698 121398 6698 0 _0221_
rlabel via2 156814 5355 156814 5355 0 _0222_
rlabel metal1 156262 3638 156262 3638 0 _0223_
rlabel metal2 156814 5984 156814 5984 0 _0224_
rlabel metal1 151708 5542 151708 5542 0 _0225_
rlabel metal3 152444 7072 152444 7072 0 _0226_
rlabel via1 142926 4114 142926 4114 0 _0227_
rlabel metal1 148442 13192 148442 13192 0 _0228_
rlabel metal2 129214 1907 129214 1907 0 _0229_
rlabel metal1 108652 9418 108652 9418 0 _0230_
rlabel metal1 119002 3502 119002 3502 0 _0231_
rlabel via1 135649 2414 135649 2414 0 _0232_
rlabel via2 143842 6341 143842 6341 0 _0233_
rlabel metal2 144946 9877 144946 9877 0 _0234_
rlabel metal2 156446 1921 156446 1921 0 _0235_
rlabel metal2 147798 1666 147798 1666 0 _0236_
rlabel metal1 132802 12954 132802 12954 0 _0237_
rlabel via2 156814 3893 156814 3893 0 _0238_
rlabel metal2 145866 4658 145866 4658 0 _0239_
rlabel metal1 150650 11322 150650 11322 0 _0240_
rlabel metal2 128570 2176 128570 2176 0 _0241_
rlabel metal2 158102 13430 158102 13430 0 _0242_
rlabel metal2 155434 10846 155434 10846 0 _0243_
rlabel metal1 143750 5168 143750 5168 0 _0244_
rlabel metal2 141450 10064 141450 10064 0 _0245_
rlabel metal1 140990 10744 140990 10744 0 _0246_
rlabel metal1 150696 9486 150696 9486 0 _0247_
rlabel metal1 143980 13158 143980 13158 0 _0248_
rlabel metal1 153548 6970 153548 6970 0 _0249_
rlabel metal1 148345 12818 148345 12818 0 _0250_
rlabel metal1 148713 7786 148713 7786 0 _0251_
rlabel metal1 148718 11526 148718 11526 0 _0252_
rlabel metal1 149592 10438 149592 10438 0 _0253_
rlabel via1 143377 5610 143377 5610 0 _0254_
rlabel metal1 140300 4726 140300 4726 0 _0255_
rlabel metal1 153594 7378 153594 7378 0 _0256_
rlabel via1 109158 12597 109158 12597 0 _0257_
rlabel metal1 126822 3706 126822 3706 0 _0258_
rlabel metal1 111182 9554 111182 9554 0 _0259_
rlabel metal1 110952 7310 110952 7310 0 _0260_
rlabel metal2 114586 8738 114586 8738 0 _0261_
rlabel metal1 113574 11730 113574 11730 0 _0262_
rlabel metal1 111228 8942 111228 8942 0 _0263_
rlabel metal1 105570 7854 105570 7854 0 _0264_
rlabel metal2 111642 11594 111642 11594 0 _0265_
rlabel metal2 108790 11526 108790 11526 0 _0266_
rlabel metal1 102810 13158 102810 13158 0 _0267_
rlabel metal1 32154 5848 32154 5848 0 _0268_
rlabel metal2 84594 10132 84594 10132 0 _0269_
rlabel metal1 112608 7990 112608 7990 0 _0270_
rlabel metal1 19458 10132 19458 10132 0 _0271_
rlabel metal2 19366 11305 19366 11305 0 _0272_
rlabel metal2 18630 11356 18630 11356 0 _0273_
rlabel metal1 18354 6290 18354 6290 0 _0274_
rlabel metal1 15686 5882 15686 5882 0 _0275_
rlabel metal2 14398 7786 14398 7786 0 _0276_
rlabel metal1 13156 12614 13156 12614 0 _0277_
rlabel metal1 12236 12614 12236 12614 0 _0278_
rlabel metal2 17250 5134 17250 5134 0 _0279_
rlabel metal1 20792 3026 20792 3026 0 _0280_
rlabel metal2 16882 4828 16882 4828 0 _0281_
rlabel metal2 15686 5202 15686 5202 0 _0282_
rlabel metal2 19826 7038 19826 7038 0 _0283_
rlabel metal2 16882 9180 16882 9180 0 _0284_
rlabel metal2 17710 5100 17710 5100 0 _0285_
rlabel metal1 12742 4794 12742 4794 0 _0286_
rlabel metal1 14628 4794 14628 4794 0 _0287_
rlabel metal1 16606 8058 16606 8058 0 _0288_
rlabel metal1 18078 2414 18078 2414 0 _0289_
rlabel metal1 18124 6902 18124 6902 0 _0290_
rlabel metal2 21298 7140 21298 7140 0 _0291_
rlabel metal1 25806 3706 25806 3706 0 _0292_
rlabel metal2 21666 9622 21666 9622 0 _0293_
rlabel metal1 23506 5678 23506 5678 0 _0294_
rlabel metal1 26634 4794 26634 4794 0 _0295_
rlabel metal1 19596 9554 19596 9554 0 _0296_
rlabel metal1 11730 2482 11730 2482 0 _0297_
rlabel metal1 5014 2618 5014 2618 0 _0298_
rlabel metal1 5290 4590 5290 4590 0 _0299_
rlabel metal2 4830 7548 4830 7548 0 _0300_
rlabel metal2 4462 11764 4462 11764 0 _0301_
rlabel metal1 5290 7378 5290 7378 0 _0302_
rlabel metal1 11822 11118 11822 11118 0 _0303_
rlabel metal1 6072 5678 6072 5678 0 _0304_
rlabel metal1 8740 4114 8740 4114 0 _0305_
rlabel metal1 13984 7378 13984 7378 0 _0306_
rlabel metal2 11822 7786 11822 7786 0 _0307_
rlabel metal1 16652 10030 16652 10030 0 _0308_
rlabel metal2 13570 3196 13570 3196 0 _0309_
rlabel metal1 13340 4794 13340 4794 0 _0310_
rlabel metal2 15410 10132 15410 10132 0 _0311_
rlabel metal2 13570 8874 13570 8874 0 _0312_
rlabel metal2 12190 6698 12190 6698 0 _0313_
rlabel metal2 21206 7854 21206 7854 0 _0314_
rlabel metal1 16790 5882 16790 5882 0 _0315_
rlabel metal1 10994 11764 10994 11764 0 _0316_
rlabel metal1 16422 3706 16422 3706 0 _0317_
rlabel metal2 23966 6834 23966 6834 0 _0318_
rlabel metal1 45678 2380 45678 2380 0 _0319_
rlabel metal2 53774 5610 53774 5610 0 _0320_
rlabel metal2 50462 9520 50462 9520 0 _0321_
rlabel metal2 46690 7004 46690 7004 0 _0322_
rlabel metal2 50462 10812 50462 10812 0 _0323_
rlabel metal1 40802 10064 40802 10064 0 _0324_
rlabel metal2 42642 11577 42642 11577 0 _0325_
rlabel metal1 36984 3706 36984 3706 0 _0326_
rlabel metal1 43378 2618 43378 2618 0 _0327_
rlabel metal1 38594 7888 38594 7888 0 _0328_
rlabel metal2 39330 8058 39330 8058 0 _0329_
rlabel via2 89286 13243 89286 13243 0 _0330_
rlabel metal1 37628 10778 37628 10778 0 _0331_
rlabel metal2 33166 7888 33166 7888 0 _0332_
rlabel metal2 37858 6256 37858 6256 0 _0333_
rlabel metal2 35374 8942 35374 8942 0 _0334_
rlabel metal1 35144 5202 35144 5202 0 _0335_
rlabel metal1 32706 7854 32706 7854 0 _0336_
rlabel metal1 30636 4590 30636 4590 0 _0337_
rlabel metal1 32752 3162 32752 3162 0 _0338_
rlabel metal1 31878 11084 31878 11084 0 _0339_
rlabel metal2 27186 9996 27186 9996 0 _0340_
rlabel metal1 36524 7378 36524 7378 0 _0341_
rlabel metal1 40802 13294 40802 13294 0 _0342_
rlabel metal1 40112 13158 40112 13158 0 _0343_
rlabel metal1 44436 8466 44436 8466 0 _0344_
rlabel metal1 45908 4590 45908 4590 0 _0345_
rlabel metal2 47978 5916 47978 5916 0 _0346_
rlabel metal1 45218 8976 45218 8976 0 _0347_
rlabel metal2 36570 7548 36570 7548 0 _0348_
rlabel metal1 40940 6426 40940 6426 0 _0349_
rlabel metal1 47518 9690 47518 9690 0 _0350_
rlabel metal2 54234 5916 54234 5916 0 _0351_
rlabel metal2 45402 11305 45402 11305 0 _0352_
rlabel metal1 36248 12614 36248 12614 0 _0353_
rlabel metal2 48714 7276 48714 7276 0 _0354_
rlabel metal1 57270 8908 57270 8908 0 _0355_
rlabel metal1 41216 8466 41216 8466 0 _0356_
rlabel metal1 42366 13294 42366 13294 0 _0357_
rlabel metal1 55844 8942 55844 8942 0 _0358_
rlabel metal1 52670 7854 52670 7854 0 _0359_
rlabel metal1 65458 3502 65458 3502 0 _0360_
rlabel metal2 58650 6154 58650 6154 0 _0361_
rlabel metal2 51014 6256 51014 6256 0 _0362_
rlabel metal1 56534 6188 56534 6188 0 _0363_
rlabel metal1 51658 10030 51658 10030 0 _0364_
rlabel metal2 56120 13226 56120 13226 0 _0365_
rlabel metal2 58098 10030 58098 10030 0 _0366_
rlabel metal1 52348 10234 52348 10234 0 _0367_
rlabel metal1 58788 12410 58788 12410 0 _0368_
rlabel metal1 59156 7378 59156 7378 0 _0369_
rlabel metal1 63940 13158 63940 13158 0 _0370_
rlabel metal2 64630 8908 64630 8908 0 _0371_
rlabel metal2 53406 6460 53406 6460 0 _0372_
rlabel metal2 54970 8330 54970 8330 0 _0373_
rlabel metal1 56948 8466 56948 8466 0 _0374_
rlabel metal2 56856 9622 56856 9622 0 _0375_
rlabel metal1 55338 9554 55338 9554 0 _0376_
rlabel metal1 64170 9554 64170 9554 0 _0377_
rlabel metal2 67482 9078 67482 9078 0 _0378_
rlabel metal2 57546 9724 57546 9724 0 _0379_
rlabel metal2 60582 9452 60582 9452 0 _0380_
rlabel metal2 63434 8636 63434 8636 0 _0381_
rlabel metal1 66976 7378 66976 7378 0 _0382_
rlabel metal1 76866 9554 76866 9554 0 _0383_
rlabel metal1 73370 4590 73370 4590 0 _0384_
rlabel metal1 67620 11118 67620 11118 0 _0385_
rlabel metal1 74106 12614 74106 12614 0 _0386_
rlabel metal1 79212 4114 79212 4114 0 _0387_
rlabel metal2 72726 8738 72726 8738 0 _0388_
rlabel metal1 75164 8942 75164 8942 0 _0389_
rlabel metal2 84318 4794 84318 4794 0 _0390_
rlabel metal1 87124 7854 87124 7854 0 _0391_
rlabel metal1 81558 4794 81558 4794 0 _0392_
rlabel metal2 76314 8330 76314 8330 0 _0393_
rlabel metal1 75072 8058 75072 8058 0 _0394_
rlabel metal2 83858 9452 83858 9452 0 _0395_
rlabel metal1 82110 10676 82110 10676 0 _0396_
rlabel metal2 88090 13464 88090 13464 0 _0397_
rlabel metal1 84916 12614 84916 12614 0 _0398_
rlabel metal1 108100 8942 108100 8942 0 _0399_
rlabel metal2 98762 10370 98762 10370 0 _0400_
rlabel metal1 82340 11730 82340 11730 0 _0401_
rlabel metal2 105662 10812 105662 10812 0 _0402_
rlabel metal2 111090 7378 111090 7378 0 _0403_
rlabel metal1 98532 12206 98532 12206 0 _0404_
rlabel metal1 91632 12614 91632 12614 0 _0405_
rlabel metal2 93150 5644 93150 5644 0 _0406_
rlabel metal2 95358 8092 95358 8092 0 _0407_
rlabel metal1 112378 8806 112378 8806 0 _0408_
rlabel metal2 119646 9996 119646 9996 0 _0409_
rlabel metal2 118174 10234 118174 10234 0 _0410_
rlabel metal1 117668 7854 117668 7854 0 _0411_
rlabel metal1 123740 7854 123740 7854 0 _0412_
rlabel metal1 121900 10166 121900 10166 0 _0413_
rlabel metal1 108744 8466 108744 8466 0 _0414_
rlabel metal2 118358 6800 118358 6800 0 _0415_
rlabel metal2 115506 4012 115506 4012 0 _0416_
rlabel metal1 117116 11186 117116 11186 0 _0417_
rlabel metal1 114632 9418 114632 9418 0 _0418_
rlabel via1 133170 2363 133170 2363 0 _0419_
rlabel metal2 125074 4692 125074 4692 0 _0420_
rlabel metal1 128524 10642 128524 10642 0 _0421_
rlabel metal2 114126 8636 114126 8636 0 _0422_
rlabel metal1 128018 11764 128018 11764 0 _0423_
rlabel metal2 130226 2689 130226 2689 0 _0424_
rlabel metal1 113114 5202 113114 5202 0 _0425_
rlabel metal1 132848 7922 132848 7922 0 _0426_
rlabel metal1 130272 5678 130272 5678 0 _0427_
rlabel metal1 132526 11322 132526 11322 0 _0428_
rlabel metal1 132756 3502 132756 3502 0 _0429_
rlabel metal1 131376 2482 131376 2482 0 _0430_
rlabel metal2 127374 10098 127374 10098 0 _0431_
rlabel metal1 127282 5338 127282 5338 0 _0432_
rlabel metal1 131560 3162 131560 3162 0 _0433_
rlabel metal2 120566 11084 120566 11084 0 _0434_
rlabel metal1 119232 4182 119232 4182 0 _0435_
rlabel metal2 127006 9860 127006 9860 0 _0436_
rlabel metal1 127788 7514 127788 7514 0 _0437_
rlabel metal1 122590 7786 122590 7786 0 _0438_
rlabel metal2 118542 6205 118542 6205 0 _0439_
rlabel metal1 126914 10438 126914 10438 0 _0440_
rlabel metal1 131514 7514 131514 7514 0 _0441_
rlabel metal1 155986 10574 155986 10574 0 _0442_
rlabel metal1 156814 2618 156814 2618 0 _0443_
rlabel metal1 155066 2312 155066 2312 0 _0444_
rlabel metal2 159206 8738 159206 8738 0 _0445_
rlabel metal2 157734 5406 157734 5406 0 _0446_
rlabel metal2 150006 14178 150006 14178 0 _0447_
rlabel metal2 157182 8058 157182 8058 0 _0448_
rlabel metal1 157826 11764 157826 11764 0 _0449_
rlabel metal2 158470 8432 158470 8432 0 _0450_
rlabel metal2 158286 4930 158286 4930 0 _0451_
rlabel metal1 146602 10200 146602 10200 0 _0452_
rlabel metal2 118174 5848 118174 5848 0 _0453_
rlabel metal1 157251 9350 157251 9350 0 _0454_
rlabel metal1 154284 6290 154284 6290 0 _0455_
rlabel metal2 130870 7123 130870 7123 0 _0456_
rlabel metal2 148258 10030 148258 10030 0 _0457_
rlabel metal2 156170 6154 156170 6154 0 _0458_
rlabel metal1 152214 8058 152214 8058 0 _0459_
rlabel metal2 147568 2414 147568 2414 0 _0460_
rlabel metal1 152260 3094 152260 3094 0 _0461_
rlabel metal1 141634 8942 141634 8942 0 _0462_
rlabel metal1 140438 2414 140438 2414 0 _0463_
rlabel metal2 118266 5100 118266 5100 0 _0464_
rlabel metal1 118726 2992 118726 2992 0 _0465_
rlabel metal2 118634 4896 118634 4896 0 _0466_
rlabel metal2 120842 6324 120842 6324 0 _0467_
rlabel metal1 122544 6834 122544 6834 0 _0468_
rlabel metal1 156032 3162 156032 3162 0 _0469_
rlabel metal2 156998 5338 156998 5338 0 _0470_
rlabel metal1 156722 6290 156722 6290 0 _0471_
rlabel metal1 155066 11050 155066 11050 0 _0472_
rlabel metal2 157550 6460 157550 6460 0 _0473_
rlabel metal2 157918 8330 157918 8330 0 _0474_
rlabel metal1 131192 8262 131192 8262 0 _0475_
rlabel metal2 152168 12954 152168 12954 0 _0476_
rlabel metal1 150144 3026 150144 3026 0 _0477_
rlabel metal1 117254 9486 117254 9486 0 _0478_
rlabel metal2 125810 8364 125810 8364 0 _0479_
rlabel metal2 135378 7582 135378 7582 0 _0480_
rlabel metal2 140162 6970 140162 6970 0 _0481_
rlabel metal2 157826 6868 157826 6868 0 _0482_
rlabel metal1 156630 3060 156630 3060 0 _0483_
rlabel metal2 158562 7038 158562 7038 0 _0484_
rlabel metal1 155296 4114 155296 4114 0 _0485_
rlabel metal2 132894 6392 132894 6392 0 _0486_
rlabel metal1 156768 4114 156768 4114 0 _0487_
rlabel metal1 156860 4590 156860 4590 0 _0488_
rlabel metal1 147890 7922 147890 7922 0 _0489_
rlabel metal1 157090 5576 157090 5576 0 _0490_
rlabel metal1 158286 12852 158286 12852 0 _0491_
rlabel metal2 157090 4012 157090 4012 0 _0492_
rlabel metal1 158240 6290 158240 6290 0 _0493_
rlabel metal2 144670 6528 144670 6528 0 _0494_
rlabel metal2 141174 11084 141174 11084 0 _0495_
rlabel metal1 151708 6766 151708 6766 0 _0496_
rlabel metal1 157228 2482 157228 2482 0 _0497_
rlabel metal1 149822 8602 149822 8602 0 _0498_
rlabel metal1 157136 6766 157136 6766 0 _0499_
rlabel metal1 152030 12172 152030 12172 0 _0500_
rlabel metal2 157734 9520 157734 9520 0 _0501_
rlabel metal2 153318 11798 153318 11798 0 _0502_
rlabel metal1 150788 3162 150788 3162 0 _0503_
rlabel metal1 139610 6766 139610 6766 0 _0504_
rlabel metal1 139794 4590 139794 4590 0 _0505_
rlabel metal1 155710 4114 155710 4114 0 _0506_
rlabel metal2 154606 3876 154606 3876 0 _0507_
rlabel metal1 117714 8296 117714 8296 0 _0508_
rlabel metal2 156354 4522 156354 4522 0 _0509_
rlabel metal1 158010 12750 158010 12750 0 _0510_
rlabel metal2 157826 9350 157826 9350 0 _0511_
rlabel metal2 153134 4624 153134 4624 0 _0512_
rlabel via2 154698 10013 154698 10013 0 _0513_
rlabel metal1 153778 3026 153778 3026 0 _0514_
rlabel via3 155963 5644 155963 5644 0 _0515_
rlabel metal1 140852 7922 140852 7922 0 _0516_
rlabel metal1 133078 4216 133078 4216 0 _0517_
rlabel metal2 157366 6766 157366 6766 0 _0518_
rlabel via1 155158 3043 155158 3043 0 _0519_
rlabel metal1 151064 6290 151064 6290 0 _0520_
rlabel metal1 153134 6290 153134 6290 0 _0521_
rlabel metal1 151892 5678 151892 5678 0 _0522_
rlabel metal1 154284 9078 154284 9078 0 _0523_
rlabel metal1 156032 2414 156032 2414 0 _0524_
rlabel via2 152858 3723 152858 3723 0 _0525_
rlabel metal1 152214 6766 152214 6766 0 _0526_
rlabel viali 151018 6764 151018 6764 0 _0527_
rlabel metal1 154100 5814 154100 5814 0 _0528_
rlabel metal2 153962 4590 153962 4590 0 _0529_
rlabel metal1 155342 2516 155342 2516 0 _0530_
rlabel metal2 154974 2247 154974 2247 0 _0531_
rlabel metal1 153042 2346 153042 2346 0 _0532_
rlabel metal1 143566 8942 143566 8942 0 _0533_
rlabel metal2 136850 6222 136850 6222 0 _0534_
rlabel metal2 139794 6460 139794 6460 0 _0535_
rlabel metal2 140530 6460 140530 6460 0 _0536_
rlabel metal1 139426 4794 139426 4794 0 _0537_
rlabel metal1 143566 8568 143566 8568 0 _0538_
rlabel metal1 150052 2346 150052 2346 0 _0539_
rlabel metal2 81282 6698 81282 6698 0 clknet_0_sclk
rlabel metal2 21390 7854 21390 7854 0 clknet_1_0__leaf_sclk
rlabel metal1 94070 5644 94070 5644 0 clknet_1_1__leaf_sclk
rlabel metal1 19458 9078 19458 9078 0 clknet_leaf_0_sclk
rlabel metal1 52026 6970 52026 6970 0 clknet_leaf_10_sclk
rlabel metal1 15686 12954 15686 12954 0 clknet_leaf_1_sclk
rlabel metal1 38318 11322 38318 11322 0 clknet_leaf_2_sclk
rlabel metal1 112424 12750 112424 12750 0 clknet_leaf_3_sclk
rlabel metal1 117392 9690 117392 9690 0 clknet_leaf_4_sclk
rlabel metal1 150328 2618 150328 2618 0 clknet_leaf_5_sclk
rlabel metal1 129536 4590 129536 4590 0 clknet_leaf_6_sclk
rlabel metal2 96278 3332 96278 3332 0 clknet_leaf_7_sclk
rlabel metal1 63526 2550 63526 2550 0 clknet_leaf_8_sclk
rlabel metal1 24518 2482 24518 2482 0 clknet_leaf_9_sclk
rlabel metal1 8832 13498 8832 13498 0 dq[0]
rlabel metal1 64906 12410 64906 12410 0 dq[100]
rlabel metal2 65458 14127 65458 14127 0 dq[101]
rlabel metal2 66102 14127 66102 14127 0 dq[102]
rlabel metal1 66240 13498 66240 13498 0 dq[103]
rlabel metal2 67022 14120 67022 14120 0 dq[104]
rlabel metal1 67620 12954 67620 12954 0 dq[105]
rlabel metal1 67896 13498 67896 13498 0 dq[106]
rlabel metal1 68770 12410 68770 12410 0 dq[107]
rlabel metal1 69046 13498 69046 13498 0 dq[108]
rlabel metal1 69920 12410 69920 12410 0 dq[109]
rlabel metal1 13478 13158 13478 13158 0 dq[10]
rlabel metal1 69736 13498 69736 13498 0 dq[110]
rlabel metal2 70886 14392 70886 14392 0 dq[111]
rlabel metal2 71346 14399 71346 14399 0 dq[112]
rlabel metal2 72082 14399 72082 14399 0 dq[113]
rlabel metal1 72680 12954 72680 12954 0 dq[114]
rlabel metal2 72818 14399 72818 14399 0 dq[115]
rlabel metal1 74152 12954 74152 12954 0 dq[116]
rlabel metal2 73922 14399 73922 14399 0 dq[117]
rlabel metal2 74658 14399 74658 14399 0 dq[118]
rlabel metal1 75440 12954 75440 12954 0 dq[119]
rlabel metal1 14628 13498 14628 13498 0 dq[11]
rlabel metal2 75486 14399 75486 14399 0 dq[120]
rlabel metal1 76498 12954 76498 12954 0 dq[121]
rlabel metal1 76590 13498 76590 13498 0 dq[122]
rlabel metal1 77740 12954 77740 12954 0 dq[123]
rlabel metal2 78062 14392 78062 14392 0 dq[124]
rlabel metal2 78798 14127 78798 14127 0 dq[125]
rlabel metal1 79074 13498 79074 13498 0 dq[126]
rlabel metal2 79810 14399 79810 14399 0 dq[127]
rlabel metal1 80362 13498 80362 13498 0 dq[128]
rlabel metal1 81144 13498 81144 13498 0 dq[129]
rlabel metal1 15594 12070 15594 12070 0 dq[12]
rlabel metal1 81742 13430 81742 13430 0 dq[130]
rlabel metal1 82386 13498 82386 13498 0 dq[131]
rlabel metal1 82754 12954 82754 12954 0 dq[132]
rlabel metal1 83490 13498 83490 13498 0 dq[133]
rlabel metal1 83766 12954 83766 12954 0 dq[134]
rlabel metal2 84134 14392 84134 14392 0 dq[135]
rlabel metal1 85054 13498 85054 13498 0 dq[136]
rlabel metal1 85330 12410 85330 12410 0 dq[137]
rlabel metal1 86204 12410 86204 12410 0 dq[138]
rlabel metal1 87354 12954 87354 12954 0 dq[139]
rlabel metal1 16468 12954 16468 12954 0 dq[13]
rlabel metal1 87170 11866 87170 11866 0 dq[140]
rlabel metal1 89102 12920 89102 12920 0 dq[141]
rlabel metal2 87998 13984 87998 13984 0 dq[142]
rlabel metal2 88826 14399 88826 14399 0 dq[143]
rlabel metal2 89148 12444 89148 12444 0 dq[144]
rlabel metal1 90252 12342 90252 12342 0 dq[145]
rlabel metal2 93242 12517 93242 12517 0 dq[146]
rlabel metal1 92644 13498 92644 13498 0 dq[147]
rlabel metal1 93150 13158 93150 13158 0 dq[148]
rlabel metal1 92690 12070 92690 12070 0 dq[149]
rlabel metal2 17526 14127 17526 14127 0 dq[14]
rlabel metal1 93334 12954 93334 12954 0 dq[150]
rlabel metal1 94484 13430 94484 13430 0 dq[151]
rlabel metal1 93886 11594 93886 11594 0 dq[152]
rlabel metal1 96324 13430 96324 13430 0 dq[153]
rlabel metal1 94806 11866 94806 11866 0 dq[154]
rlabel metal1 96370 13498 96370 13498 0 dq[155]
rlabel metal1 97382 12920 97382 12920 0 dq[156]
rlabel metal1 96554 12410 96554 12410 0 dq[157]
rlabel metal1 97750 13430 97750 13430 0 dq[158]
rlabel metal1 97934 12954 97934 12954 0 dq[159]
rlabel metal1 17572 13498 17572 13498 0 dq[15]
rlabel via1 98026 13515 98026 13515 0 dq[160]
rlabel metal2 98486 14358 98486 14358 0 dq[161]
rlabel metal2 99038 14222 99038 14222 0 dq[162]
rlabel metal1 99958 12682 99958 12682 0 dq[163]
rlabel metal1 100556 12954 100556 12954 0 dq[164]
rlabel metal1 101200 12682 101200 12682 0 dq[165]
rlabel metal1 102212 13430 102212 13430 0 dq[166]
rlabel metal1 102120 12954 102120 12954 0 dq[167]
rlabel metal1 102902 12954 102902 12954 0 dq[168]
rlabel metal1 103730 13498 103730 13498 0 dq[169]
rlabel metal1 18216 13498 18216 13498 0 dq[16]
rlabel metal1 104420 13430 104420 13430 0 dq[170]
rlabel metal1 104282 12954 104282 12954 0 dq[171]
rlabel metal1 105478 13498 105478 13498 0 dq[172]
rlabel metal1 105248 12410 105248 12410 0 dq[173]
rlabel metal1 105846 12410 105846 12410 0 dq[174]
rlabel metal1 106950 12614 106950 12614 0 dq[175]
rlabel metal1 106950 12410 106950 12410 0 dq[176]
rlabel metal1 107824 12954 107824 12954 0 dq[177]
rlabel metal1 108606 13464 108606 13464 0 dq[178]
rlabel metal2 108422 14120 108422 14120 0 dq[179]
rlabel metal2 18722 14127 18722 14127 0 dq[17]
rlabel metal2 108974 14392 108974 14392 0 dq[180]
rlabel metal1 110492 13430 110492 13430 0 dq[181]
rlabel metal2 110177 15300 110177 15300 0 dq[182]
rlabel metal1 111458 13498 111458 13498 0 dq[183]
rlabel metal1 112286 13430 112286 13430 0 dq[184]
rlabel metal1 112010 12410 112010 12410 0 dq[185]
rlabel metal1 112608 12954 112608 12954 0 dq[186]
rlabel metal1 113298 13498 113298 13498 0 dq[187]
rlabel metal2 113666 14127 113666 14127 0 dq[188]
rlabel metal1 114448 13498 114448 13498 0 dq[189]
rlabel metal1 19136 13498 19136 13498 0 dq[18]
rlabel metal1 115460 13430 115460 13430 0 dq[190]
rlabel metal2 115145 15300 115145 15300 0 dq[191]
rlabel metal1 117070 13430 117070 13430 0 dq[192]
rlabel metal2 116334 13685 116334 13685 0 dq[193]
rlabel metal1 117438 13498 117438 13498 0 dq[194]
rlabel metal1 117898 13396 117898 13396 0 dq[195]
rlabel metal1 118174 12954 118174 12954 0 dq[196]
rlabel metal2 118358 14392 118358 14392 0 dq[197]
rlabel metal1 119968 13430 119968 13430 0 dq[198]
rlabel metal1 119876 12954 119876 12954 0 dq[199]
rlabel metal1 19780 12954 19780 12954 0 dq[19]
rlabel metal1 9844 12954 9844 12954 0 dq[1]
rlabel metal1 120428 12954 120428 12954 0 dq[200]
rlabel metal1 121026 13498 121026 13498 0 dq[201]
rlabel metal1 121302 12954 121302 12954 0 dq[202]
rlabel metal1 121716 12410 121716 12410 0 dq[203]
rlabel metal1 123326 12614 123326 12614 0 dq[204]
rlabel metal1 123970 13498 123970 13498 0 dq[205]
rlabel metal1 124246 12954 124246 12954 0 dq[206]
rlabel metal2 123878 13853 123878 13853 0 dq[207]
rlabel metal1 125304 13430 125304 13430 0 dq[208]
rlabel metal1 125580 12614 125580 12614 0 dq[209]
rlabel metal2 20601 15300 20601 15300 0 dq[20]
rlabel metal1 126086 13498 126086 13498 0 dq[210]
rlabel metal1 126914 13430 126914 13430 0 dq[211]
rlabel metal1 127834 13464 127834 13464 0 dq[212]
rlabel metal1 127512 12410 127512 12410 0 dq[213]
rlabel metal2 128018 14399 128018 14399 0 dq[214]
rlabel metal2 128294 14120 128294 14120 0 dq[215]
rlabel metal1 129582 13430 129582 13430 0 dq[216]
rlabel metal1 130042 12954 130042 12954 0 dq[217]
rlabel metal1 130502 13498 130502 13498 0 dq[218]
rlabel metal1 130778 12954 130778 12954 0 dq[219]
rlabel metal1 20562 13430 20562 13430 0 dq[21]
rlabel metal1 131468 13498 131468 13498 0 dq[220]
rlabel metal2 131882 14127 131882 14127 0 dq[221]
rlabel metal1 132756 13498 132756 13498 0 dq[222]
rlabel metal1 133216 13430 133216 13430 0 dq[223]
rlabel metal1 134182 13430 134182 13430 0 dq[224]
rlabel metal1 133998 12954 133998 12954 0 dq[225]
rlabel metal1 134918 13498 134918 13498 0 dq[226]
rlabel metal1 135240 12954 135240 12954 0 dq[227]
rlabel metal1 136022 13498 136022 13498 0 dq[228]
rlabel metal1 136712 13498 136712 13498 0 dq[229]
rlabel metal1 21206 13498 21206 13498 0 dq[22]
rlabel metal1 136712 12954 136712 12954 0 dq[230]
rlabel metal2 137126 14392 137126 14392 0 dq[231]
rlabel metal2 137954 14127 137954 14127 0 dq[232]
rlabel metal1 138506 13498 138506 13498 0 dq[233]
rlabel metal1 139242 13498 139242 13498 0 dq[234]
rlabel metal1 139564 12954 139564 12954 0 dq[235]
rlabel metal1 140254 13498 140254 13498 0 dq[236]
rlabel metal1 141082 13498 141082 13498 0 dq[237]
rlabel metal1 141726 13430 141726 13430 0 dq[238]
rlabel metal2 141443 15300 141443 15300 0 dq[239]
rlabel via1 22034 13413 22034 13413 0 dq[23]
rlabel metal1 142554 12954 142554 12954 0 dq[240]
rlabel metal1 140714 12614 140714 12614 0 dq[241]
rlabel metal1 145084 12410 145084 12410 0 dq[242]
rlabel metal2 148350 11968 148350 11968 0 dq[243]
rlabel metal2 144302 14137 144302 14137 0 dq[244]
rlabel metal2 144854 13746 144854 13746 0 dq[245]
rlabel metal2 153594 13634 153594 13634 0 dq[246]
rlabel metal2 154330 14246 154330 14246 0 dq[247]
rlabel metal2 154422 14110 154422 14110 0 dq[248]
rlabel metal1 156032 13498 156032 13498 0 dq[249]
rlabel metal1 22954 12410 22954 12410 0 dq[24]
rlabel metal1 156354 13430 156354 13430 0 dq[250]
rlabel metal2 156170 13362 156170 13362 0 dq[251]
rlabel metal1 155526 12342 155526 12342 0 dq[252]
rlabel metal1 157642 13192 157642 13192 0 dq[253]
rlabel metal1 156860 12954 156860 12954 0 dq[254]
rlabel metal2 150321 15300 150321 15300 0 dq[255]
rlabel metal1 23046 12954 23046 12954 0 dq[25]
rlabel metal1 23184 13498 23184 13498 0 dq[26]
rlabel metal1 24196 12410 24196 12410 0 dq[27]
rlabel metal1 24150 12954 24150 12954 0 dq[28]
rlabel metal1 24196 13430 24196 13430 0 dq[29]
rlabel metal2 10619 15300 10619 15300 0 dq[2]
rlabel metal1 23966 13192 23966 13192 0 dq[30]
rlabel metal2 26450 14127 26450 14127 0 dq[31]
rlabel metal2 27278 13848 27278 13848 0 dq[32]
rlabel metal1 27922 12410 27922 12410 0 dq[33]
rlabel metal1 27876 13498 27876 13498 0 dq[34]
rlabel metal1 28658 13498 28658 13498 0 dq[35]
rlabel metal1 29716 12410 29716 12410 0 dq[36]
rlabel metal2 29854 13957 29854 13957 0 dq[37]
rlabel metal1 29854 13498 29854 13498 0 dq[38]
rlabel metal1 31418 11866 31418 11866 0 dq[39]
rlabel metal2 10074 13702 10074 13702 0 dq[3]
rlabel metal2 31694 13848 31694 13848 0 dq[40]
rlabel metal2 32522 14127 32522 14127 0 dq[41]
rlabel metal2 32798 14392 32798 14392 0 dq[42]
rlabel metal2 33534 14127 33534 14127 0 dq[43]
rlabel metal1 33994 12410 33994 12410 0 dq[44]
rlabel metal1 33948 13498 33948 13498 0 dq[45]
rlabel metal2 35105 15300 35105 15300 0 dq[46]
rlabel metal1 34500 13430 34500 13430 0 dq[47]
rlabel metal1 36248 12410 36248 12410 0 dq[48]
rlabel metal1 36754 12954 36754 12954 0 dq[49]
rlabel metal1 11040 12954 11040 12954 0 dq[4]
rlabel metal1 37306 12410 37306 12410 0 dq[50]
rlabel metal1 37858 12954 37858 12954 0 dq[51]
rlabel metal1 38456 12410 38456 12410 0 dq[52]
rlabel metal1 38732 12954 38732 12954 0 dq[53]
rlabel metal1 38640 13498 38640 13498 0 dq[54]
rlabel metal1 39698 12410 39698 12410 0 dq[55]
rlabel metal2 40671 15300 40671 15300 0 dq[56]
rlabel metal1 38732 13158 38732 13158 0 dq[57]
rlabel metal2 41630 14120 41630 14120 0 dq[58]
rlabel metal1 40802 12648 40802 12648 0 dq[59]
rlabel metal1 11316 13498 11316 13498 0 dq[5]
rlabel metal1 39330 13192 39330 13192 0 dq[60]
rlabel metal1 42596 11866 42596 11866 0 dq[61]
rlabel metal2 43601 15300 43601 15300 0 dq[62]
rlabel metal1 42964 11526 42964 11526 0 dq[63]
rlabel metal1 45034 10778 45034 10778 0 dq[64]
rlabel metal1 42642 13192 42642 13192 0 dq[65]
rlabel metal1 44436 11594 44436 11594 0 dq[66]
rlabel metal1 46368 10234 46368 10234 0 dq[67]
rlabel metal1 43884 12342 43884 12342 0 dq[68]
rlabel metal1 44390 11832 44390 11832 0 dq[69]
rlabel viali 12634 11526 12634 11526 0 dq[6]
rlabel metal1 45908 11866 45908 11866 0 dq[70]
rlabel metal3 46276 12444 46276 12444 0 dq[71]
rlabel metal2 49358 13853 49358 13853 0 dq[72]
rlabel metal1 46828 12614 46828 12614 0 dq[73]
rlabel metal2 50462 13853 50462 13853 0 dq[74]
rlabel metal1 49726 11866 49726 11866 0 dq[75]
rlabel metal2 51421 15300 51421 15300 0 dq[76]
rlabel metal1 52118 11628 52118 11628 0 dq[77]
rlabel metal1 51888 10778 51888 10778 0 dq[78]
rlabel metal2 53321 15300 53321 15300 0 dq[79]
rlabel metal2 13478 13984 13478 13984 0 dq[7]
rlabel metal1 50830 12308 50830 12308 0 dq[80]
rlabel metal2 54326 14120 54326 14120 0 dq[81]
rlabel metal1 52302 12070 52302 12070 0 dq[82]
rlabel metal2 55331 15300 55331 15300 0 dq[83]
rlabel metal2 56127 15300 56127 15300 0 dq[84]
rlabel metal1 56718 9690 56718 9690 0 dq[85]
rlabel metal2 56849 15300 56849 15300 0 dq[86]
rlabel metal1 53866 12614 53866 12614 0 dq[87]
rlabel metal2 58335 15300 58335 15300 0 dq[88]
rlabel metal1 58880 10166 58880 10166 0 dq[89]
rlabel metal1 13846 12410 13846 12410 0 dq[8]
rlabel metal1 58604 11322 58604 11322 0 dq[90]
rlabel metal1 59938 10166 59938 10166 0 dq[91]
rlabel metal2 60451 15300 60451 15300 0 dq[92]
rlabel metal2 60030 11594 60030 11594 0 dq[93]
rlabel metal2 61502 14120 61502 14120 0 dq[94]
rlabel metal1 62330 11322 62330 11322 0 dq[95]
rlabel metal1 63020 11866 63020 11866 0 dq[96]
rlabel metal2 63211 15300 63211 15300 0 dq[97]
rlabel metal2 63763 15300 63763 15300 0 dq[98]
rlabel metal2 63894 14127 63894 14127 0 dq[99]
rlabel metal1 12558 13464 12558 13464 0 dq[9]
rlabel metal2 1610 9775 1610 9775 0 latch
rlabel metal2 13662 10540 13662 10540 0 net1
rlabel metal1 68126 12818 68126 12818 0 net10
rlabel metal1 117392 12614 117392 12614 0 net100
rlabel metal1 114816 12818 114816 12818 0 net101
rlabel metal1 114724 13294 114724 13294 0 net102
rlabel metal1 18906 13260 18906 13260 0 net103
rlabel metal2 112930 13396 112930 13396 0 net104
rlabel metal2 118036 12580 118036 12580 0 net105
rlabel via1 117346 13277 117346 13277 0 net106
rlabel metal2 152674 13668 152674 13668 0 net107
rlabel metal1 152628 11866 152628 11866 0 net108
rlabel metal2 150834 3060 150834 3060 0 net109
rlabel metal1 72634 2618 72634 2618 0 net11
rlabel metal2 152674 10591 152674 10591 0 net110
rlabel metal2 128938 7888 128938 7888 0 net111
rlabel metal3 123648 12988 123648 12988 0 net112
rlabel metal2 130410 13311 130410 13311 0 net113
rlabel metal1 19642 12852 19642 12852 0 net114
rlabel metal1 12926 12818 12926 12818 0 net115
rlabel metal1 130318 4012 130318 4012 0 net116
rlabel metal1 131468 8602 131468 8602 0 net117
rlabel metal1 122544 12886 122544 12886 0 net118
rlabel via2 150834 7531 150834 7531 0 net119
rlabel metal1 73462 12104 73462 12104 0 net12
rlabel metal2 153778 2261 153778 2261 0 net120
rlabel metal2 129582 13532 129582 13532 0 net121
rlabel metal2 128846 12988 128846 12988 0 net122
rlabel metal2 128478 12342 128478 12342 0 net123
rlabel metal2 130042 12461 130042 12461 0 net124
rlabel metal1 126546 12886 126546 12886 0 net125
rlabel metal1 21022 11696 21022 11696 0 net126
rlabel metal2 130686 11577 130686 11577 0 net127
rlabel metal2 131790 11169 131790 11169 0 net128
rlabel metal1 128708 13294 128708 13294 0 net129
rlabel metal2 73738 9928 73738 9928 0 net13
rlabel metal2 127466 8092 127466 8092 0 net130
rlabel metal1 132204 11526 132204 11526 0 net131
rlabel metal1 140760 12954 140760 12954 0 net132
rlabel via2 140806 6613 140806 6613 0 net133
rlabel metal1 131698 12410 131698 12410 0 net134
rlabel metal1 132388 13294 132388 13294 0 net135
rlabel metal1 133078 12852 133078 12852 0 net136
rlabel metal1 19826 13294 19826 13294 0 net137
rlabel metal2 132020 13294 132020 13294 0 net138
rlabel metal1 131146 12750 131146 12750 0 net139
rlabel metal2 67942 9452 67942 9452 0 net14
rlabel metal1 123878 13328 123878 13328 0 net140
rlabel metal1 129766 12716 129766 12716 0 net141
rlabel metal1 134090 13294 134090 13294 0 net142
rlabel metal1 119048 12818 119048 12818 0 net143
rlabel metal2 135562 10795 135562 10795 0 net144
rlabel metal1 129858 12648 129858 12648 0 net145
rlabel metal1 135976 11050 135976 11050 0 net146
rlabel metal1 129214 12784 129214 12784 0 net147
rlabel metal1 20424 13294 20424 13294 0 net148
rlabel metal2 136666 12631 136666 12631 0 net149
rlabel metal2 7866 13600 7866 13600 0 net15
rlabel metal2 113574 2720 113574 2720 0 net150
rlabel metal1 137586 10234 137586 10234 0 net151
rlabel via2 116150 12597 116150 12597 0 net152
rlabel metal2 139426 8636 139426 8636 0 net153
rlabel metal1 130318 10744 130318 10744 0 net154
rlabel metal1 137402 10472 137402 10472 0 net155
rlabel metal1 136850 9656 136850 9656 0 net156
rlabel metal2 134734 6545 134734 6545 0 net157
rlabel metal2 117990 13022 117990 13022 0 net158
rlabel metal2 21574 13294 21574 13294 0 net159
rlabel metal2 77786 12342 77786 12342 0 net16
rlabel metal2 135562 12784 135562 12784 0 net160
rlabel via2 150834 12699 150834 12699 0 net161
rlabel metal1 152398 12342 152398 12342 0 net162
rlabel metal1 133216 9690 133216 9690 0 net163
rlabel metal3 135884 2652 135884 2652 0 net164
rlabel via2 131146 9061 131146 9061 0 net165
rlabel metal2 153410 13804 153410 13804 0 net166
rlabel metal1 149776 3706 149776 3706 0 net167
rlabel metal2 154882 13838 154882 13838 0 net168
rlabel metal2 155986 13668 155986 13668 0 net169
rlabel metal1 70794 13294 70794 13294 0 net17
rlabel metal1 31878 8296 31878 8296 0 net170
rlabel metal2 156722 13940 156722 13940 0 net171
rlabel metal2 156078 13498 156078 13498 0 net172
rlabel metal1 153180 11526 153180 11526 0 net173
rlabel metal2 157458 14008 157458 14008 0 net174
rlabel via2 156722 12835 156722 12835 0 net175
rlabel metal1 154974 12410 154974 12410 0 net176
rlabel metal1 37996 6630 37996 6630 0 net177
rlabel metal1 22586 13328 22586 13328 0 net178
rlabel metal1 31418 10540 31418 10540 0 net179
rlabel metal1 71622 13294 71622 13294 0 net18
rlabel metal1 22724 12750 22724 12750 0 net180
rlabel metal1 32338 7412 32338 7412 0 net181
rlabel metal2 10350 9197 10350 9197 0 net182
rlabel metal2 23782 12954 23782 12954 0 net183
rlabel metal1 35144 10778 35144 10778 0 net184
rlabel metal1 25806 10438 25806 10438 0 net185
rlabel metal1 40526 2822 40526 2822 0 net186
rlabel metal1 27508 13294 27508 13294 0 net187
rlabel metal1 19366 11866 19366 11866 0 net188
rlabel metal1 18814 10710 18814 10710 0 net189
rlabel metal2 75762 12954 75762 12954 0 net19
rlabel metal1 26634 12682 26634 12682 0 net190
rlabel metal1 19688 3706 19688 3706 0 net191
rlabel metal1 29486 9078 29486 9078 0 net192
rlabel metal1 19734 2618 19734 2618 0 net193
rlabel metal1 32522 12138 32522 12138 0 net194
rlabel metal2 27692 12988 27692 12988 0 net195
rlabel metal1 32568 3638 32568 3638 0 net196
rlabel metal1 33764 12070 33764 12070 0 net197
rlabel metal1 40342 12240 40342 12240 0 net198
rlabel metal1 33626 13328 33626 13328 0 net199
rlabel metal1 6992 2346 6992 2346 0 net2
rlabel metal1 73600 12750 73600 12750 0 net20
rlabel metal1 36938 12750 36938 12750 0 net200
rlabel metal1 34592 13294 34592 13294 0 net201
rlabel metal1 34638 11322 34638 11322 0 net202
rlabel metal1 34086 12716 34086 12716 0 net203
rlabel metal2 19550 4352 19550 4352 0 net204
rlabel metal1 37904 12206 37904 12206 0 net205
rlabel metal1 37260 12818 37260 12818 0 net206
rlabel metal1 36984 12682 36984 12682 0 net207
rlabel metal2 39882 13124 39882 13124 0 net208
rlabel metal1 38042 13362 38042 13362 0 net209
rlabel metal1 73462 13294 73462 13294 0 net21
rlabel metal2 39238 11866 39238 11866 0 net210
rlabel metal2 41446 10676 41446 10676 0 net211
rlabel metal2 38778 12857 38778 12857 0 net212
rlabel metal2 35466 13022 35466 13022 0 net213
rlabel metal3 40572 12308 40572 12308 0 net214
rlabel metal1 16790 7752 16790 7752 0 net215
rlabel metal1 39606 11866 39606 11866 0 net216
rlabel metal1 44436 13158 44436 13158 0 net217
rlabel metal2 49450 8840 49450 8840 0 net218
rlabel metal1 42458 11730 42458 11730 0 net219
rlabel metal2 74842 12699 74842 12699 0 net22
rlabel metal2 47886 10200 47886 10200 0 net220
rlabel metal1 41262 13328 41262 13328 0 net221
rlabel metal2 42826 9894 42826 9894 0 net222
rlabel metal1 46782 10098 46782 10098 0 net223
rlabel metal1 32982 11288 32982 11288 0 net224
rlabel metal1 35742 9010 35742 9010 0 net225
rlabel metal1 13524 12614 13524 12614 0 net226
rlabel metal2 56810 4624 56810 4624 0 net227
rlabel metal1 40388 10234 40388 10234 0 net228
rlabel metal1 58742 9350 58742 9350 0 net229
rlabel metal2 79994 13311 79994 13311 0 net23
rlabel metal1 53544 11322 53544 11322 0 net230
rlabel metal2 73186 4250 73186 4250 0 net231
rlabel metal1 48898 11730 48898 11730 0 net232
rlabel metal2 51198 9690 51198 9690 0 net233
rlabel metal1 50186 7990 50186 7990 0 net234
rlabel metal1 50370 3706 50370 3706 0 net235
rlabel via1 53866 8942 53866 8942 0 net236
rlabel metal2 32430 2176 32430 2176 0 net237
rlabel metal1 54317 6154 54317 6154 0 net238
rlabel metal2 66286 3536 66286 3536 0 net239
rlabel metal1 74980 13294 74980 13294 0 net24
rlabel metal2 51658 12410 51658 12410 0 net240
rlabel metal2 53590 11220 53590 11220 0 net241
rlabel metal1 54694 5338 54694 5338 0 net242
rlabel metal2 46966 13226 46966 13226 0 net243
rlabel metal2 54326 12036 54326 12036 0 net244
rlabel metal1 55936 12954 55936 12954 0 net245
rlabel metal1 55430 13430 55430 13430 0 net246
rlabel metal2 58834 10642 58834 10642 0 net247
rlabel metal1 13524 12206 13524 12206 0 net248
rlabel metal1 57638 10778 57638 10778 0 net249
rlabel metal1 75213 12750 75213 12750 0 net25
rlabel metal1 59846 10064 59846 10064 0 net250
rlabel metal2 60122 11662 60122 11662 0 net251
rlabel metal1 59846 11152 59846 11152 0 net252
rlabel metal1 58742 12784 58742 12784 0 net253
rlabel metal1 62744 12614 62744 12614 0 net254
rlabel metal1 59570 12648 59570 12648 0 net255
rlabel metal2 62514 11356 62514 11356 0 net256
rlabel metal1 62238 12104 62238 12104 0 net257
rlabel metal1 64262 12818 64262 12818 0 net258
rlabel metal2 17066 5814 17066 5814 0 net259
rlabel metal1 21850 13430 21850 13430 0 net26
rlabel metal2 116978 13044 116978 13044 0 net260
rlabel metal1 18538 2618 18538 2618 0 net261
rlabel metal1 28980 12818 28980 12818 0 net262
rlabel metal1 30130 5134 30130 5134 0 net263
rlabel metal1 34178 12682 34178 12682 0 net264
rlabel metal1 38042 6834 38042 6834 0 net265
rlabel metal1 42504 12614 42504 12614 0 net266
rlabel metal1 42136 8942 42136 8942 0 net267
rlabel metal1 21666 11050 21666 11050 0 net268
rlabel metal1 55522 8466 55522 8466 0 net269
rlabel metal1 75348 13294 75348 13294 0 net27
rlabel metal1 53866 12818 53866 12818 0 net270
rlabel metal1 52946 10540 52946 10540 0 net271
rlabel metal2 57270 12036 57270 12036 0 net272
rlabel metal1 58190 12376 58190 12376 0 net273
rlabel metal1 74658 2414 74658 2414 0 net274
rlabel metal2 76222 11526 76222 11526 0 net275
rlabel metal1 80822 12750 80822 12750 0 net276
rlabel metal1 54740 9146 54740 9146 0 net277
rlabel metal1 90804 11662 90804 11662 0 net278
rlabel metal1 88964 13294 88964 13294 0 net279
rlabel metal1 84640 3638 84640 3638 0 net28
rlabel metal1 95496 12818 95496 12818 0 net280
rlabel metal1 116472 13158 116472 13158 0 net281
rlabel metal1 110308 11118 110308 11118 0 net282
rlabel metal1 129030 7990 129030 7990 0 net283
rlabel metal1 121762 11118 121762 11118 0 net284
rlabel metal1 136022 9962 136022 9962 0 net285
rlabel metal2 133170 11696 133170 11696 0 net286
rlabel metal1 136390 10438 136390 10438 0 net287
rlabel metal1 152306 3570 152306 3570 0 net288
rlabel metal1 154054 12852 154054 12852 0 net289
rlabel metal1 76774 13294 76774 13294 0 net29
rlabel metal1 155342 9962 155342 9962 0 net290
rlabel via1 132802 6222 132802 6222 0 net291
rlabel metal1 115736 13294 115736 13294 0 net292
rlabel metal2 9338 8398 9338 8398 0 net3
rlabel metal1 81282 12920 81282 12920 0 net30
rlabel metal1 76452 13226 76452 13226 0 net31
rlabel metal1 79074 11866 79074 11866 0 net32
rlabel metal1 83490 6154 83490 6154 0 net33
rlabel metal1 72266 12920 72266 12920 0 net34
rlabel metal1 80868 13294 80868 13294 0 net35
rlabel metal1 81236 13294 81236 13294 0 net36
rlabel metal1 18860 4590 18860 4590 0 net37
rlabel metal1 83076 9418 83076 9418 0 net38
rlabel metal1 83030 13328 83030 13328 0 net39
rlabel metal1 9522 13260 9522 13260 0 net4
rlabel metal2 83214 13124 83214 13124 0 net40
rlabel metal1 84226 13294 84226 13294 0 net41
rlabel metal1 91172 7990 91172 7990 0 net42
rlabel metal1 88090 13498 88090 13498 0 net43
rlabel metal1 86986 13294 86986 13294 0 net44
rlabel metal2 82110 13226 82110 13226 0 net45
rlabel metal1 85928 11866 85928 11866 0 net46
rlabel metal2 87906 13260 87906 13260 0 net47
rlabel metal1 22080 7242 22080 7242 0 net48
rlabel metal1 75026 10200 75026 10200 0 net49
rlabel metal2 65826 11356 65826 11356 0 net5
rlabel metal1 89286 12784 89286 12784 0 net50
rlabel metal1 89562 12818 89562 12818 0 net51
rlabel metal2 90850 13498 90850 13498 0 net52
rlabel metal1 83536 12138 83536 12138 0 net53
rlabel metal1 87998 9146 87998 9146 0 net54
rlabel metal2 93426 12767 93426 12767 0 net55
rlabel metal1 96968 11730 96968 11730 0 net56
rlabel metal2 109618 12512 109618 12512 0 net57
rlabel metal2 70610 11424 70610 11424 0 net58
rlabel metal1 20194 12648 20194 12648 0 net59
rlabel metal1 64676 12682 64676 12682 0 net6
rlabel metal1 94392 9622 94392 9622 0 net60
rlabel metal2 95910 13345 95910 13345 0 net61
rlabel metal1 96002 9078 96002 9078 0 net62
rlabel via2 97014 13277 97014 13277 0 net63
rlabel metal1 96278 11254 96278 11254 0 net64
rlabel metal2 97750 13209 97750 13209 0 net65
rlabel metal1 97566 12784 97566 12784 0 net66
rlabel metal2 97014 12444 97014 12444 0 net67
rlabel metal1 96876 12682 96876 12682 0 net68
rlabel metal1 94852 12682 94852 12682 0 net69
rlabel metal1 71898 12648 71898 12648 0 net7
rlabel metal2 17434 13498 17434 13498 0 net70
rlabel metal1 79626 10472 79626 10472 0 net71
rlabel via1 98486 7803 98486 7803 0 net72
rlabel metal1 110078 12376 110078 12376 0 net73
rlabel metal1 99958 7990 99958 7990 0 net74
rlabel metal1 101246 12818 101246 12818 0 net75
rlabel metal2 133170 12801 133170 12801 0 net76
rlabel metal2 104098 13090 104098 13090 0 net77
rlabel metal1 116058 6324 116058 6324 0 net78
rlabel metal1 116150 6392 116150 6392 0 net79
rlabel metal1 65826 13396 65826 13396 0 net8
rlabel metal1 97106 6120 97106 6120 0 net80
rlabel metal1 18400 13294 18400 13294 0 net81
rlabel metal2 109710 13498 109710 13498 0 net82
rlabel metal2 96922 7412 96922 7412 0 net83
rlabel metal1 93518 12682 93518 12682 0 net84
rlabel metal1 101982 3706 101982 3706 0 net85
rlabel metal1 113850 11696 113850 11696 0 net86
rlabel metal1 107962 12818 107962 12818 0 net87
rlabel metal1 111182 11560 111182 11560 0 net88
rlabel metal1 114678 3706 114678 3706 0 net89
rlabel metal2 76130 3264 76130 3264 0 net9
rlabel metal1 109986 13294 109986 13294 0 net90
rlabel metal1 113298 12750 113298 12750 0 net91
rlabel metal1 19688 12750 19688 12750 0 net92
rlabel metal1 112194 13158 112194 13158 0 net93
rlabel metal1 112976 12614 112976 12614 0 net94
rlabel metal1 114218 12070 114218 12070 0 net95
rlabel metal1 112838 13226 112838 13226 0 net96
rlabel metal1 111734 13362 111734 13362 0 net97
rlabel metal1 113666 12206 113666 12206 0 net98
rlabel metal1 115736 12954 115736 12954 0 net99
rlabel metal2 1702 2193 1702 2193 0 rst_n
rlabel via2 4094 13821 4094 13821 0 sclk
rlabel metal2 1610 6103 1610 6103 0 sdi
rlabel metal2 158286 8143 158286 8143 0 sdo
rlabel metal1 25448 12818 25448 12818 0 sr\[0\]
rlabel metal1 72542 10676 72542 10676 0 sr\[100\]
rlabel metal2 73738 7820 73738 7820 0 sr\[101\]
rlabel metal2 72358 8840 72358 8840 0 sr\[102\]
rlabel metal1 57806 13226 57806 13226 0 sr\[103\]
rlabel metal1 73232 5610 73232 5610 0 sr\[104\]
rlabel metal1 73830 10064 73830 10064 0 sr\[105\]
rlabel metal1 75409 2346 75409 2346 0 sr\[106\]
rlabel via1 87910 8534 87910 8534 0 sr\[107\]
rlabel metal2 91954 5576 91954 5576 0 sr\[108\]
rlabel metal1 74750 5542 74750 5542 0 sr\[109\]
rlabel metal1 19228 3910 19228 3910 0 sr\[10\]
rlabel metal1 75118 7854 75118 7854 0 sr\[110\]
rlabel metal2 84318 9078 84318 9078 0 sr\[111\]
rlabel via1 93697 8874 93697 8874 0 sr\[112\]
rlabel metal1 84916 12818 84916 12818 0 sr\[113\]
rlabel metal1 104052 8466 104052 8466 0 sr\[114\]
rlabel metal2 94530 5066 94530 5066 0 sr\[115\]
rlabel metal2 89930 11968 89930 11968 0 sr\[116\]
rlabel metal1 93794 11832 93794 11832 0 sr\[117\]
rlabel via1 93886 5797 93886 5797 0 sr\[118\]
rlabel metal1 76554 6290 76554 6290 0 sr\[119\]
rlabel metal1 17388 8466 17388 8466 0 sr\[11\]
rlabel metal1 89194 12886 89194 12886 0 sr\[120\]
rlabel metal1 92690 6290 92690 6290 0 sr\[121\]
rlabel metal2 94346 9554 94346 9554 0 sr\[122\]
rlabel metal2 89010 12937 89010 12937 0 sr\[123\]
rlabel metal2 74750 9809 74750 9809 0 sr\[124\]
rlabel metal1 96186 12342 96186 12342 0 sr\[125\]
rlabel metal1 87783 6358 87783 6358 0 sr\[126\]
rlabel metal1 71755 12818 71755 12818 0 sr\[127\]
rlabel metal2 79166 11152 79166 11152 0 sr\[128\]
rlabel metal1 70973 6358 70973 6358 0 sr\[129\]
rlabel metal2 16974 5780 16974 5780 0 sr\[12\]
rlabel metal1 95717 9520 95717 9520 0 sr\[130\]
rlabel metal1 56248 12818 56248 12818 0 sr\[131\]
rlabel metal2 88642 13328 88642 13328 0 sr\[132\]
rlabel metal1 115460 9350 115460 9350 0 sr\[133\]
rlabel metal1 95910 7990 95910 7990 0 sr\[134\]
rlabel metal1 90865 11050 90865 11050 0 sr\[135\]
rlabel metal2 99038 7684 99038 7684 0 sr\[136\]
rlabel via2 129582 2499 129582 2499 0 sr\[137\]
rlabel metal1 91402 5032 91402 5032 0 sr\[138\]
rlabel metal2 73002 11305 73002 11305 0 sr\[139\]
rlabel metal1 21344 3706 21344 3706 0 sr\[13\]
rlabel metal2 70518 10387 70518 10387 0 sr\[140\]
rlabel metal2 74842 3689 74842 3689 0 sr\[141\]
rlabel metal1 90574 7990 90574 7990 0 sr\[142\]
rlabel metal2 96830 11509 96830 11509 0 sr\[143\]
rlabel via1 81369 12818 81369 12818 0 sr\[144\]
rlabel metal2 93242 8160 93242 8160 0 sr\[145\]
rlabel metal2 92874 10693 92874 10693 0 sr\[146\]
rlabel metal1 74934 5236 74934 5236 0 sr\[147\]
rlabel metal1 111243 11050 111243 11050 0 sr\[148\]
rlabel metal1 75026 11866 75026 11866 0 sr\[149\]
rlabel metal1 15732 6698 15732 6698 0 sr\[14\]
rlabel metal1 94162 9350 94162 9350 0 sr\[150\]
rlabel metal2 59570 9894 59570 9894 0 sr\[151\]
rlabel metal2 98210 6630 98210 6630 0 sr\[152\]
rlabel metal2 154330 2533 154330 2533 0 sr\[153\]
rlabel metal1 146924 6970 146924 6970 0 sr\[154\]
rlabel metal1 150098 2890 150098 2890 0 sr\[155\]
rlabel metal2 155526 7276 155526 7276 0 sr\[156\]
rlabel metal4 151892 4692 151892 4692 0 sr\[157\]
rlabel metal1 97980 12886 97980 12886 0 sr\[158\]
rlabel metal2 92782 9945 92782 9945 0 sr\[159\]
rlabel metal2 17250 10115 17250 10115 0 sr\[15\]
rlabel metal2 77878 9741 77878 9741 0 sr\[160\]
rlabel metal2 93518 5117 93518 5117 0 sr\[161\]
rlabel metal3 153755 7004 153755 7004 0 sr\[162\]
rlabel metal1 98946 7752 98946 7752 0 sr\[163\]
rlabel metal2 131054 4590 131054 4590 0 sr\[164\]
rlabel metal1 148994 8330 148994 8330 0 sr\[165\]
rlabel metal2 129398 11458 129398 11458 0 sr\[166\]
rlabel metal1 117714 5848 117714 5848 0 sr\[167\]
rlabel metal1 132480 6698 132480 6698 0 sr\[168\]
rlabel via2 91494 6307 91494 6307 0 sr\[169\]
rlabel metal1 20286 6188 20286 6188 0 sr\[16\]
rlabel metal2 128938 4607 128938 4607 0 sr\[170\]
rlabel metal1 94530 3128 94530 3128 0 sr\[171\]
rlabel metal2 117438 2329 117438 2329 0 sr\[172\]
rlabel metal1 106766 3978 106766 3978 0 sr\[173\]
rlabel metal2 118450 5780 118450 5780 0 sr\[174\]
rlabel metal1 119186 5610 119186 5610 0 sr\[175\]
rlabel metal1 118082 11662 118082 11662 0 sr\[176\]
rlabel metal1 116763 3434 116763 3434 0 sr\[177\]
rlabel metal1 154688 7854 154688 7854 0 sr\[178\]
rlabel metal1 152214 9928 152214 9928 0 sr\[179\]
rlabel via1 21661 4522 21661 4522 0 sr\[17\]
rlabel metal2 153502 11679 153502 11679 0 sr\[180\]
rlabel metal4 148028 8636 148028 8636 0 sr\[181\]
rlabel metal1 129720 5338 129720 5338 0 sr\[182\]
rlabel metal2 128386 8415 128386 8415 0 sr\[183\]
rlabel metal2 110078 5338 110078 5338 0 sr\[184\]
rlabel via1 127921 5678 127921 5678 0 sr\[185\]
rlabel metal2 125626 10846 125626 10846 0 sr\[186\]
rlabel metal1 121030 3434 121030 3434 0 sr\[187\]
rlabel metal1 136022 2278 136022 2278 0 sr\[188\]
rlabel via1 115878 6290 115878 6290 0 sr\[189\]
rlabel metal1 25070 5338 25070 5338 0 sr\[18\]
rlabel metal1 129168 5338 129168 5338 0 sr\[190\]
rlabel metal1 151804 10642 151804 10642 0 sr\[191\]
rlabel metal1 153732 4590 153732 4590 0 sr\[192\]
rlabel metal1 153732 13158 153732 13158 0 sr\[193\]
rlabel metal1 147016 5882 147016 5882 0 sr\[194\]
rlabel metal1 146234 4454 146234 4454 0 sr\[195\]
rlabel metal1 153184 10642 153184 10642 0 sr\[196\]
rlabel metal2 155618 5134 155618 5134 0 sr\[197\]
rlabel metal1 150746 9962 150746 9962 0 sr\[198\]
rlabel metal1 154698 12784 154698 12784 0 sr\[199\]
rlabel metal2 28566 10370 28566 10370 0 sr\[19\]
rlabel metal1 18446 10608 18446 10608 0 sr\[1\]
rlabel metal1 135562 4012 135562 4012 0 sr\[200\]
rlabel metal2 135378 10302 135378 10302 0 sr\[201\]
rlabel metal1 132664 6766 132664 6766 0 sr\[202\]
rlabel metal1 150746 7446 150746 7446 0 sr\[203\]
rlabel metal2 156170 9299 156170 9299 0 sr\[204\]
rlabel metal1 155342 12206 155342 12206 0 sr\[205\]
rlabel metal2 155710 12925 155710 12925 0 sr\[206\]
rlabel viali 152218 11050 152218 11050 0 sr\[207\]
rlabel metal1 144394 8976 144394 8976 0 sr\[208\]
rlabel metal2 130870 8160 130870 8160 0 sr\[209\]
rlabel metal2 23414 8840 23414 8840 0 sr\[20\]
rlabel metal2 147706 6817 147706 6817 0 sr\[210\]
rlabel metal2 147890 3621 147890 3621 0 sr\[211\]
rlabel via2 145498 3077 145498 3077 0 sr\[212\]
rlabel metal1 155066 6324 155066 6324 0 sr\[213\]
rlabel metal1 155296 4590 155296 4590 0 sr\[214\]
rlabel metal2 142554 13158 142554 13158 0 sr\[215\]
rlabel metal2 143106 6086 143106 6086 0 sr\[216\]
rlabel metal1 145268 7242 145268 7242 0 sr\[217\]
rlabel metal2 154698 4437 154698 4437 0 sr\[218\]
rlabel metal2 136942 3196 136942 3196 0 sr\[219\]
rlabel metal1 36666 5678 36666 5678 0 sr\[21\]
rlabel metal1 136620 7446 136620 7446 0 sr\[220\]
rlabel metal1 130410 4488 130410 4488 0 sr\[221\]
rlabel via2 156998 8483 156998 8483 0 sr\[222\]
rlabel metal1 131284 7990 131284 7990 0 sr\[223\]
rlabel metal1 132066 5066 132066 5066 0 sr\[224\]
rlabel metal2 118358 9656 118358 9656 0 sr\[225\]
rlabel metal1 131606 6222 131606 6222 0 sr\[226\]
rlabel metal2 149638 2193 149638 2193 0 sr\[227\]
rlabel metal2 123878 2108 123878 2108 0 sr\[228\]
rlabel metal2 135332 5882 135332 5882 0 sr\[229\]
rlabel metal1 38134 9112 38134 9112 0 sr\[22\]
rlabel metal1 128754 9384 128754 9384 0 sr\[230\]
rlabel metal4 147844 7004 147844 7004 0 sr\[231\]
rlabel metal2 136114 2179 136114 2179 0 sr\[232\]
rlabel metal2 156078 9129 156078 9129 0 sr\[233\]
rlabel metal2 155158 2040 155158 2040 0 sr\[234\]
rlabel metal2 134090 9758 134090 9758 0 sr\[235\]
rlabel metal1 142278 7242 142278 7242 0 sr\[236\]
rlabel via1 122134 10642 122134 10642 0 sr\[237\]
rlabel metal1 137862 2414 137862 2414 0 sr\[238\]
rlabel metal2 133262 11356 133262 11356 0 sr\[239\]
rlabel metal1 6026 2482 6026 2482 0 sr\[23\]
rlabel metal1 136528 12274 136528 12274 0 sr\[240\]
rlabel metal2 147062 11526 147062 11526 0 sr\[241\]
rlabel metal2 129582 6868 129582 6868 0 sr\[242\]
rlabel metal2 129490 5525 129490 5525 0 sr\[243\]
rlabel metal2 118174 4590 118174 4590 0 sr\[244\]
rlabel metal1 106536 11118 106536 11118 0 sr\[245\]
rlabel metal1 114816 6766 114816 6766 0 sr\[246\]
rlabel metal1 113528 2414 113528 2414 0 sr\[247\]
rlabel metal1 112838 10438 112838 10438 0 sr\[248\]
rlabel metal1 97934 8908 97934 8908 0 sr\[249\]
rlabel metal1 32706 8398 32706 8398 0 sr\[24\]
rlabel metal1 113850 11050 113850 11050 0 sr\[250\]
rlabel metal1 111044 11866 111044 11866 0 sr\[251\]
rlabel metal1 98486 6188 98486 6188 0 sr\[252\]
rlabel metal2 98394 10268 98394 10268 0 sr\[253\]
rlabel metal1 98486 7888 98486 7888 0 sr\[254\]
rlabel metal1 17158 7922 17158 7922 0 sr\[25\]
rlabel metal1 21666 12376 21666 12376 0 sr\[26\]
rlabel metal2 5198 10030 5198 10030 0 sr\[27\]
rlabel metal1 11592 2414 11592 2414 0 sr\[28\]
rlabel metal2 20286 11288 20286 11288 0 sr\[29\]
rlabel metal1 18584 8602 18584 8602 0 sr\[2\]
rlabel metal1 49634 2618 49634 2618 0 sr\[30\]
rlabel metal2 12466 11424 12466 11424 0 sr\[31\]
rlabel metal1 16468 9418 16468 9418 0 sr\[32\]
rlabel metal1 16606 2958 16606 2958 0 sr\[33\]
rlabel metal2 15226 3400 15226 3400 0 sr\[34\]
rlabel metal1 16176 11798 16176 11798 0 sr\[35\]
rlabel metal1 17326 10710 17326 10710 0 sr\[36\]
rlabel metal2 11454 6052 11454 6052 0 sr\[37\]
rlabel metal1 17986 8976 17986 8976 0 sr\[38\]
rlabel metal2 20286 5916 20286 5916 0 sr\[39\]
rlabel metal1 21032 2414 21032 2414 0 sr\[3\]
rlabel metal1 13478 11798 13478 11798 0 sr\[40\]
rlabel metal1 16514 10166 16514 10166 0 sr\[41\]
rlabel metal1 19136 7174 19136 7174 0 sr\[42\]
rlabel metal2 54142 8126 54142 8126 0 sr\[43\]
rlabel metal1 48948 13226 48948 13226 0 sr\[44\]
rlabel metal2 36202 13498 36202 13498 0 sr\[45\]
rlabel metal2 39790 8857 39790 8857 0 sr\[46\]
rlabel metal1 54238 8534 54238 8534 0 sr\[47\]
rlabel metal1 40710 11764 40710 11764 0 sr\[48\]
rlabel metal1 31786 11152 31786 11152 0 sr\[49\]
rlabel metal1 16054 8364 16054 8364 0 sr\[4\]
rlabel metal1 45908 2482 45908 2482 0 sr\[50\]
rlabel metal2 37582 10234 37582 10234 0 sr\[51\]
rlabel metal1 34300 12886 34300 12886 0 sr\[52\]
rlabel metal2 35374 6256 35374 6256 0 sr\[53\]
rlabel metal1 33856 6766 33856 6766 0 sr\[54\]
rlabel metal1 40480 6154 40480 6154 0 sr\[55\]
rlabel metal1 40434 8330 40434 8330 0 sr\[56\]
rlabel metal2 32982 5440 32982 5440 0 sr\[57\]
rlabel metal1 27922 13430 27922 13430 0 sr\[58\]
rlabel metal1 33396 3026 33396 3026 0 sr\[59\]
rlabel metal1 15364 12886 15364 12886 0 sr\[5\]
rlabel metal1 35190 11696 35190 11696 0 sr\[60\]
rlabel metal1 36708 13158 36708 13158 0 sr\[61\]
rlabel metal2 33902 10064 33902 10064 0 sr\[62\]
rlabel metal1 40296 13294 40296 13294 0 sr\[63\]
rlabel metal1 54602 13430 54602 13430 0 sr\[64\]
rlabel metal1 44436 6766 44436 6766 0 sr\[65\]
rlabel metal1 43143 7854 43143 7854 0 sr\[66\]
rlabel via1 60586 12818 60586 12818 0 sr\[67\]
rlabel metal2 36570 9996 36570 9996 0 sr\[68\]
rlabel metal1 32430 6222 32430 6222 0 sr\[69\]
rlabel metal1 14172 12886 14172 12886 0 sr\[6\]
rlabel metal1 47794 9078 47794 9078 0 sr\[70\]
rlabel metal1 50876 6086 50876 6086 0 sr\[71\]
rlabel metal2 60030 9078 60030 9078 0 sr\[72\]
rlabel metal1 53866 11016 53866 11016 0 sr\[73\]
rlabel metal2 58650 11169 58650 11169 0 sr\[74\]
rlabel metal1 48525 12818 48525 12818 0 sr\[75\]
rlabel metal1 41998 9418 41998 9418 0 sr\[76\]
rlabel viali 51014 11119 51014 11119 0 sr\[77\]
rlabel metal2 51750 5389 51750 5389 0 sr\[78\]
rlabel metal1 65458 2550 65458 2550 0 sr\[79\]
rlabel metal2 31786 2142 31786 2142 0 sr\[7\]
rlabel metal2 60490 5304 60490 5304 0 sr\[80\]
rlabel metal1 57408 3366 57408 3366 0 sr\[81\]
rlabel metal1 51662 12818 51662 12818 0 sr\[82\]
rlabel metal1 56856 12206 56856 12206 0 sr\[83\]
rlabel metal2 58834 6596 58834 6596 0 sr\[84\]
rlabel metal2 52026 11084 52026 11084 0 sr\[85\]
rlabel metal2 47334 11628 47334 11628 0 sr\[86\]
rlabel metal2 60674 9180 60674 9180 0 sr\[87\]
rlabel metal1 54137 13226 54137 13226 0 sr\[88\]
rlabel metal1 52297 11050 52297 11050 0 sr\[89\]
rlabel metal2 21482 6528 21482 6528 0 sr\[8\]
rlabel metal1 55108 6834 55108 6834 0 sr\[90\]
rlabel metal2 54050 10914 54050 10914 0 sr\[91\]
rlabel metal1 56534 8840 56534 8840 0 sr\[92\]
rlabel metal2 55706 11492 55706 11492 0 sr\[93\]
rlabel metal1 59984 2618 59984 2618 0 sr\[94\]
rlabel metal1 63158 12716 63158 12716 0 sr\[95\]
rlabel metal2 61226 8840 61226 8840 0 sr\[96\]
rlabel metal1 60306 11730 60306 11730 0 sr\[97\]
rlabel metal1 63250 10064 63250 10064 0 sr\[98\]
rlabel metal1 66842 9962 66842 9962 0 sr\[99\]
rlabel metal1 16192 6154 16192 6154 0 sr\[9\]
<< properties >>
string FIXED_BBOX 0 0 160000 16000
<< end >>
