magic
tech sky130A
magscale 1 2
timestamp 1672297736
<< locali >>
rect 2700 -3420 2820 -3400
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
<< viali >>
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
<< metal1 >>
rect 2700 -3420 2820 -3400
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3780 3060 -3420
rect 2940 -3800 3060 -3780
rect -1200 -4440 -1120 -4430
rect -1200 -4500 -1190 -4440
rect -1130 -4500 -1120 -4440
rect -1200 -4510 -1120 -4500
rect -4369 -7084 -4329 -6884
rect -4301 -7084 -4261 -6884
<< via1 >>
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
rect -1190 -4500 -1130 -4440
<< metal2 >>
rect -5500 580 -5240 600
rect -5500 120 -5480 580
rect -5260 120 -5240 580
rect -5500 -2820 -5240 120
rect -2600 0 2000 100
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 2400 -3000 2540 -2980
rect 2400 -3080 2420 -3000
rect 1860 -3140 2060 -3100
rect 2120 -3140 2420 -3080
rect 2520 -3140 2540 -3000
rect 2120 -3160 2540 -3140
rect 2700 -3420 2820 -3400
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3780 3060 -3420
rect 2940 -3800 3060 -3780
rect -1400 -4440 -1120 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1190 -4440
rect -1130 -4500 -1120 -4440
rect -1400 -4510 -1120 -4500
rect -2840 -6200 -2340 -5800
rect -2840 -6500 -1600 -6200
rect -2840 -6700 -2340 -6500
rect -4200 -6952 -4120 -6843
rect -4200 -7008 -4014 -6952
rect -3320 -7000 -1600 -6700
rect 1600 -7000 2000 -5800
rect -4200 -7084 -4120 -7008
rect -3000 -7100 -1200 -7000
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via2 >>
rect -5480 120 -5260 580
rect -2500 -500 1900 0
rect 2420 -3140 2520 -3000
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
rect -1390 -4500 -1230 -4440
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< metal3 >>
rect -5500 580 -5240 600
rect -5500 120 -5480 580
rect -5260 120 -5240 580
rect -5500 100 -5240 120
rect -2600 0 2000 100
rect -7600 -7100 -4800 -200
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 2400 -3000 2540 -2980
rect 2400 -3140 2420 -3000
rect 2520 -3140 2540 -3000
rect 2700 -3100 4300 700
rect 2400 -3160 2540 -3140
rect 2600 -3231 2820 -3220
rect 1904 -3305 2820 -3231
rect 2600 -3320 2820 -3305
rect 2700 -3420 2820 -3320
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3620 3060 -3420
rect 3380 -3520 4300 -3100
rect 3380 -3620 3400 -3520
rect 3040 -3740 3400 -3620
rect 3040 -3780 3060 -3740
rect 2940 -3800 3060 -3780
rect 3380 -3840 3400 -3740
rect 4280 -3840 4300 -3520
rect 3380 -3860 4300 -3840
rect -660 -4200 -620 -4180
rect 120 -4200 160 -4180
rect -1400 -4440 -1220 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1220 -4440
rect -3600 -5700 -2800 -5600
rect -1400 -5700 -1220 -4500
rect -3600 -5800 -1220 -5700
rect -3000 -6000 -1220 -5800
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 -1200 -7000
rect -4900 -7600 -4600 -7300
rect -4900 -7700 -4800 -7600
rect -7600 -7800 -4800 -7700
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via3 >>
rect -5480 120 -5260 580
rect -2500 -500 1900 0
rect 2420 -3140 2520 -3000
rect 3400 -3840 4280 -3520
rect -7500 -7700 -4900 -7100
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< mimcap >>
rect 2800 560 4200 600
rect -7500 -340 -4900 -300
rect -7500 -6460 -7460 -340
rect -4940 -6460 -4900 -340
rect 2800 -2960 2840 560
rect 4160 -2960 4200 560
rect 2800 -3000 4200 -2960
rect -7500 -6500 -4900 -6460
<< mimcapcontact >>
rect -7460 -6460 -4940 -340
rect 2840 -2960 4160 560
<< metal4 >>
rect -7400 580 2000 600
rect -7400 120 -5480 580
rect -5260 120 2000 580
rect -7400 100 2000 120
rect -7400 -200 -5000 100
rect -2600 0 2000 100
rect -7600 -340 -4800 -200
rect -7600 -6460 -7460 -340
rect -4940 -6460 -4800 -340
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 2700 560 4300 700
rect 2700 -2960 2840 560
rect 4160 -2960 4300 560
rect 2700 -2980 4300 -2960
rect 2400 -3000 4300 -2980
rect 2400 -3140 2420 -3000
rect 2520 -3100 4300 -3000
rect 2520 -3140 2540 -3100
rect 2400 -3160 2540 -3140
rect 3380 -3520 4300 -3500
rect 3380 -3840 3400 -3520
rect 4280 -3840 4300 -3520
rect 3380 -3860 4300 -3840
rect -7600 -6600 -4800 -6460
rect -7600 -7100 -4800 -7000
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 2000 -7000
rect -3000 -7300 -2900 -7100
rect -4900 -7700 -2900 -7300
rect -1300 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect -7600 -7800 2000 -7700
<< via4 >>
rect 3420 -3820 4260 -3540
rect -7500 -7700 -4900 -7100
<< mimcap2 >>
rect 2800 560 4200 600
rect -7500 -340 -4900 -300
rect -7500 -6460 -7460 -340
rect -4940 -6460 -4900 -340
rect 2800 -2960 2840 560
rect 4160 -2960 4200 560
rect 2800 -3000 4200 -2960
rect -7500 -6500 -4900 -6460
<< mimcap2contact >>
rect -7460 -6460 -4940 -340
rect 2840 -2960 4160 560
<< metal5 >>
rect 2700 560 4300 700
rect -7600 -340 -4800 -200
rect -7600 -6460 -7460 -340
rect -4940 -6460 -4800 -340
rect 2700 -2960 2840 560
rect 4160 -2960 4300 560
rect 2700 -3100 4300 -2960
rect 3380 -3540 4300 -3100
rect 3380 -3820 3420 -3540
rect 4260 -3820 4300 -3540
rect 3380 -3860 4300 -3820
rect -7600 -7100 -4800 -6460
rect -7600 -7700 -7500 -7100
rect -4900 -7700 -4800 -7100
rect -7600 -7800 -4800 -7700
use cmota_1_flat_1  cmota_1_flat_1_0
timestamp 1671334909
transform 1 0 -2836 0 1 -3200
box -164 -3800 5363 2800
use gated_iref_fix  gated_iref_fix_0
timestamp 1672205966
transform 0 1 -4300 1 0 -7948
box 940 -2420 7820 1220
use sky130_fd_pr__res_high_po_0p69_N63KD6  sky130_fd_pr__res_high_po_0p69_N63KD6_0
timestamp 1671858438
transform 1 0 2879 0 -1 -3778
box -352 -564 352 564
<< labels >>
rlabel metal4 -3840 -7800 -3660 -7300 1 VLO
rlabel metal4 -4220 320 -3840 600 1 VHI
rlabel metal3 -660 -4200 -620 -4180 1 VIN
rlabel metal3 120 -4200 160 -4180 1 VIP
rlabel metal2 1860 -3140 2060 -3100 1 VOP
rlabel metal1 -4369 -7084 -4329 -7044 1 S
rlabel metal1 -4301 -7084 -4261 -7044 1 SBAR
rlabel metal2 -4200 -7084 -4120 -7004 1 VREF
<< end >>
