magic
tech sky130A
magscale 1 2
timestamp 1672206264
<< nwell >>
rect 2001 1514 2113 1614
rect 2538 1519 2909 1531
rect 2538 1514 3180 1519
rect 2001 1488 3180 1514
rect 2001 1430 2113 1488
rect 2882 1212 3180 1488
<< locali >>
rect 2286 2472 2392 2568
rect 2295 1856 2401 1952
rect 10180 1930 10280 1950
rect 10120 1850 10200 1930
rect 10260 1850 10280 1930
rect 10180 1830 10280 1850
rect 10180 1240 10280 1260
rect 3421 1140 3529 1236
rect 10180 1220 10200 1240
rect 10160 1160 10200 1220
rect 10260 1160 10280 1240
rect 10180 1140 10280 1160
rect 39160 1008 39260 1210
rect 38946 470 39260 1008
rect 38946 380 39170 470
rect 39250 380 39260 470
rect 45074 487 45176 494
rect 45074 453 45130 487
rect 45164 453 45176 487
rect 45074 446 45176 453
rect 38946 -126 39260 380
rect 45089 300 45137 365
rect 45100 173 45137 300
rect 39160 -320 39260 -126
rect 45074 -525 45176 -518
rect 45074 -559 45130 -525
rect 45164 -559 45176 -525
rect 45074 -566 45176 -559
rect 45089 -712 45137 -647
rect 10514 -793 10616 -786
rect 10514 -827 10570 -793
rect 10604 -827 10616 -793
rect 10514 -834 10616 -827
rect 45100 -839 45137 -712
rect 10529 -980 10577 -915
rect 10540 -1107 10577 -980
<< viali >>
rect 10200 1850 10260 1930
rect 10200 1160 10260 1240
rect 39170 380 39250 470
rect 45130 453 45164 487
rect 45130 -559 45164 -525
rect 10570 -827 10604 -793
<< metal1 >>
rect 11463 5180 11503 6156
rect 11050 5140 11503 5180
rect 11050 4920 11090 5140
rect 11531 5100 11571 6156
rect 47771 5310 47811 6160
rect 11210 5060 11571 5100
rect 45790 5270 47811 5310
rect 11210 4920 11250 5060
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 10180 1930 10280 1950
rect 10180 1850 10200 1930
rect 10260 1850 10280 1930
rect 10180 1830 10280 1850
rect 10180 1240 10280 1260
rect 1880 1220 2020 1240
rect 1880 1120 1900 1220
rect 2000 1120 2020 1220
rect 1880 1100 2020 1120
rect 2240 1220 2380 1240
rect 2240 1120 2260 1220
rect 2360 1120 2380 1220
rect 2240 1100 2380 1120
rect 2620 1220 2760 1240
rect 2620 1120 2640 1220
rect 2740 1120 2760 1220
rect 10180 1160 10200 1240
rect 10260 1160 10280 1240
rect 10180 1140 10280 1160
rect 2620 1100 2760 1120
rect 39370 980 39390 1040
rect 39770 980 39790 1040
rect 39900 980 39920 1040
rect 40300 980 40320 1040
rect 1680 920 3287 954
rect 1680 858 1740 920
rect 1720 800 1740 858
rect 1820 860 2080 920
rect 1820 858 2040 860
rect 1820 800 1840 858
rect 1720 780 1840 800
rect 2060 800 2080 860
rect 2160 858 3287 920
rect 2160 800 2180 858
rect 39370 820 39390 880
rect 39770 820 39790 880
rect 39900 820 39920 880
rect 40300 820 40320 880
rect 44580 860 44840 880
rect 2060 780 2180 800
rect 39370 650 39390 710
rect 39770 650 39790 710
rect 39900 650 39920 710
rect 40300 650 40320 710
rect 8100 520 8120 620
rect 8260 520 8280 620
rect 39370 490 39390 550
rect 39770 490 39790 550
rect 44580 540 44600 860
rect 44720 540 44740 860
rect 39150 480 39270 490
rect 39900 480 39920 540
rect 40300 480 40320 540
rect 44580 520 44740 540
rect 38930 470 39270 480
rect 38930 380 39170 470
rect 39250 380 39270 470
rect 38930 370 39270 380
rect 39150 360 39270 370
rect 39370 320 39390 380
rect 39770 320 39790 380
rect 39900 310 39920 370
rect 40300 310 40320 370
rect 8020 280 8360 300
rect 8020 200 8040 280
rect 8340 200 8360 280
rect 8020 180 8360 200
rect 39370 160 39390 220
rect 39770 160 39790 220
rect 39900 210 40320 211
rect 39900 150 39920 210
rect 40300 150 40320 210
rect 39900 50 40320 51
rect 39370 -10 39390 50
rect 39770 -10 39790 50
rect 39900 -10 39920 50
rect 40300 -10 40320 50
rect 39900 -120 40320 -119
rect 39370 -180 39390 -120
rect 39770 -180 39790 -120
rect 39900 -180 39920 -120
rect 40300 -180 40320 -120
rect 10020 -420 10280 -400
rect 10780 -420 10980 -400
rect 10020 -740 10040 -420
rect 10160 -740 10280 -420
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10020 -760 10280 -740
rect 10780 -740 10800 -420
rect 10960 -740 10980 -420
rect 10780 -760 10980 -740
rect 45310 860 45540 880
rect 45520 540 45540 860
rect 45310 520 45540 540
rect 45106 494 45112 505
rect 45074 453 45112 494
rect 45164 494 45170 505
rect 45164 453 45176 494
rect 45074 446 45176 453
rect 45310 230 45440 520
rect 45040 150 45200 160
rect 45040 40 45050 150
rect 45190 40 45200 150
rect 45040 30 45200 40
rect 45060 -210 45190 -200
rect 45060 -340 45070 -210
rect 45180 -340 45190 -210
rect 45060 -350 45190 -340
rect 44740 -612 44840 -430
rect 45106 -518 45112 -507
rect 45074 -559 45112 -518
rect 45164 -518 45170 -507
rect 45320 -512 45440 230
rect 45790 200 45830 5270
rect 47839 5220 47879 6160
rect 45880 5180 47879 5220
rect 45880 650 45920 5180
rect 45880 610 46010 650
rect 45970 500 46010 610
rect 45940 490 46040 500
rect 45940 410 45950 490
rect 46030 410 46040 490
rect 45940 400 46040 410
rect 45760 190 45860 200
rect 45760 110 45770 190
rect 45850 110 45860 190
rect 45760 100 45860 110
rect 45164 -559 45176 -518
rect 45074 -566 45176 -559
rect 10546 -786 10552 -775
rect 10514 -827 10552 -786
rect 10604 -786 10610 -775
rect 10604 -827 10616 -786
rect 10514 -834 10616 -827
rect 11200 -790 11300 -780
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 10480 -1130 10640 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 10480 -1250 10640 -1240
rect 11230 -1210 11270 -880
rect 11380 -1090 11480 -1080
rect 11380 -1170 11390 -1090
rect 11470 -1110 11480 -1090
rect 11470 -1150 11571 -1110
rect 11470 -1170 11480 -1150
rect 11380 -1180 11480 -1170
rect 11230 -1250 11503 -1210
rect 10500 -1490 10630 -1480
rect 10500 -1620 10510 -1490
rect 10620 -1620 10630 -1490
rect 10500 -1630 10630 -1620
rect 11463 -2760 11503 -1250
rect 11531 -2760 11571 -1150
rect 45310 -782 45440 -512
rect 45760 -522 45860 -512
rect 45760 -602 45770 -522
rect 45850 -540 45860 -522
rect 45850 -580 46110 -540
rect 45850 -602 45860 -580
rect 45760 -612 45860 -602
rect 45790 -620 45830 -612
rect 45040 -862 45200 -852
rect 45040 -972 45050 -862
rect 45190 -972 45200 -862
rect 45040 -982 45200 -972
rect 44740 -1160 44840 -1112
rect 45320 -1460 45440 -782
rect 45940 -822 46040 -812
rect 45940 -902 45950 -822
rect 46030 -902 46040 -822
rect 45940 -910 46040 -902
rect 45940 -912 46000 -910
rect 45960 -1890 46000 -912
rect 46070 -1810 46110 -580
rect 46070 -1850 47879 -1810
rect 45960 -1930 47811 -1890
rect 47771 -2760 47811 -1930
rect 47839 -2756 47879 -1850
<< via1 >>
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 10200 1850 10260 1930
rect 1900 1120 2000 1220
rect 2260 1120 2360 1220
rect 2640 1120 2740 1220
rect 10200 1160 10260 1240
rect 39390 980 39770 1040
rect 39920 980 40300 1040
rect 1740 800 1820 920
rect 2080 800 2160 920
rect 39390 820 39770 880
rect 39920 820 40300 880
rect 39390 650 39770 710
rect 39920 650 40300 710
rect 8120 520 8260 620
rect 39390 490 39770 550
rect 44600 540 44720 860
rect 39920 480 40300 540
rect 39390 320 39770 380
rect 39920 310 40300 370
rect 8040 200 8340 280
rect 39390 160 39770 220
rect 39920 150 40300 210
rect 39390 -10 39770 50
rect 39920 -10 40300 50
rect 39390 -180 39770 -120
rect 39920 -180 40300 -120
rect 10040 -740 10160 -420
rect 10500 -700 10620 -440
rect 10800 -740 10960 -420
rect 44740 -430 44840 860
rect 45310 540 45520 860
rect 45112 487 45164 505
rect 45112 453 45130 487
rect 45130 453 45164 487
rect 45050 40 45190 150
rect 45070 -340 45180 -210
rect 45112 -525 45164 -507
rect 45950 410 46030 490
rect 45770 110 45850 190
rect 45112 -559 45130 -525
rect 45130 -559 45164 -525
rect 10552 -793 10604 -775
rect 10552 -827 10570 -793
rect 10570 -827 10604 -793
rect 11210 -870 11290 -790
rect 10490 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 10510 -1620 10620 -1490
rect 44740 -1112 44840 -612
rect 45770 -602 45850 -522
rect 45050 -972 45190 -862
rect 45950 -902 46030 -822
<< metal2 >>
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11322 4770 11402 6196
rect 47950 6060 48200 6290
rect 48048 5001 48131 6060
rect 46218 4918 48131 5001
rect 11320 4760 11420 4770
rect 11320 4680 11330 4760
rect 11410 4680 11420 4760
rect 11320 4670 11420 4680
rect 9240 4260 14440 4280
rect 9240 2960 9260 4260
rect 14420 3960 14440 4260
rect 9460 3940 14440 3960
rect 9460 3880 10460 3940
rect 9460 2960 9480 3880
rect 9240 2940 9480 2960
rect 9240 2880 9440 2940
rect 1920 2540 2040 2560
rect 1920 2460 1940 2540
rect 2020 2460 2367 2540
rect 1920 2440 2040 2460
rect 1920 1960 2040 1980
rect 1920 1880 1940 1960
rect 2020 1880 2347 1960
rect 10180 1930 10280 1950
rect 1920 1860 2040 1880
rect 10180 1850 10200 1930
rect 10260 1850 10280 1930
rect 10180 1830 10280 1850
rect 5208 1750 5238 1786
rect 5046 1650 5084 1700
rect 8928 1252 8966 1302
rect 10180 1240 10280 1260
rect 1880 1220 2020 1240
rect 1880 1120 1900 1220
rect 2000 1120 2020 1220
rect 1880 1100 2020 1120
rect 2240 1220 2380 1240
rect 2240 1120 2260 1220
rect 2360 1120 2380 1220
rect 2240 1040 2380 1120
rect 2240 960 2260 1040
rect 2360 960 2380 1040
rect 2240 940 2380 960
rect 2620 1220 2760 1240
rect 2620 1120 2640 1220
rect 2740 1120 2760 1220
rect 1720 920 1840 940
rect 1720 800 1740 920
rect 1820 800 1840 920
rect 1720 780 1840 800
rect 2060 920 2180 940
rect 2060 800 2080 920
rect 2160 800 2180 920
rect 2060 780 2180 800
rect 2620 860 2760 1120
rect 2620 780 2640 860
rect 2740 780 2760 860
rect 2620 760 2760 780
rect 8200 620 8240 1220
rect 10180 1160 10200 1240
rect 10260 1160 10280 1240
rect 10180 1140 10280 1160
rect 39900 1040 40320 1050
rect 39370 1030 39390 1040
rect 39140 990 39390 1030
rect 11070 920 11390 940
rect 8100 600 8120 620
rect 7730 540 8120 600
rect 1560 -850 1660 -840
rect 7730 -850 7790 540
rect 8100 520 8120 540
rect 8260 520 8280 620
rect 8020 280 8360 300
rect 8020 200 8040 280
rect 8340 200 8360 280
rect 8020 180 8360 200
rect 9880 120 10080 880
rect 11070 840 11090 920
rect 11190 840 11390 920
rect 11070 820 11390 840
rect 39140 809 39180 990
rect 39370 980 39390 990
rect 39770 980 39790 1040
rect 39900 980 39920 1040
rect 40300 980 40320 1040
rect 39900 970 40320 980
rect 39900 880 40320 890
rect 39370 870 39390 880
rect 39018 769 39180 809
rect 39210 830 39390 870
rect 39210 689 39250 830
rect 39370 820 39390 830
rect 39770 820 39790 880
rect 39900 820 39920 880
rect 40300 820 40320 880
rect 39900 810 40320 820
rect 44580 860 44840 880
rect 39900 710 40320 720
rect 39370 700 39390 710
rect 39018 649 39250 689
rect 39280 660 39390 700
rect 39280 619 39320 660
rect 39370 650 39390 660
rect 39770 650 39790 710
rect 39900 650 39920 710
rect 40300 650 40320 710
rect 39900 640 40320 650
rect 39018 579 39320 619
rect 39370 549 39390 550
rect 39018 509 39390 549
rect 39370 490 39390 509
rect 39770 490 39790 550
rect 39900 540 40320 550
rect 39900 480 39920 540
rect 40300 480 40320 540
rect 44580 540 44600 860
rect 44720 540 44740 860
rect 44580 520 44740 540
rect 39018 439 39330 479
rect 39900 470 40320 480
rect 39018 369 39260 409
rect 39018 299 39190 339
rect 39018 229 39120 269
rect 9880 100 14400 120
rect 9880 -180 9900 100
rect 14380 -180 14400 100
rect 39080 -130 39120 229
rect 39150 40 39190 299
rect 39220 210 39260 369
rect 39290 370 39330 439
rect 39370 370 39390 380
rect 39290 330 39390 370
rect 39370 320 39390 330
rect 39770 320 39790 380
rect 39900 370 40320 380
rect 39900 310 39920 370
rect 40300 310 40320 370
rect 39900 300 40320 310
rect 39370 210 39390 220
rect 39220 170 39390 210
rect 39370 160 39390 170
rect 39770 160 39790 220
rect 39900 210 40320 220
rect 39900 150 39920 210
rect 40300 150 40320 210
rect 39900 140 40320 150
rect 44510 150 44650 160
rect 39900 50 40320 60
rect 39370 40 39390 50
rect 39150 0 39390 40
rect 39370 -10 39390 0
rect 39770 -10 39790 50
rect 39900 -10 39920 50
rect 40300 -10 40320 50
rect 44510 40 44520 150
rect 44640 40 44650 150
rect 44510 30 44650 40
rect 39900 -20 40320 -10
rect 39900 -120 40320 -110
rect 39370 -130 39390 -120
rect 39080 -170 39390 -130
rect 39370 -180 39390 -170
rect 39770 -180 39790 -120
rect 39900 -180 39920 -120
rect 40300 -180 40320 -120
rect 9880 -200 14400 -180
rect 39900 -190 40320 -180
rect 10020 -420 10280 -400
rect 10780 -420 10980 -400
rect 10020 -740 10040 -420
rect 10160 -740 10280 -420
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10020 -760 10280 -740
rect 10780 -740 10800 -420
rect 10960 -740 10980 -420
rect 10780 -760 10980 -740
rect 45310 860 45540 880
rect 45520 540 45540 860
rect 45310 520 45540 540
rect 45106 494 45112 505
rect 45074 453 45112 494
rect 45164 494 45170 505
rect 45164 480 45176 494
rect 45940 490 46040 500
rect 45164 453 45520 480
rect 45074 450 45520 453
rect 45074 446 45440 450
rect 45110 440 45440 446
rect 45430 390 45440 440
rect 45510 390 45520 450
rect 45940 410 45950 490
rect 46030 410 46040 490
rect 45940 400 46040 410
rect 45430 380 45520 390
rect 45760 190 45860 200
rect 45040 150 45200 160
rect 45040 40 45050 150
rect 45190 40 45200 150
rect 45760 110 45770 190
rect 45850 110 45860 190
rect 45760 100 45860 110
rect 45040 30 45200 40
rect 46218 -30 46301 4918
rect 46210 -200 46310 -30
rect 45060 -210 45190 -200
rect 45060 -340 45070 -210
rect 45180 -340 45190 -210
rect 45870 -210 46310 -200
rect 45870 -290 45880 -210
rect 45960 -282 46310 -210
rect 45960 -290 45970 -282
rect 45870 -300 45970 -290
rect 45060 -350 45190 -340
rect 44740 -612 44840 -430
rect 45106 -518 45112 -507
rect 45074 -559 45112 -518
rect 45164 -518 45170 -507
rect 45164 -532 45176 -518
rect 45760 -522 45860 -512
rect 45164 -559 45520 -532
rect 45074 -562 45520 -559
rect 45074 -566 45440 -562
rect 45110 -572 45440 -566
rect 10546 -786 10552 -775
rect 10514 -827 10552 -786
rect 10604 -786 10610 -775
rect 10604 -800 10616 -786
rect 11200 -790 11300 -780
rect 10604 -827 10960 -800
rect 10514 -830 10960 -827
rect 10514 -834 10880 -830
rect 10550 -840 10880 -834
rect 1560 -860 7790 -850
rect 1560 -940 1580 -860
rect 1640 -910 7790 -860
rect 10870 -890 10880 -840
rect 10950 -890 10960 -830
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 44510 -862 44650 -852
rect 10870 -900 10960 -890
rect 1640 -940 1660 -910
rect 1560 -960 1660 -940
rect 44510 -972 44520 -862
rect 44640 -972 44650 -862
rect 44510 -982 44650 -972
rect 11380 -1090 11480 -1080
rect 10480 -1130 10640 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 11380 -1170 11390 -1090
rect 11470 -1170 11480 -1090
rect 45430 -622 45440 -572
rect 45510 -622 45520 -562
rect 45760 -602 45770 -522
rect 45850 -602 45860 -522
rect 45760 -612 45860 -602
rect 45430 -632 45520 -622
rect 45940 -822 46040 -812
rect 45040 -862 45200 -852
rect 45040 -972 45050 -862
rect 45190 -972 45200 -862
rect 45940 -902 45950 -822
rect 46030 -902 46040 -822
rect 45940 -910 46040 -902
rect 45940 -912 46000 -910
rect 45040 -982 45200 -972
rect 44740 -1160 44840 -1112
rect 11380 -1180 11480 -1170
rect 10480 -1250 10640 -1240
rect 10500 -1490 10630 -1480
rect 10500 -1620 10510 -1490
rect 10620 -1620 10630 -1490
rect 11310 -1490 11410 -1480
rect 11310 -1570 11320 -1490
rect 11400 -1570 11410 -1490
rect 11310 -1580 11410 -1570
rect 10500 -1630 10630 -1620
rect 1720 -2600 5860 -2580
rect 1720 -2780 1760 -2600
rect 1820 -2780 2080 -2600
rect 2140 -2780 5860 -2600
rect 1720 -2800 5860 -2780
rect 11321 -2800 11404 -1580
rect 46219 -1689 46302 -282
rect 46219 -1772 48141 -1689
rect 48058 -2690 48141 -1772
rect 11321 -2831 11440 -2800
rect 11402 -2859 11440 -2831
rect 47940 -2870 48200 -2690
rect 48978 -10423 49064 -6157
<< via2 >>
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 11330 4680 11410 4760
rect 9260 3960 14420 4260
rect 9260 2960 9460 3960
rect 1940 2460 2020 2540
rect 1940 1880 2020 1960
rect 10200 1850 10260 1930
rect 1900 1120 2000 1220
rect 2260 960 2360 1040
rect 1740 800 1820 920
rect 2080 800 2160 920
rect 2640 780 2740 860
rect 10200 1160 10260 1240
rect 8040 200 8340 280
rect 11090 840 11190 920
rect 39920 980 40300 1040
rect 39920 820 40300 880
rect 39920 650 40300 710
rect 39920 480 40300 540
rect 44600 540 44720 860
rect 9900 -180 14380 100
rect 39920 310 40300 370
rect 39920 150 40300 210
rect 39920 -10 40300 50
rect 44520 40 44640 150
rect 39920 -180 40300 -120
rect 10040 -740 10160 -420
rect 10500 -700 10620 -440
rect 10880 -740 10960 -420
rect 45330 540 45520 860
rect 45440 390 45510 450
rect 45950 410 46030 490
rect 45050 40 45190 150
rect 45770 110 45850 190
rect 45070 -340 45180 -210
rect 45880 -290 45960 -210
rect 1580 -940 1640 -860
rect 10880 -890 10950 -830
rect 11210 -870 11290 -790
rect 44520 -972 44640 -862
rect 10490 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 45440 -622 45510 -562
rect 45770 -602 45850 -522
rect 45050 -972 45190 -862
rect 45950 -902 46030 -822
rect 10510 -1620 10620 -1490
rect 11320 -1570 11400 -1490
rect 1760 -2780 1820 -2600
rect 2080 -2780 2140 -2600
<< metal3 >>
rect 54430 10250 54630 10260
rect 54430 10120 54440 10250
rect 54510 10120 54630 10250
rect 54430 10110 54630 10120
rect 50680 9040 50920 9050
rect 7300 7240 7500 9020
rect -1020 7180 -520 7240
rect -40 7180 7500 7240
rect -1020 7100 7500 7180
rect -1020 7040 -520 7100
rect -40 7040 7500 7100
rect -1020 -7320 -820 7040
rect 8480 5180 8680 9020
rect 50680 8940 50690 9040
rect 50910 8940 50920 9040
rect 50680 8930 50920 8940
rect 8480 4980 14900 5180
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11320 4760 11420 4770
rect 11320 4680 11330 4760
rect 11410 4680 11420 4760
rect 11320 4670 11420 4680
rect -380 4440 -180 4460
rect -380 4280 -360 4440
rect -200 4280 -180 4440
rect -380 4260 -180 4280
rect 8600 4260 14440 4280
rect -340 2560 -220 4260
rect 8600 3960 8620 4260
rect 14420 3960 14440 4260
rect 8600 3940 9260 3960
rect 9240 2960 9260 3940
rect 9460 3940 14440 3960
rect 9460 2960 9480 3940
rect 9240 2920 9480 2960
rect 14700 2660 14900 4980
rect 14600 2620 15000 2660
rect -340 2540 2040 2560
rect -340 2460 1940 2540
rect 2020 2460 2040 2540
rect -340 2440 2040 2460
rect 14600 2300 14640 2620
rect 14960 2300 15000 2620
rect 14600 2260 15000 2300
rect 13520 1980 14460 2040
rect -340 1960 2040 1980
rect -340 1880 1940 1960
rect 2020 1880 2040 1960
rect 10280 1950 14460 1980
rect 40000 1950 40600 2000
rect -340 1860 2040 1880
rect 10180 1930 13620 1950
rect -340 0 -220 1860
rect 10180 1850 10200 1930
rect 10260 1880 13620 1930
rect 10260 1850 10280 1880
rect 10180 1830 10280 1850
rect 10970 1410 11730 1510
rect 10180 1240 10280 1260
rect 1880 1220 3121 1240
rect 1880 1120 1900 1220
rect 2000 1120 3121 1220
rect 10180 1160 10200 1240
rect 10260 1230 10280 1240
rect 10970 1230 11070 1410
rect 10260 1160 11070 1230
rect 10180 1140 11070 1160
rect 10280 1130 11070 1140
rect 11630 1160 11730 1410
rect 13748 1160 13808 1540
rect 14400 1410 14460 1950
rect 14260 1350 14460 1410
rect 39150 1900 40600 1950
rect 39150 1700 40100 1900
rect 40500 1700 40600 1900
rect 39150 1650 40600 1700
rect 1880 1100 2020 1120
rect 1720 920 1840 940
rect 1720 800 1740 920
rect 1820 800 1840 920
rect 1720 780 1840 800
rect -380 -20 -180 0
rect -380 -180 -360 -20
rect -200 -180 -180 -20
rect -380 -200 -180 -180
rect 1560 -860 1660 -840
rect 1560 -940 1580 -860
rect 1640 -940 1660 -860
rect 1560 -6680 1660 -940
rect 1740 -2600 1840 780
rect 1740 -2780 1760 -2600
rect 1820 -2780 1840 -2600
rect 1740 -6680 1840 -2780
rect 1900 -6680 2000 1100
rect 11630 1060 13830 1160
rect 2240 1040 2780 1060
rect 2240 960 2260 1040
rect 2360 960 2780 1040
rect 2240 940 2780 960
rect 2060 920 2180 940
rect 2060 800 2080 920
rect 2160 800 2180 920
rect 2060 780 2180 800
rect 2060 -2600 2160 780
rect 2060 -2780 2080 -2600
rect 2140 -2780 2160 -2600
rect 2060 -6680 2160 -2780
rect 2240 -6680 2360 940
rect 11070 920 11210 940
rect 2620 860 2900 880
rect 2620 840 2640 860
rect 1580 -7320 1640 -6680
rect 1760 -7320 1820 -6680
rect 1920 -7320 1980 -6680
rect 2080 -7320 2140 -6680
rect 2300 -7320 2360 -6680
rect -1020 -7520 1480 -7320
rect 1360 -9060 1480 -7520
rect 1560 -9060 1660 -7320
rect 1740 -9060 1840 -7320
rect 1900 -9060 2000 -7320
rect 2060 -9060 2160 -7320
rect 2240 -9060 2360 -7320
rect 2420 780 2640 840
rect 2740 780 2900 860
rect 11070 840 11090 920
rect 11190 840 11210 920
rect 11070 820 11210 840
rect 2420 760 2900 780
rect 2420 -6680 2540 760
rect 39150 589 39450 1650
rect 40000 1600 40600 1650
rect 39900 1040 40320 1050
rect 39900 980 39920 1040
rect 40300 980 40530 1040
rect 39900 970 40320 980
rect 39900 880 40320 890
rect 39900 820 39920 880
rect 40300 820 40530 880
rect 44580 860 44740 880
rect 39900 810 40320 820
rect 39900 710 40320 720
rect 39900 650 39920 710
rect 40300 650 40530 710
rect 39900 640 40320 650
rect 8020 280 8360 300
rect 8020 200 8040 280
rect 8340 200 8360 280
rect 8020 180 8360 200
rect 14380 120 14700 580
rect 38550 289 39450 589
rect 39900 540 40320 550
rect 44580 540 44600 860
rect 44720 540 44740 860
rect 39900 480 39920 540
rect 40300 480 40530 540
rect 44580 520 44740 540
rect 45310 860 45540 880
rect 45310 540 45330 860
rect 45520 540 45540 860
rect 45310 520 45540 540
rect 45940 490 46040 500
rect 39900 470 40320 480
rect 45430 450 45620 460
rect 45430 380 45440 450
rect 45610 380 45620 450
rect 45940 410 45950 490
rect 46030 410 46040 490
rect 45940 400 46040 410
rect 39900 370 40320 380
rect 45430 370 45620 380
rect 39900 310 39920 370
rect 40300 310 40530 370
rect 39900 300 40320 310
rect 9880 100 14700 120
rect 9880 -180 9900 100
rect 14380 -180 14700 100
rect 9880 -200 14700 -180
rect 10020 -420 10180 -400
rect 10860 -420 10980 -200
rect 10020 -740 10040 -420
rect 10160 -740 10180 -420
rect 10480 -440 10640 -420
rect 10480 -540 10500 -440
rect 10020 -760 10180 -740
rect 10240 -650 10500 -540
rect 10240 -980 10300 -650
rect 10480 -700 10500 -650
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10860 -740 10880 -420
rect 10960 -740 10980 -420
rect 10860 -760 10980 -740
rect 11200 -790 11300 -780
rect 10870 -830 11060 -820
rect 10870 -900 10880 -830
rect 11050 -900 11060 -830
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 39150 -850 39450 289
rect 39900 210 40320 220
rect 39900 150 39920 210
rect 40300 150 40530 210
rect 45760 190 45860 200
rect 44510 150 45200 160
rect 39900 140 40320 150
rect 39900 50 40320 60
rect 39900 -10 39920 50
rect 40300 -10 40530 50
rect 44510 40 44520 150
rect 44640 40 45050 150
rect 45190 40 45200 150
rect 45760 110 45770 190
rect 45850 110 45860 190
rect 45760 100 45860 110
rect 44510 30 45200 40
rect 39900 -20 40320 -10
rect 39900 -120 40320 -110
rect 39900 -180 39920 -120
rect 40300 -180 40530 -120
rect 39900 -190 40320 -180
rect 45060 -210 45190 -200
rect 45060 -340 45070 -210
rect 45180 -340 45190 -210
rect 45870 -210 45970 -200
rect 45870 -290 45880 -210
rect 45960 -290 45970 -210
rect 45870 -300 45970 -290
rect 45060 -350 45190 -340
rect 45760 -522 45860 -512
rect 45430 -562 45620 -552
rect 45430 -632 45440 -562
rect 45610 -632 45620 -562
rect 45760 -602 45770 -522
rect 45850 -602 45860 -522
rect 45760 -612 45860 -602
rect 45430 -642 45620 -632
rect 40000 -850 40600 -800
rect 10870 -910 11060 -900
rect 39150 -900 40600 -850
rect 45940 -822 46040 -812
rect 2780 -1100 10300 -980
rect 14600 -1040 15000 -1000
rect 11380 -1090 11480 -1080
rect 2600 -4120 2720 -4100
rect 2600 -4280 2620 -4120
rect 2700 -4280 2720 -4120
rect 2600 -6680 2720 -4280
rect 2780 -6680 2900 -1100
rect 10480 -1130 10640 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 11380 -1170 11390 -1090
rect 11470 -1170 11480 -1090
rect 11380 -1180 11480 -1170
rect 10480 -1250 10640 -1240
rect 3000 -1251 10640 -1250
rect 2960 -1370 10640 -1251
rect 14600 -1360 14640 -1040
rect 14960 -1360 15000 -1040
rect 39150 -1100 40100 -900
rect 40500 -1100 40600 -900
rect 44510 -862 45200 -852
rect 44510 -972 44520 -862
rect 44640 -972 45050 -862
rect 45190 -972 45200 -862
rect 45940 -902 45950 -822
rect 46030 -902 46040 -822
rect 45940 -910 46040 -902
rect 45940 -912 46000 -910
rect 44510 -982 45200 -972
rect 39150 -1150 40600 -1100
rect 40000 -1200 40600 -1150
rect 2960 -6680 3080 -1370
rect 14600 -1400 15000 -1360
rect 3140 -1490 10630 -1480
rect 3140 -1600 10510 -1490
rect 3140 -6680 3260 -1600
rect 10500 -1620 10510 -1600
rect 10620 -1620 10630 -1490
rect 11310 -1490 11410 -1480
rect 11310 -1570 11320 -1490
rect 11400 -1570 11410 -1490
rect 11310 -1580 11410 -1570
rect 10500 -1630 10630 -1620
rect 14700 -1700 14900 -1400
rect 7700 -1900 14900 -1700
rect 7700 -5600 7900 -1900
rect 8100 -5420 8300 -5400
rect 8100 -5580 8120 -5420
rect 8280 -5580 8300 -5420
rect 8100 -5600 8300 -5580
rect 50680 -5540 50920 -5530
rect 50680 -5640 50690 -5540
rect 50910 -5640 50920 -5540
rect 50680 -5650 50920 -5640
rect 2420 -7320 2480 -6680
rect 2630 -7320 2690 -6680
rect 2810 -7320 2870 -6680
rect 2990 -7320 3050 -6680
rect 3170 -7320 3230 -6680
rect 54430 -6720 54630 -6710
rect 54430 -6850 54440 -6720
rect 54510 -6850 54630 -6720
rect 54430 -6860 54630 -6850
rect 2420 -9060 2540 -7320
rect 2600 -9060 2720 -7320
rect 2780 -9060 2900 -7320
rect 2960 -9060 3080 -7320
rect 3140 -9060 3260 -7320
<< via3 >>
rect 54440 10120 54510 10250
rect 50690 8940 50910 9040
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 11330 4680 11410 4760
rect -360 4280 -200 4440
rect 8620 3960 9260 4260
rect 9260 3960 9580 4260
rect 14640 2300 14960 2620
rect 40100 1700 40500 1900
rect -360 -180 -200 -20
rect 11090 840 11190 920
rect 8040 200 8340 280
rect 44600 540 44720 860
rect 45330 540 45520 860
rect 45440 390 45510 450
rect 45510 390 45610 450
rect 45440 380 45610 390
rect 45950 410 46030 490
rect 12020 -180 12780 100
rect 10040 -740 10160 -420
rect 10500 -700 10620 -440
rect 10880 -890 10950 -830
rect 10950 -890 11050 -830
rect 10880 -900 11050 -890
rect 11210 -870 11290 -790
rect 45050 40 45190 150
rect 45770 110 45850 190
rect 45070 -340 45180 -210
rect 45880 -290 45960 -210
rect 45440 -622 45510 -562
rect 45510 -622 45610 -562
rect 45440 -632 45610 -622
rect 45770 -602 45850 -522
rect 2620 -4280 2700 -4120
rect 10490 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 14640 -1360 14960 -1040
rect 40100 -1100 40500 -900
rect 45050 -972 45190 -862
rect 45950 -902 46030 -822
rect 10510 -1620 10620 -1490
rect 11320 -1570 11400 -1490
rect 8120 -5580 8280 -5420
rect 50690 -5640 50910 -5540
rect 54440 -6850 54510 -6720
<< metal4 >>
rect 3400 13800 4600 14000
rect 3400 13200 3600 13800
rect 4400 13200 6600 13800
rect 14200 13700 44860 13800
rect 3400 13000 4600 13200
rect 14200 12600 43100 13700
rect 44100 12600 44860 13700
rect 14200 12500 44860 12600
rect -360 10300 5140 10460
rect -360 4460 -200 10300
rect 54300 10250 54520 10260
rect 54300 10180 54440 10250
rect 54290 10120 54440 10180
rect 54510 10120 54520 10250
rect 54290 10110 54520 10120
rect 0 9800 100 10100
rect 200 9800 300 10100
rect 400 9800 500 10100
rect 600 9900 900 10100
rect 600 9800 700 9900
rect 800 9800 900 9900
rect 50145 10025 53285 10095
rect 50145 9050 50215 10025
rect 50145 9040 50920 9050
rect 50145 8980 50690 9040
rect 50680 8940 50690 8980
rect 50910 8940 50920 9040
rect 50680 8930 50920 8940
rect 40000 6100 45100 6200
rect 40000 5500 40100 6100
rect 41100 5500 45100 6100
rect 40000 5400 45100 5500
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11060 4460 11120 4820
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11180 4580 11240 4820
rect 11320 4760 11990 4770
rect 11320 4680 11330 4760
rect 11410 4680 11990 4760
rect 11320 4670 11990 4680
rect 11180 4520 11620 4580
rect -380 4440 -180 4460
rect -380 4280 -360 4440
rect -200 4280 -180 4440
rect 11060 4400 11490 4460
rect -380 4260 -180 4280
rect 8600 4260 9600 4280
rect 8600 3960 8620 4260
rect 9580 3960 9600 4260
rect 8600 3940 9600 3960
rect 10500 920 11210 940
rect 10500 840 11090 920
rect 11190 840 11210 920
rect 10500 820 11210 840
rect 8020 280 8360 300
rect 8020 200 8040 280
rect 8020 20 8060 200
rect 8340 20 8360 280
rect 8020 0 8360 20
rect -380 -20 -180 0
rect -380 -180 -360 -20
rect -200 -180 -180 -20
rect -380 -200 -180 -180
rect -360 -6920 -200 -200
rect 9900 -420 10180 -400
rect 10500 -420 10620 820
rect 11430 680 11490 4400
rect 11240 620 11490 680
rect 9900 -740 9920 -420
rect 10160 -740 10180 -420
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 9900 -760 10180 -740
rect 11240 -780 11300 620
rect 11560 560 11620 4520
rect 11200 -790 11300 -780
rect 11200 -820 11210 -790
rect 10870 -830 11210 -820
rect 10870 -900 10880 -830
rect 11050 -870 11210 -830
rect 11290 -870 11300 -790
rect 11050 -880 11300 -870
rect 11420 500 11620 560
rect 11050 -900 11060 -880
rect 10870 -910 11060 -900
rect 11420 -1080 11480 500
rect 11890 370 11990 4670
rect 14600 2620 15000 2660
rect 14600 2300 14640 2620
rect 14960 2300 15000 2620
rect 14600 2220 15000 2300
rect 14800 1700 15100 2200
rect 40000 2100 40600 2200
rect 40000 1700 40100 2100
rect 40500 1885 40600 2100
rect 40500 1700 45540 1885
rect 40000 1655 45540 1700
rect 40000 1600 40600 1655
rect 44460 860 44740 880
rect 44460 540 44480 860
rect 44720 540 44740 860
rect 44460 520 44740 540
rect 45310 860 45540 1655
rect 45310 540 45330 860
rect 45520 540 45540 860
rect 45310 520 45540 540
rect 45940 490 46040 500
rect 45940 460 45950 490
rect 45430 450 45950 460
rect 45430 380 45440 450
rect 45610 410 45950 450
rect 46030 410 46040 490
rect 45610 400 46040 410
rect 45610 380 45620 400
rect 45430 370 45620 380
rect 11380 -1090 11480 -1080
rect 11380 -1120 11390 -1090
rect 10480 -1130 11390 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1170 11390 -1130
rect 11470 -1170 11480 -1090
rect 10630 -1180 11480 -1170
rect 11790 270 11990 370
rect 10630 -1240 10640 -1180
rect 10480 -1250 10640 -1240
rect 11790 -1480 11890 270
rect 45760 190 45860 200
rect 45760 160 45770 190
rect 45040 150 45770 160
rect 11980 100 12820 120
rect 11980 -180 12020 100
rect 12780 -180 12820 100
rect 45040 40 45050 150
rect 45190 110 45770 150
rect 45850 110 45860 190
rect 45190 100 45860 110
rect 45190 40 45200 100
rect 45040 30 45200 40
rect 11980 -200 12820 -180
rect 41410 -200 41510 -190
rect 41410 -210 46140 -200
rect 41410 -300 45070 -210
rect 40000 -900 40600 -800
rect 14600 -1040 15000 -1000
rect 14600 -1360 14640 -1040
rect 14960 -1360 15000 -1040
rect 14600 -1400 15000 -1360
rect 40000 -1300 40100 -900
rect 40500 -1300 40600 -900
rect 40000 -1400 40600 -1300
rect 10500 -1490 11890 -1480
rect 10500 -1620 10510 -1490
rect 10620 -1570 11320 -1490
rect 11400 -1570 11890 -1490
rect 10620 -1580 11890 -1570
rect 10620 -1620 10630 -1580
rect 10500 -1630 10630 -1620
rect 11790 -1690 11890 -1580
rect 41410 -1610 41510 -300
rect 45060 -340 45070 -300
rect 45180 -290 45880 -210
rect 45960 -290 46140 -210
rect 45180 -300 46140 -290
rect 45180 -340 45190 -300
rect 45060 -350 45190 -340
rect 45760 -522 45860 -512
rect 45760 -552 45770 -522
rect 45430 -562 45770 -552
rect 45430 -632 45440 -562
rect 45610 -602 45770 -562
rect 45850 -602 45860 -522
rect 45610 -612 45860 -602
rect 45610 -632 45620 -612
rect 45430 -642 45620 -632
rect 45940 -822 46040 -812
rect 45940 -852 45950 -822
rect 45040 -862 45950 -852
rect 45040 -972 45050 -862
rect 45190 -902 45950 -862
rect 46030 -902 46040 -822
rect 45190 -910 46040 -902
rect 45190 -912 46000 -910
rect 45190 -972 45200 -912
rect 45040 -982 45200 -972
rect 11790 -1790 15230 -1690
rect 2600 -4120 7000 -4100
rect 2600 -4280 2620 -4120
rect 2700 -4280 7000 -4120
rect 2600 -4300 7000 -4280
rect 6800 -5400 7000 -4300
rect 6800 -5420 8300 -5400
rect 6800 -5580 8120 -5420
rect 8280 -5580 8300 -5420
rect 6800 -5600 8300 -5580
rect 0 -6600 100 -6400
rect 200 -6600 300 -6400
rect 0 -6700 300 -6600
rect 400 -6700 500 -6400
rect 600 -6700 700 -6400
rect 800 -6600 1100 -6400
rect 800 -6700 900 -6600
rect 1000 -6700 1100 -6600
rect -360 -7080 5200 -6920
rect 15130 -7690 15230 -1790
rect 39330 -1710 41510 -1610
rect 39330 -7690 39430 -1710
rect 40000 -2100 44540 -2000
rect 40000 -2700 40100 -2100
rect 41100 -2700 44540 -2100
rect 40000 -2800 44540 -2700
rect 50680 -5540 50920 -5530
rect 50680 -5580 50690 -5540
rect 50145 -5640 50690 -5580
rect 50910 -5640 50920 -5540
rect 50145 -5650 50920 -5640
rect 50145 -6625 50215 -5650
rect 50145 -6695 53285 -6625
rect 54290 -6720 54520 -6710
rect 54290 -6780 54440 -6720
rect 54300 -6850 54440 -6780
rect 54510 -6850 54520 -6720
rect 54300 -6860 54520 -6850
rect 15130 -7790 39430 -7690
rect 14200 -9200 45000 -9100
rect 3400 -9800 4600 -9600
rect 3400 -10400 3600 -9800
rect 4400 -10400 6600 -9800
rect 14200 -10300 43100 -9200
rect 44100 -10300 45000 -9200
rect 14200 -10400 45000 -10300
rect 3400 -10600 4600 -10400
<< via4 >>
rect 3600 13200 4400 13800
rect 43100 12600 44100 13700
rect 40100 5500 41100 6100
rect 8640 3960 9560 4260
rect 8060 200 8340 260
rect 8060 20 8340 200
rect 9920 -740 10040 -420
rect 10040 -740 10160 -420
rect 40100 1900 40500 2100
rect 40100 1700 40500 1900
rect 44480 540 44600 860
rect 44600 540 44720 860
rect 12020 -180 12780 100
rect 40100 -1100 40500 -900
rect 40100 -1300 40500 -1100
rect 40100 -2700 41100 -2100
rect 3600 -10400 4400 -9800
rect 43100 -10300 44100 -9200
<< metal5 >>
rect 3400 13800 4600 15000
rect 3400 13200 3600 13800
rect 4400 13200 4600 13800
rect 3400 5400 4600 13200
rect 12000 5400 13200 15000
rect 3400 4800 9600 5400
rect 8600 4260 9600 4800
rect 8600 3960 8640 4260
rect 9560 3960 9600 4260
rect 8600 300 9600 3960
rect 8020 260 9600 300
rect 8020 20 8060 260
rect 8340 20 9600 260
rect 8020 -20 9600 20
rect 8600 -380 9600 -20
rect 11600 5000 13200 5400
rect 40000 6100 41200 15000
rect 40000 5500 40100 6100
rect 41100 5500 41200 6100
rect 11600 120 12800 5000
rect 40000 2100 41200 5500
rect 40000 1700 40100 2100
rect 40500 1700 41200 2100
rect 11600 100 12820 120
rect 11600 -180 12020 100
rect 12780 -180 12820 100
rect 11600 -200 12820 -180
rect 8600 -420 10200 -380
rect 8600 -740 9920 -420
rect 10160 -740 10200 -420
rect 8600 -780 10200 -740
rect 8600 -1000 9600 -780
rect 3400 -1600 9600 -1000
rect 11600 -1600 12800 -200
rect 40000 -900 41200 1700
rect 40000 -1300 40100 -900
rect 40500 -1300 41200 -900
rect 3400 -9800 4600 -1600
rect 11600 -2000 13200 -1600
rect 3400 -10400 3600 -9800
rect 4400 -10400 4600 -9800
rect 3400 -13000 4600 -10400
rect 12000 -13000 13200 -2000
rect 40000 -2100 41200 -1300
rect 40000 -2700 40100 -2100
rect 41100 -2700 41200 -2100
rect 40000 -13000 41200 -2700
rect 43000 13700 44200 15000
rect 43000 12600 43100 13700
rect 44100 12600 44200 13700
rect 43000 900 44200 12600
rect 43000 860 44760 900
rect 43000 540 44480 860
rect 44720 540 44760 860
rect 43000 500 44760 540
rect 43000 -9200 44200 500
rect 43000 -10300 43100 -9200
rect 44100 -10300 44200 -9200
rect 43000 -13000 44200 -10300
<< comment >>
rect -102 3247 -92 3251
use cmota_gb_rp_gp  cmota_gb_rp_gp_0
timestamp 1672206111
transform -1 0 7802 0 -1 -9800
box -7000 -7800 2802 600
use cmota_gb_rp_gp  cmota_gb_rp_gp_1
timestamp 1672206111
transform -1 0 7802 0 1 13200
box -7000 -7800 2802 600
use cmota_gb_rp_gp  cmota_gb_rp_gp_2
timestamp 1672206111
transform 1 0 51540 0 -1 -9800
box -7000 -7800 2802 600
use cmota_gb_rp_gp  cmota_gb_rp_gp_3
timestamp 1672206111
transform 1 0 51540 0 1 13200
box -7000 -7800 2802 600
use isrc  isrc_0
timestamp 1671401643
transform 1 0 10508 0 1 -1702
box -200 1760 4090 5700
use sky130_fd_pr__res_xhigh_po_0p35_KD7HM5  sky130_fd_pr__res_xhigh_po_0p35_KD7HM5_0
timestamp 1671931150
transform 0 1 39845 -1 0 429
box -782 -648 782 648
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 0 -1 10792 1 0 -998
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1670771148
transform 0 -1 45352 1 0 -730
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1670771148
transform 0 -1 45352 1 0 282
box -38 -48 314 592
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 2135 0 -1 2212
box -38 -49 230 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_1
timestamp 1670771148
transform 1 0 3287 0 1 880
box -38 -49 230 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_2
timestamp 1670771148
transform 1 0 2135 0 1 2212
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 3191 0 1 880
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1670771148
transform 1 0 9815 0 1 2212
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1670771148
transform 1 0 2039 0 1 2212
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_4
timestamp 1670771148
transform 1 0 2039 0 -1 2212
box -38 -49 134 715
use sky130hd_esd  sky130hd_esd_0
timestamp 1671850507
transform 1 0 2243 0 1 918
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_1
timestamp 1671850507
transform 1 0 7746 0 -1 796
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_2
timestamp 1671850507
transform 1 0 1875 0 1 918
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_3
timestamp 1671850507
transform 0 -1 10780 -1 0 -94
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_4
timestamp 1671850507
transform 0 -1 10780 -1 0 -1106
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_5
timestamp 1671850507
transform 0 -1 10780 -1 0 -738
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_6
timestamp 1671850507
transform 1 0 1507 0 1 918
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_7
timestamp 1671850507
transform 0 -1 45340 -1 0 542
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_9
timestamp 1671850507
transform 0 -1 45340 -1 0 -470
box 222 -60 666 580
use sky130hd_esd  sky130hd_esd_10
timestamp 1671850507
transform 0 -1 45340 -1 0 174
box 222 -60 666 580
use swcap_array_1  swcap_array_1_0
timestamp 1671395052
transform 0 -1 37998 1 0 -171
box -6569 -1080 7773 23570
use twcon  twcon_0
timestamp 1671985581
transform 1 0 5207 0 1 880
box -5309 -1622 5030 3682
<< labels >>
rlabel metal3 1900 -9060 2000 -8860 1 CLKIN
port 6 n
rlabel metal3 40500 980 40530 1040 1 B0
port 8 n
rlabel metal3 40500 820 40530 880 1 B1
port 9 n
rlabel metal3 40500 650 40530 710 1 B2
port 10 n
rlabel metal3 40500 480 40530 540 1 B3
port 11 n
rlabel metal3 40500 310 40530 370 1 B4
port 12 n
rlabel metal3 40500 150 40530 210 1 B5
port 13 n
rlabel metal3 40500 -10 40530 50 1 B6
port 14 n
rlabel metal3 40500 -180 40530 -120 1 B7
port 15 n
rlabel metal5 3400 -13000 4600 -12400 1 VHI
port 16 n
rlabel metal5 12000 -13000 13200 -12400 1 VLO
port 17 n
rlabel metal4 14800 1700 15100 2200 1 VOUT
port 18 n
rlabel metal3 2420 -9060 2540 -8860 1 C50
port 4 n
rlabel metal3 2240 -9060 2360 -8860 1 C100
port 5 n
rlabel metal3 2780 -9060 2900 -8860 1 IREF
port 2 n
rlabel metal3 2600 -9060 2720 -8860 1 ULIM
port 3 n
rlabel metal3 2960 -9060 3080 -8860 1 OPAEN
port 21 n
rlabel metal3 10360 1890 10450 1960 1 GP
port 22 n
rlabel metal3 10390 1150 10440 1200 1 GN
port 23 n
rlabel metal4 -360 10300 -200 10460 1 LLIM_A
port 24 n
rlabel metal4 -360 -7080 -200 -6920 1 ULIM_A
port 25 n
rlabel metal2 5208 1750 5238 1786 1 MUX_OUT
port 26 n
rlabel metal2 8928 1252 8966 1302 1 UPDN
port 27 n
rlabel metal2 5046 1650 5084 1700 1 ENCLK
port 28 n
rlabel metal3 3140 -9060 3260 -8860 1 VREF_OPA
port 29 n
rlabel metal3 1360 -9060 1480 -8860 1 LLIM
port 7 n
rlabel metal3 1560 -9060 1660 -8860 1 RSTB
port 30 n
rlabel metal3 44510 30 44650 160 1 GATE1
rlabel metal3 44520 -970 44650 -860 1 GATE2
rlabel metal3 54530 10120 54620 10250 1 OUT1
rlabel metal3 54530 -6850 54620 -6720 1 OUT2
<< end >>
