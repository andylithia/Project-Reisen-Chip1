magic
tech sky130A
magscale 1 2
timestamp 1671820621
<< obsli1 >>
rect 1104 2159 158884 13617
<< obsm1 >>
rect 1104 960 159514 15088
<< metal2 >>
rect 9586 15200 9642 16000
rect 10138 15200 10194 16000
rect 10690 15200 10746 16000
rect 11242 15200 11298 16000
rect 11794 15200 11850 16000
rect 12346 15200 12402 16000
rect 12898 15200 12954 16000
rect 13450 15200 13506 16000
rect 14002 15200 14058 16000
rect 14554 15200 14610 16000
rect 15106 15200 15162 16000
rect 15658 15200 15714 16000
rect 16210 15200 16266 16000
rect 16762 15200 16818 16000
rect 17314 15200 17370 16000
rect 17866 15200 17922 16000
rect 18418 15200 18474 16000
rect 18970 15200 19026 16000
rect 19522 15200 19578 16000
rect 20074 15200 20130 16000
rect 20626 15200 20682 16000
rect 21178 15200 21234 16000
rect 21730 15200 21786 16000
rect 22282 15200 22338 16000
rect 22834 15200 22890 16000
rect 23386 15200 23442 16000
rect 23938 15200 23994 16000
rect 24490 15200 24546 16000
rect 25042 15200 25098 16000
rect 25594 15200 25650 16000
rect 26146 15200 26202 16000
rect 26698 15200 26754 16000
rect 27250 15200 27306 16000
rect 27802 15200 27858 16000
rect 28354 15200 28410 16000
rect 28906 15200 28962 16000
rect 29458 15200 29514 16000
rect 30010 15200 30066 16000
rect 30562 15200 30618 16000
rect 31114 15200 31170 16000
rect 31666 15200 31722 16000
rect 32218 15200 32274 16000
rect 32770 15200 32826 16000
rect 33322 15200 33378 16000
rect 33874 15200 33930 16000
rect 34426 15200 34482 16000
rect 34978 15200 35034 16000
rect 35530 15200 35586 16000
rect 36082 15200 36138 16000
rect 36634 15200 36690 16000
rect 37186 15200 37242 16000
rect 37738 15200 37794 16000
rect 38290 15200 38346 16000
rect 38842 15200 38898 16000
rect 39394 15200 39450 16000
rect 39946 15200 40002 16000
rect 40498 15200 40554 16000
rect 41050 15200 41106 16000
rect 41602 15200 41658 16000
rect 42154 15200 42210 16000
rect 42706 15200 42762 16000
rect 43258 15200 43314 16000
rect 43810 15200 43866 16000
rect 44362 15200 44418 16000
rect 44914 15200 44970 16000
rect 45466 15200 45522 16000
rect 46018 15200 46074 16000
rect 46570 15200 46626 16000
rect 47122 15200 47178 16000
rect 47674 15200 47730 16000
rect 48226 15200 48282 16000
rect 48778 15200 48834 16000
rect 49330 15200 49386 16000
rect 49882 15200 49938 16000
rect 50434 15200 50490 16000
rect 50986 15200 51042 16000
rect 51538 15200 51594 16000
rect 52090 15200 52146 16000
rect 52642 15200 52698 16000
rect 53194 15200 53250 16000
rect 53746 15200 53802 16000
rect 54298 15200 54354 16000
rect 54850 15200 54906 16000
rect 55402 15200 55458 16000
rect 55954 15200 56010 16000
rect 56506 15200 56562 16000
rect 57058 15200 57114 16000
rect 57610 15200 57666 16000
rect 58162 15200 58218 16000
rect 58714 15200 58770 16000
rect 59266 15200 59322 16000
rect 59818 15200 59874 16000
rect 60370 15200 60426 16000
rect 60922 15200 60978 16000
rect 61474 15200 61530 16000
rect 62026 15200 62082 16000
rect 62578 15200 62634 16000
rect 63130 15200 63186 16000
rect 63682 15200 63738 16000
rect 64234 15200 64290 16000
rect 64786 15200 64842 16000
rect 65338 15200 65394 16000
rect 65890 15200 65946 16000
rect 66442 15200 66498 16000
rect 66994 15200 67050 16000
rect 67546 15200 67602 16000
rect 68098 15200 68154 16000
rect 68650 15200 68706 16000
rect 69202 15200 69258 16000
rect 69754 15200 69810 16000
rect 70306 15200 70362 16000
rect 70858 15200 70914 16000
rect 71410 15200 71466 16000
rect 71962 15200 72018 16000
rect 72514 15200 72570 16000
rect 73066 15200 73122 16000
rect 73618 15200 73674 16000
rect 74170 15200 74226 16000
rect 74722 15200 74778 16000
rect 75274 15200 75330 16000
rect 75826 15200 75882 16000
rect 76378 15200 76434 16000
rect 76930 15200 76986 16000
rect 77482 15200 77538 16000
rect 78034 15200 78090 16000
rect 78586 15200 78642 16000
rect 79138 15200 79194 16000
rect 79690 15200 79746 16000
rect 80242 15200 80298 16000
rect 80794 15200 80850 16000
rect 81346 15200 81402 16000
rect 81898 15200 81954 16000
rect 82450 15200 82506 16000
rect 83002 15200 83058 16000
rect 83554 15200 83610 16000
rect 84106 15200 84162 16000
rect 84658 15200 84714 16000
rect 85210 15200 85266 16000
rect 85762 15200 85818 16000
rect 86314 15200 86370 16000
rect 86866 15200 86922 16000
rect 87418 15200 87474 16000
rect 87970 15200 88026 16000
rect 88522 15200 88578 16000
rect 89074 15200 89130 16000
rect 89626 15200 89682 16000
rect 90178 15200 90234 16000
rect 90730 15200 90786 16000
rect 91282 15200 91338 16000
rect 91834 15200 91890 16000
rect 92386 15200 92442 16000
rect 92938 15200 92994 16000
rect 93490 15200 93546 16000
rect 94042 15200 94098 16000
rect 94594 15200 94650 16000
rect 95146 15200 95202 16000
rect 95698 15200 95754 16000
rect 96250 15200 96306 16000
rect 96802 15200 96858 16000
rect 97354 15200 97410 16000
rect 97906 15200 97962 16000
rect 98458 15200 98514 16000
rect 99010 15200 99066 16000
rect 99562 15200 99618 16000
rect 100114 15200 100170 16000
rect 100666 15200 100722 16000
rect 101218 15200 101274 16000
rect 101770 15200 101826 16000
rect 102322 15200 102378 16000
rect 102874 15200 102930 16000
rect 103426 15200 103482 16000
rect 103978 15200 104034 16000
rect 104530 15200 104586 16000
rect 105082 15200 105138 16000
rect 105634 15200 105690 16000
rect 106186 15200 106242 16000
rect 106738 15200 106794 16000
rect 107290 15200 107346 16000
rect 107842 15200 107898 16000
rect 108394 15200 108450 16000
rect 108946 15200 109002 16000
rect 109498 15200 109554 16000
rect 110050 15200 110106 16000
rect 110602 15200 110658 16000
rect 111154 15200 111210 16000
rect 111706 15200 111762 16000
rect 112258 15200 112314 16000
rect 112810 15200 112866 16000
rect 113362 15200 113418 16000
rect 113914 15200 113970 16000
rect 114466 15200 114522 16000
rect 115018 15200 115074 16000
rect 115570 15200 115626 16000
rect 116122 15200 116178 16000
rect 116674 15200 116730 16000
rect 117226 15200 117282 16000
rect 117778 15200 117834 16000
rect 118330 15200 118386 16000
rect 118882 15200 118938 16000
rect 119434 15200 119490 16000
rect 119986 15200 120042 16000
rect 120538 15200 120594 16000
rect 121090 15200 121146 16000
rect 121642 15200 121698 16000
rect 122194 15200 122250 16000
rect 122746 15200 122802 16000
rect 123298 15200 123354 16000
rect 123850 15200 123906 16000
rect 124402 15200 124458 16000
rect 124954 15200 125010 16000
rect 125506 15200 125562 16000
rect 126058 15200 126114 16000
rect 126610 15200 126666 16000
rect 127162 15200 127218 16000
rect 127714 15200 127770 16000
rect 128266 15200 128322 16000
rect 128818 15200 128874 16000
rect 129370 15200 129426 16000
rect 129922 15200 129978 16000
rect 130474 15200 130530 16000
rect 131026 15200 131082 16000
rect 131578 15200 131634 16000
rect 132130 15200 132186 16000
rect 132682 15200 132738 16000
rect 133234 15200 133290 16000
rect 133786 15200 133842 16000
rect 134338 15200 134394 16000
rect 134890 15200 134946 16000
rect 135442 15200 135498 16000
rect 135994 15200 136050 16000
rect 136546 15200 136602 16000
rect 137098 15200 137154 16000
rect 137650 15200 137706 16000
rect 138202 15200 138258 16000
rect 138754 15200 138810 16000
rect 139306 15200 139362 16000
rect 139858 15200 139914 16000
rect 140410 15200 140466 16000
rect 140962 15200 141018 16000
rect 141514 15200 141570 16000
rect 142066 15200 142122 16000
rect 142618 15200 142674 16000
rect 143170 15200 143226 16000
rect 143722 15200 143778 16000
rect 144274 15200 144330 16000
rect 144826 15200 144882 16000
rect 145378 15200 145434 16000
rect 145930 15200 145986 16000
rect 146482 15200 146538 16000
rect 147034 15200 147090 16000
rect 147586 15200 147642 16000
rect 148138 15200 148194 16000
rect 148690 15200 148746 16000
rect 149242 15200 149298 16000
rect 149794 15200 149850 16000
rect 150346 15200 150402 16000
<< obsm2 >>
rect 1582 15144 9530 15314
rect 9698 15144 10082 15314
rect 10250 15144 10634 15314
rect 10802 15144 11186 15314
rect 11354 15144 11738 15314
rect 11906 15144 12290 15314
rect 12458 15144 12842 15314
rect 13010 15144 13394 15314
rect 13562 15144 13946 15314
rect 14114 15144 14498 15314
rect 14666 15144 15050 15314
rect 15218 15144 15602 15314
rect 15770 15144 16154 15314
rect 16322 15144 16706 15314
rect 16874 15144 17258 15314
rect 17426 15144 17810 15314
rect 17978 15144 18362 15314
rect 18530 15144 18914 15314
rect 19082 15144 19466 15314
rect 19634 15144 20018 15314
rect 20186 15144 20570 15314
rect 20738 15144 21122 15314
rect 21290 15144 21674 15314
rect 21842 15144 22226 15314
rect 22394 15144 22778 15314
rect 22946 15144 23330 15314
rect 23498 15144 23882 15314
rect 24050 15144 24434 15314
rect 24602 15144 24986 15314
rect 25154 15144 25538 15314
rect 25706 15144 26090 15314
rect 26258 15144 26642 15314
rect 26810 15144 27194 15314
rect 27362 15144 27746 15314
rect 27914 15144 28298 15314
rect 28466 15144 28850 15314
rect 29018 15144 29402 15314
rect 29570 15144 29954 15314
rect 30122 15144 30506 15314
rect 30674 15144 31058 15314
rect 31226 15144 31610 15314
rect 31778 15144 32162 15314
rect 32330 15144 32714 15314
rect 32882 15144 33266 15314
rect 33434 15144 33818 15314
rect 33986 15144 34370 15314
rect 34538 15144 34922 15314
rect 35090 15144 35474 15314
rect 35642 15144 36026 15314
rect 36194 15144 36578 15314
rect 36746 15144 37130 15314
rect 37298 15144 37682 15314
rect 37850 15144 38234 15314
rect 38402 15144 38786 15314
rect 38954 15144 39338 15314
rect 39506 15144 39890 15314
rect 40058 15144 40442 15314
rect 40610 15144 40994 15314
rect 41162 15144 41546 15314
rect 41714 15144 42098 15314
rect 42266 15144 42650 15314
rect 42818 15144 43202 15314
rect 43370 15144 43754 15314
rect 43922 15144 44306 15314
rect 44474 15144 44858 15314
rect 45026 15144 45410 15314
rect 45578 15144 45962 15314
rect 46130 15144 46514 15314
rect 46682 15144 47066 15314
rect 47234 15144 47618 15314
rect 47786 15144 48170 15314
rect 48338 15144 48722 15314
rect 48890 15144 49274 15314
rect 49442 15144 49826 15314
rect 49994 15144 50378 15314
rect 50546 15144 50930 15314
rect 51098 15144 51482 15314
rect 51650 15144 52034 15314
rect 52202 15144 52586 15314
rect 52754 15144 53138 15314
rect 53306 15144 53690 15314
rect 53858 15144 54242 15314
rect 54410 15144 54794 15314
rect 54962 15144 55346 15314
rect 55514 15144 55898 15314
rect 56066 15144 56450 15314
rect 56618 15144 57002 15314
rect 57170 15144 57554 15314
rect 57722 15144 58106 15314
rect 58274 15144 58658 15314
rect 58826 15144 59210 15314
rect 59378 15144 59762 15314
rect 59930 15144 60314 15314
rect 60482 15144 60866 15314
rect 61034 15144 61418 15314
rect 61586 15144 61970 15314
rect 62138 15144 62522 15314
rect 62690 15144 63074 15314
rect 63242 15144 63626 15314
rect 63794 15144 64178 15314
rect 64346 15144 64730 15314
rect 64898 15144 65282 15314
rect 65450 15144 65834 15314
rect 66002 15144 66386 15314
rect 66554 15144 66938 15314
rect 67106 15144 67490 15314
rect 67658 15144 68042 15314
rect 68210 15144 68594 15314
rect 68762 15144 69146 15314
rect 69314 15144 69698 15314
rect 69866 15144 70250 15314
rect 70418 15144 70802 15314
rect 70970 15144 71354 15314
rect 71522 15144 71906 15314
rect 72074 15144 72458 15314
rect 72626 15144 73010 15314
rect 73178 15144 73562 15314
rect 73730 15144 74114 15314
rect 74282 15144 74666 15314
rect 74834 15144 75218 15314
rect 75386 15144 75770 15314
rect 75938 15144 76322 15314
rect 76490 15144 76874 15314
rect 77042 15144 77426 15314
rect 77594 15144 77978 15314
rect 78146 15144 78530 15314
rect 78698 15144 79082 15314
rect 79250 15144 79634 15314
rect 79802 15144 80186 15314
rect 80354 15144 80738 15314
rect 80906 15144 81290 15314
rect 81458 15144 81842 15314
rect 82010 15144 82394 15314
rect 82562 15144 82946 15314
rect 83114 15144 83498 15314
rect 83666 15144 84050 15314
rect 84218 15144 84602 15314
rect 84770 15144 85154 15314
rect 85322 15144 85706 15314
rect 85874 15144 86258 15314
rect 86426 15144 86810 15314
rect 86978 15144 87362 15314
rect 87530 15144 87914 15314
rect 88082 15144 88466 15314
rect 88634 15144 89018 15314
rect 89186 15144 89570 15314
rect 89738 15144 90122 15314
rect 90290 15144 90674 15314
rect 90842 15144 91226 15314
rect 91394 15144 91778 15314
rect 91946 15144 92330 15314
rect 92498 15144 92882 15314
rect 93050 15144 93434 15314
rect 93602 15144 93986 15314
rect 94154 15144 94538 15314
rect 94706 15144 95090 15314
rect 95258 15144 95642 15314
rect 95810 15144 96194 15314
rect 96362 15144 96746 15314
rect 96914 15144 97298 15314
rect 97466 15144 97850 15314
rect 98018 15144 98402 15314
rect 98570 15144 98954 15314
rect 99122 15144 99506 15314
rect 99674 15144 100058 15314
rect 100226 15144 100610 15314
rect 100778 15144 101162 15314
rect 101330 15144 101714 15314
rect 101882 15144 102266 15314
rect 102434 15144 102818 15314
rect 102986 15144 103370 15314
rect 103538 15144 103922 15314
rect 104090 15144 104474 15314
rect 104642 15144 105026 15314
rect 105194 15144 105578 15314
rect 105746 15144 106130 15314
rect 106298 15144 106682 15314
rect 106850 15144 107234 15314
rect 107402 15144 107786 15314
rect 107954 15144 108338 15314
rect 108506 15144 108890 15314
rect 109058 15144 109442 15314
rect 109610 15144 109994 15314
rect 110162 15144 110546 15314
rect 110714 15144 111098 15314
rect 111266 15144 111650 15314
rect 111818 15144 112202 15314
rect 112370 15144 112754 15314
rect 112922 15144 113306 15314
rect 113474 15144 113858 15314
rect 114026 15144 114410 15314
rect 114578 15144 114962 15314
rect 115130 15144 115514 15314
rect 115682 15144 116066 15314
rect 116234 15144 116618 15314
rect 116786 15144 117170 15314
rect 117338 15144 117722 15314
rect 117890 15144 118274 15314
rect 118442 15144 118826 15314
rect 118994 15144 119378 15314
rect 119546 15144 119930 15314
rect 120098 15144 120482 15314
rect 120650 15144 121034 15314
rect 121202 15144 121586 15314
rect 121754 15144 122138 15314
rect 122306 15144 122690 15314
rect 122858 15144 123242 15314
rect 123410 15144 123794 15314
rect 123962 15144 124346 15314
rect 124514 15144 124898 15314
rect 125066 15144 125450 15314
rect 125618 15144 126002 15314
rect 126170 15144 126554 15314
rect 126722 15144 127106 15314
rect 127274 15144 127658 15314
rect 127826 15144 128210 15314
rect 128378 15144 128762 15314
rect 128930 15144 129314 15314
rect 129482 15144 129866 15314
rect 130034 15144 130418 15314
rect 130586 15144 130970 15314
rect 131138 15144 131522 15314
rect 131690 15144 132074 15314
rect 132242 15144 132626 15314
rect 132794 15144 133178 15314
rect 133346 15144 133730 15314
rect 133898 15144 134282 15314
rect 134450 15144 134834 15314
rect 135002 15144 135386 15314
rect 135554 15144 135938 15314
rect 136106 15144 136490 15314
rect 136658 15144 137042 15314
rect 137210 15144 137594 15314
rect 137762 15144 138146 15314
rect 138314 15144 138698 15314
rect 138866 15144 139250 15314
rect 139418 15144 139802 15314
rect 139970 15144 140354 15314
rect 140522 15144 140906 15314
rect 141074 15144 141458 15314
rect 141626 15144 142010 15314
rect 142178 15144 142562 15314
rect 142730 15144 143114 15314
rect 143282 15144 143666 15314
rect 143834 15144 144218 15314
rect 144386 15144 144770 15314
rect 144938 15144 145322 15314
rect 145490 15144 145874 15314
rect 146042 15144 146426 15314
rect 146594 15144 146978 15314
rect 147146 15144 147530 15314
rect 147698 15144 148082 15314
rect 148250 15144 148634 15314
rect 148802 15144 149186 15314
rect 149354 15144 149738 15314
rect 149906 15144 150290 15314
rect 150458 15144 159508 15314
rect 1582 954 159508 15144
<< metal3 >>
rect 0 13744 800 13864
rect 0 9800 800 9920
rect 159200 7896 160000 8016
rect 0 5856 800 5976
rect 0 1912 800 2032
<< obsm3 >>
rect 800 13944 159331 14517
rect 880 13664 159331 13944
rect 800 10000 159331 13664
rect 880 9720 159331 10000
rect 800 8096 159331 9720
rect 800 7816 159120 8096
rect 800 6056 159331 7816
rect 880 5776 159331 6056
rect 800 2112 159331 5776
rect 880 1832 159331 2112
rect 800 987 159331 1832
<< metal4 >>
rect 20666 2128 20986 13648
rect 40388 2128 40708 13648
rect 60111 2128 60431 13648
rect 79833 2128 80153 13648
rect 99556 2128 99876 13648
rect 119278 2128 119598 13648
rect 139001 2128 139321 13648
rect 158723 2128 159043 13648
<< obsm4 >>
rect 124259 13728 156893 14517
rect 124259 2048 138921 13728
rect 139401 2048 156893 13728
rect 124259 1123 156893 2048
<< labels >>
rlabel metal2 s 9586 15200 9642 16000 6 dq[0]
port 1 nsew signal output
rlabel metal2 s 64786 15200 64842 16000 6 dq[100]
port 2 nsew signal output
rlabel metal2 s 65338 15200 65394 16000 6 dq[101]
port 3 nsew signal output
rlabel metal2 s 65890 15200 65946 16000 6 dq[102]
port 4 nsew signal output
rlabel metal2 s 66442 15200 66498 16000 6 dq[103]
port 5 nsew signal output
rlabel metal2 s 66994 15200 67050 16000 6 dq[104]
port 6 nsew signal output
rlabel metal2 s 67546 15200 67602 16000 6 dq[105]
port 7 nsew signal output
rlabel metal2 s 68098 15200 68154 16000 6 dq[106]
port 8 nsew signal output
rlabel metal2 s 68650 15200 68706 16000 6 dq[107]
port 9 nsew signal output
rlabel metal2 s 69202 15200 69258 16000 6 dq[108]
port 10 nsew signal output
rlabel metal2 s 69754 15200 69810 16000 6 dq[109]
port 11 nsew signal output
rlabel metal2 s 15106 15200 15162 16000 6 dq[10]
port 12 nsew signal output
rlabel metal2 s 70306 15200 70362 16000 6 dq[110]
port 13 nsew signal output
rlabel metal2 s 70858 15200 70914 16000 6 dq[111]
port 14 nsew signal output
rlabel metal2 s 71410 15200 71466 16000 6 dq[112]
port 15 nsew signal output
rlabel metal2 s 71962 15200 72018 16000 6 dq[113]
port 16 nsew signal output
rlabel metal2 s 72514 15200 72570 16000 6 dq[114]
port 17 nsew signal output
rlabel metal2 s 73066 15200 73122 16000 6 dq[115]
port 18 nsew signal output
rlabel metal2 s 73618 15200 73674 16000 6 dq[116]
port 19 nsew signal output
rlabel metal2 s 74170 15200 74226 16000 6 dq[117]
port 20 nsew signal output
rlabel metal2 s 74722 15200 74778 16000 6 dq[118]
port 21 nsew signal output
rlabel metal2 s 75274 15200 75330 16000 6 dq[119]
port 22 nsew signal output
rlabel metal2 s 15658 15200 15714 16000 6 dq[11]
port 23 nsew signal output
rlabel metal2 s 75826 15200 75882 16000 6 dq[120]
port 24 nsew signal output
rlabel metal2 s 76378 15200 76434 16000 6 dq[121]
port 25 nsew signal output
rlabel metal2 s 76930 15200 76986 16000 6 dq[122]
port 26 nsew signal output
rlabel metal2 s 77482 15200 77538 16000 6 dq[123]
port 27 nsew signal output
rlabel metal2 s 78034 15200 78090 16000 6 dq[124]
port 28 nsew signal output
rlabel metal2 s 78586 15200 78642 16000 6 dq[125]
port 29 nsew signal output
rlabel metal2 s 79138 15200 79194 16000 6 dq[126]
port 30 nsew signal output
rlabel metal2 s 79690 15200 79746 16000 6 dq[127]
port 31 nsew signal output
rlabel metal2 s 80242 15200 80298 16000 6 dq[128]
port 32 nsew signal output
rlabel metal2 s 80794 15200 80850 16000 6 dq[129]
port 33 nsew signal output
rlabel metal2 s 16210 15200 16266 16000 6 dq[12]
port 34 nsew signal output
rlabel metal2 s 81346 15200 81402 16000 6 dq[130]
port 35 nsew signal output
rlabel metal2 s 81898 15200 81954 16000 6 dq[131]
port 36 nsew signal output
rlabel metal2 s 82450 15200 82506 16000 6 dq[132]
port 37 nsew signal output
rlabel metal2 s 83002 15200 83058 16000 6 dq[133]
port 38 nsew signal output
rlabel metal2 s 83554 15200 83610 16000 6 dq[134]
port 39 nsew signal output
rlabel metal2 s 84106 15200 84162 16000 6 dq[135]
port 40 nsew signal output
rlabel metal2 s 84658 15200 84714 16000 6 dq[136]
port 41 nsew signal output
rlabel metal2 s 85210 15200 85266 16000 6 dq[137]
port 42 nsew signal output
rlabel metal2 s 85762 15200 85818 16000 6 dq[138]
port 43 nsew signal output
rlabel metal2 s 86314 15200 86370 16000 6 dq[139]
port 44 nsew signal output
rlabel metal2 s 16762 15200 16818 16000 6 dq[13]
port 45 nsew signal output
rlabel metal2 s 86866 15200 86922 16000 6 dq[140]
port 46 nsew signal output
rlabel metal2 s 87418 15200 87474 16000 6 dq[141]
port 47 nsew signal output
rlabel metal2 s 87970 15200 88026 16000 6 dq[142]
port 48 nsew signal output
rlabel metal2 s 88522 15200 88578 16000 6 dq[143]
port 49 nsew signal output
rlabel metal2 s 89074 15200 89130 16000 6 dq[144]
port 50 nsew signal output
rlabel metal2 s 89626 15200 89682 16000 6 dq[145]
port 51 nsew signal output
rlabel metal2 s 90178 15200 90234 16000 6 dq[146]
port 52 nsew signal output
rlabel metal2 s 90730 15200 90786 16000 6 dq[147]
port 53 nsew signal output
rlabel metal2 s 91282 15200 91338 16000 6 dq[148]
port 54 nsew signal output
rlabel metal2 s 91834 15200 91890 16000 6 dq[149]
port 55 nsew signal output
rlabel metal2 s 17314 15200 17370 16000 6 dq[14]
port 56 nsew signal output
rlabel metal2 s 92386 15200 92442 16000 6 dq[150]
port 57 nsew signal output
rlabel metal2 s 92938 15200 92994 16000 6 dq[151]
port 58 nsew signal output
rlabel metal2 s 93490 15200 93546 16000 6 dq[152]
port 59 nsew signal output
rlabel metal2 s 94042 15200 94098 16000 6 dq[153]
port 60 nsew signal output
rlabel metal2 s 94594 15200 94650 16000 6 dq[154]
port 61 nsew signal output
rlabel metal2 s 95146 15200 95202 16000 6 dq[155]
port 62 nsew signal output
rlabel metal2 s 95698 15200 95754 16000 6 dq[156]
port 63 nsew signal output
rlabel metal2 s 96250 15200 96306 16000 6 dq[157]
port 64 nsew signal output
rlabel metal2 s 96802 15200 96858 16000 6 dq[158]
port 65 nsew signal output
rlabel metal2 s 97354 15200 97410 16000 6 dq[159]
port 66 nsew signal output
rlabel metal2 s 17866 15200 17922 16000 6 dq[15]
port 67 nsew signal output
rlabel metal2 s 97906 15200 97962 16000 6 dq[160]
port 68 nsew signal output
rlabel metal2 s 98458 15200 98514 16000 6 dq[161]
port 69 nsew signal output
rlabel metal2 s 99010 15200 99066 16000 6 dq[162]
port 70 nsew signal output
rlabel metal2 s 99562 15200 99618 16000 6 dq[163]
port 71 nsew signal output
rlabel metal2 s 100114 15200 100170 16000 6 dq[164]
port 72 nsew signal output
rlabel metal2 s 100666 15200 100722 16000 6 dq[165]
port 73 nsew signal output
rlabel metal2 s 101218 15200 101274 16000 6 dq[166]
port 74 nsew signal output
rlabel metal2 s 101770 15200 101826 16000 6 dq[167]
port 75 nsew signal output
rlabel metal2 s 102322 15200 102378 16000 6 dq[168]
port 76 nsew signal output
rlabel metal2 s 102874 15200 102930 16000 6 dq[169]
port 77 nsew signal output
rlabel metal2 s 18418 15200 18474 16000 6 dq[16]
port 78 nsew signal output
rlabel metal2 s 103426 15200 103482 16000 6 dq[170]
port 79 nsew signal output
rlabel metal2 s 103978 15200 104034 16000 6 dq[171]
port 80 nsew signal output
rlabel metal2 s 104530 15200 104586 16000 6 dq[172]
port 81 nsew signal output
rlabel metal2 s 105082 15200 105138 16000 6 dq[173]
port 82 nsew signal output
rlabel metal2 s 105634 15200 105690 16000 6 dq[174]
port 83 nsew signal output
rlabel metal2 s 106186 15200 106242 16000 6 dq[175]
port 84 nsew signal output
rlabel metal2 s 106738 15200 106794 16000 6 dq[176]
port 85 nsew signal output
rlabel metal2 s 107290 15200 107346 16000 6 dq[177]
port 86 nsew signal output
rlabel metal2 s 107842 15200 107898 16000 6 dq[178]
port 87 nsew signal output
rlabel metal2 s 108394 15200 108450 16000 6 dq[179]
port 88 nsew signal output
rlabel metal2 s 18970 15200 19026 16000 6 dq[17]
port 89 nsew signal output
rlabel metal2 s 108946 15200 109002 16000 6 dq[180]
port 90 nsew signal output
rlabel metal2 s 109498 15200 109554 16000 6 dq[181]
port 91 nsew signal output
rlabel metal2 s 110050 15200 110106 16000 6 dq[182]
port 92 nsew signal output
rlabel metal2 s 110602 15200 110658 16000 6 dq[183]
port 93 nsew signal output
rlabel metal2 s 111154 15200 111210 16000 6 dq[184]
port 94 nsew signal output
rlabel metal2 s 111706 15200 111762 16000 6 dq[185]
port 95 nsew signal output
rlabel metal2 s 112258 15200 112314 16000 6 dq[186]
port 96 nsew signal output
rlabel metal2 s 112810 15200 112866 16000 6 dq[187]
port 97 nsew signal output
rlabel metal2 s 113362 15200 113418 16000 6 dq[188]
port 98 nsew signal output
rlabel metal2 s 113914 15200 113970 16000 6 dq[189]
port 99 nsew signal output
rlabel metal2 s 19522 15200 19578 16000 6 dq[18]
port 100 nsew signal output
rlabel metal2 s 114466 15200 114522 16000 6 dq[190]
port 101 nsew signal output
rlabel metal2 s 115018 15200 115074 16000 6 dq[191]
port 102 nsew signal output
rlabel metal2 s 115570 15200 115626 16000 6 dq[192]
port 103 nsew signal output
rlabel metal2 s 116122 15200 116178 16000 6 dq[193]
port 104 nsew signal output
rlabel metal2 s 116674 15200 116730 16000 6 dq[194]
port 105 nsew signal output
rlabel metal2 s 117226 15200 117282 16000 6 dq[195]
port 106 nsew signal output
rlabel metal2 s 117778 15200 117834 16000 6 dq[196]
port 107 nsew signal output
rlabel metal2 s 118330 15200 118386 16000 6 dq[197]
port 108 nsew signal output
rlabel metal2 s 118882 15200 118938 16000 6 dq[198]
port 109 nsew signal output
rlabel metal2 s 119434 15200 119490 16000 6 dq[199]
port 110 nsew signal output
rlabel metal2 s 20074 15200 20130 16000 6 dq[19]
port 111 nsew signal output
rlabel metal2 s 10138 15200 10194 16000 6 dq[1]
port 112 nsew signal output
rlabel metal2 s 119986 15200 120042 16000 6 dq[200]
port 113 nsew signal output
rlabel metal2 s 120538 15200 120594 16000 6 dq[201]
port 114 nsew signal output
rlabel metal2 s 121090 15200 121146 16000 6 dq[202]
port 115 nsew signal output
rlabel metal2 s 121642 15200 121698 16000 6 dq[203]
port 116 nsew signal output
rlabel metal2 s 122194 15200 122250 16000 6 dq[204]
port 117 nsew signal output
rlabel metal2 s 122746 15200 122802 16000 6 dq[205]
port 118 nsew signal output
rlabel metal2 s 123298 15200 123354 16000 6 dq[206]
port 119 nsew signal output
rlabel metal2 s 123850 15200 123906 16000 6 dq[207]
port 120 nsew signal output
rlabel metal2 s 124402 15200 124458 16000 6 dq[208]
port 121 nsew signal output
rlabel metal2 s 124954 15200 125010 16000 6 dq[209]
port 122 nsew signal output
rlabel metal2 s 20626 15200 20682 16000 6 dq[20]
port 123 nsew signal output
rlabel metal2 s 125506 15200 125562 16000 6 dq[210]
port 124 nsew signal output
rlabel metal2 s 126058 15200 126114 16000 6 dq[211]
port 125 nsew signal output
rlabel metal2 s 126610 15200 126666 16000 6 dq[212]
port 126 nsew signal output
rlabel metal2 s 127162 15200 127218 16000 6 dq[213]
port 127 nsew signal output
rlabel metal2 s 127714 15200 127770 16000 6 dq[214]
port 128 nsew signal output
rlabel metal2 s 128266 15200 128322 16000 6 dq[215]
port 129 nsew signal output
rlabel metal2 s 128818 15200 128874 16000 6 dq[216]
port 130 nsew signal output
rlabel metal2 s 129370 15200 129426 16000 6 dq[217]
port 131 nsew signal output
rlabel metal2 s 129922 15200 129978 16000 6 dq[218]
port 132 nsew signal output
rlabel metal2 s 130474 15200 130530 16000 6 dq[219]
port 133 nsew signal output
rlabel metal2 s 21178 15200 21234 16000 6 dq[21]
port 134 nsew signal output
rlabel metal2 s 131026 15200 131082 16000 6 dq[220]
port 135 nsew signal output
rlabel metal2 s 131578 15200 131634 16000 6 dq[221]
port 136 nsew signal output
rlabel metal2 s 132130 15200 132186 16000 6 dq[222]
port 137 nsew signal output
rlabel metal2 s 132682 15200 132738 16000 6 dq[223]
port 138 nsew signal output
rlabel metal2 s 133234 15200 133290 16000 6 dq[224]
port 139 nsew signal output
rlabel metal2 s 133786 15200 133842 16000 6 dq[225]
port 140 nsew signal output
rlabel metal2 s 134338 15200 134394 16000 6 dq[226]
port 141 nsew signal output
rlabel metal2 s 134890 15200 134946 16000 6 dq[227]
port 142 nsew signal output
rlabel metal2 s 135442 15200 135498 16000 6 dq[228]
port 143 nsew signal output
rlabel metal2 s 135994 15200 136050 16000 6 dq[229]
port 144 nsew signal output
rlabel metal2 s 21730 15200 21786 16000 6 dq[22]
port 145 nsew signal output
rlabel metal2 s 136546 15200 136602 16000 6 dq[230]
port 146 nsew signal output
rlabel metal2 s 137098 15200 137154 16000 6 dq[231]
port 147 nsew signal output
rlabel metal2 s 137650 15200 137706 16000 6 dq[232]
port 148 nsew signal output
rlabel metal2 s 138202 15200 138258 16000 6 dq[233]
port 149 nsew signal output
rlabel metal2 s 138754 15200 138810 16000 6 dq[234]
port 150 nsew signal output
rlabel metal2 s 139306 15200 139362 16000 6 dq[235]
port 151 nsew signal output
rlabel metal2 s 139858 15200 139914 16000 6 dq[236]
port 152 nsew signal output
rlabel metal2 s 140410 15200 140466 16000 6 dq[237]
port 153 nsew signal output
rlabel metal2 s 140962 15200 141018 16000 6 dq[238]
port 154 nsew signal output
rlabel metal2 s 141514 15200 141570 16000 6 dq[239]
port 155 nsew signal output
rlabel metal2 s 22282 15200 22338 16000 6 dq[23]
port 156 nsew signal output
rlabel metal2 s 142066 15200 142122 16000 6 dq[240]
port 157 nsew signal output
rlabel metal2 s 142618 15200 142674 16000 6 dq[241]
port 158 nsew signal output
rlabel metal2 s 143170 15200 143226 16000 6 dq[242]
port 159 nsew signal output
rlabel metal2 s 143722 15200 143778 16000 6 dq[243]
port 160 nsew signal output
rlabel metal2 s 144274 15200 144330 16000 6 dq[244]
port 161 nsew signal output
rlabel metal2 s 144826 15200 144882 16000 6 dq[245]
port 162 nsew signal output
rlabel metal2 s 145378 15200 145434 16000 6 dq[246]
port 163 nsew signal output
rlabel metal2 s 145930 15200 145986 16000 6 dq[247]
port 164 nsew signal output
rlabel metal2 s 146482 15200 146538 16000 6 dq[248]
port 165 nsew signal output
rlabel metal2 s 147034 15200 147090 16000 6 dq[249]
port 166 nsew signal output
rlabel metal2 s 22834 15200 22890 16000 6 dq[24]
port 167 nsew signal output
rlabel metal2 s 147586 15200 147642 16000 6 dq[250]
port 168 nsew signal output
rlabel metal2 s 148138 15200 148194 16000 6 dq[251]
port 169 nsew signal output
rlabel metal2 s 148690 15200 148746 16000 6 dq[252]
port 170 nsew signal output
rlabel metal2 s 149242 15200 149298 16000 6 dq[253]
port 171 nsew signal output
rlabel metal2 s 149794 15200 149850 16000 6 dq[254]
port 172 nsew signal output
rlabel metal2 s 150346 15200 150402 16000 6 dq[255]
port 173 nsew signal output
rlabel metal2 s 23386 15200 23442 16000 6 dq[25]
port 174 nsew signal output
rlabel metal2 s 23938 15200 23994 16000 6 dq[26]
port 175 nsew signal output
rlabel metal2 s 24490 15200 24546 16000 6 dq[27]
port 176 nsew signal output
rlabel metal2 s 25042 15200 25098 16000 6 dq[28]
port 177 nsew signal output
rlabel metal2 s 25594 15200 25650 16000 6 dq[29]
port 178 nsew signal output
rlabel metal2 s 10690 15200 10746 16000 6 dq[2]
port 179 nsew signal output
rlabel metal2 s 26146 15200 26202 16000 6 dq[30]
port 180 nsew signal output
rlabel metal2 s 26698 15200 26754 16000 6 dq[31]
port 181 nsew signal output
rlabel metal2 s 27250 15200 27306 16000 6 dq[32]
port 182 nsew signal output
rlabel metal2 s 27802 15200 27858 16000 6 dq[33]
port 183 nsew signal output
rlabel metal2 s 28354 15200 28410 16000 6 dq[34]
port 184 nsew signal output
rlabel metal2 s 28906 15200 28962 16000 6 dq[35]
port 185 nsew signal output
rlabel metal2 s 29458 15200 29514 16000 6 dq[36]
port 186 nsew signal output
rlabel metal2 s 30010 15200 30066 16000 6 dq[37]
port 187 nsew signal output
rlabel metal2 s 30562 15200 30618 16000 6 dq[38]
port 188 nsew signal output
rlabel metal2 s 31114 15200 31170 16000 6 dq[39]
port 189 nsew signal output
rlabel metal2 s 11242 15200 11298 16000 6 dq[3]
port 190 nsew signal output
rlabel metal2 s 31666 15200 31722 16000 6 dq[40]
port 191 nsew signal output
rlabel metal2 s 32218 15200 32274 16000 6 dq[41]
port 192 nsew signal output
rlabel metal2 s 32770 15200 32826 16000 6 dq[42]
port 193 nsew signal output
rlabel metal2 s 33322 15200 33378 16000 6 dq[43]
port 194 nsew signal output
rlabel metal2 s 33874 15200 33930 16000 6 dq[44]
port 195 nsew signal output
rlabel metal2 s 34426 15200 34482 16000 6 dq[45]
port 196 nsew signal output
rlabel metal2 s 34978 15200 35034 16000 6 dq[46]
port 197 nsew signal output
rlabel metal2 s 35530 15200 35586 16000 6 dq[47]
port 198 nsew signal output
rlabel metal2 s 36082 15200 36138 16000 6 dq[48]
port 199 nsew signal output
rlabel metal2 s 36634 15200 36690 16000 6 dq[49]
port 200 nsew signal output
rlabel metal2 s 11794 15200 11850 16000 6 dq[4]
port 201 nsew signal output
rlabel metal2 s 37186 15200 37242 16000 6 dq[50]
port 202 nsew signal output
rlabel metal2 s 37738 15200 37794 16000 6 dq[51]
port 203 nsew signal output
rlabel metal2 s 38290 15200 38346 16000 6 dq[52]
port 204 nsew signal output
rlabel metal2 s 38842 15200 38898 16000 6 dq[53]
port 205 nsew signal output
rlabel metal2 s 39394 15200 39450 16000 6 dq[54]
port 206 nsew signal output
rlabel metal2 s 39946 15200 40002 16000 6 dq[55]
port 207 nsew signal output
rlabel metal2 s 40498 15200 40554 16000 6 dq[56]
port 208 nsew signal output
rlabel metal2 s 41050 15200 41106 16000 6 dq[57]
port 209 nsew signal output
rlabel metal2 s 41602 15200 41658 16000 6 dq[58]
port 210 nsew signal output
rlabel metal2 s 42154 15200 42210 16000 6 dq[59]
port 211 nsew signal output
rlabel metal2 s 12346 15200 12402 16000 6 dq[5]
port 212 nsew signal output
rlabel metal2 s 42706 15200 42762 16000 6 dq[60]
port 213 nsew signal output
rlabel metal2 s 43258 15200 43314 16000 6 dq[61]
port 214 nsew signal output
rlabel metal2 s 43810 15200 43866 16000 6 dq[62]
port 215 nsew signal output
rlabel metal2 s 44362 15200 44418 16000 6 dq[63]
port 216 nsew signal output
rlabel metal2 s 44914 15200 44970 16000 6 dq[64]
port 217 nsew signal output
rlabel metal2 s 45466 15200 45522 16000 6 dq[65]
port 218 nsew signal output
rlabel metal2 s 46018 15200 46074 16000 6 dq[66]
port 219 nsew signal output
rlabel metal2 s 46570 15200 46626 16000 6 dq[67]
port 220 nsew signal output
rlabel metal2 s 47122 15200 47178 16000 6 dq[68]
port 221 nsew signal output
rlabel metal2 s 47674 15200 47730 16000 6 dq[69]
port 222 nsew signal output
rlabel metal2 s 12898 15200 12954 16000 6 dq[6]
port 223 nsew signal output
rlabel metal2 s 48226 15200 48282 16000 6 dq[70]
port 224 nsew signal output
rlabel metal2 s 48778 15200 48834 16000 6 dq[71]
port 225 nsew signal output
rlabel metal2 s 49330 15200 49386 16000 6 dq[72]
port 226 nsew signal output
rlabel metal2 s 49882 15200 49938 16000 6 dq[73]
port 227 nsew signal output
rlabel metal2 s 50434 15200 50490 16000 6 dq[74]
port 228 nsew signal output
rlabel metal2 s 50986 15200 51042 16000 6 dq[75]
port 229 nsew signal output
rlabel metal2 s 51538 15200 51594 16000 6 dq[76]
port 230 nsew signal output
rlabel metal2 s 52090 15200 52146 16000 6 dq[77]
port 231 nsew signal output
rlabel metal2 s 52642 15200 52698 16000 6 dq[78]
port 232 nsew signal output
rlabel metal2 s 53194 15200 53250 16000 6 dq[79]
port 233 nsew signal output
rlabel metal2 s 13450 15200 13506 16000 6 dq[7]
port 234 nsew signal output
rlabel metal2 s 53746 15200 53802 16000 6 dq[80]
port 235 nsew signal output
rlabel metal2 s 54298 15200 54354 16000 6 dq[81]
port 236 nsew signal output
rlabel metal2 s 54850 15200 54906 16000 6 dq[82]
port 237 nsew signal output
rlabel metal2 s 55402 15200 55458 16000 6 dq[83]
port 238 nsew signal output
rlabel metal2 s 55954 15200 56010 16000 6 dq[84]
port 239 nsew signal output
rlabel metal2 s 56506 15200 56562 16000 6 dq[85]
port 240 nsew signal output
rlabel metal2 s 57058 15200 57114 16000 6 dq[86]
port 241 nsew signal output
rlabel metal2 s 57610 15200 57666 16000 6 dq[87]
port 242 nsew signal output
rlabel metal2 s 58162 15200 58218 16000 6 dq[88]
port 243 nsew signal output
rlabel metal2 s 58714 15200 58770 16000 6 dq[89]
port 244 nsew signal output
rlabel metal2 s 14002 15200 14058 16000 6 dq[8]
port 245 nsew signal output
rlabel metal2 s 59266 15200 59322 16000 6 dq[90]
port 246 nsew signal output
rlabel metal2 s 59818 15200 59874 16000 6 dq[91]
port 247 nsew signal output
rlabel metal2 s 60370 15200 60426 16000 6 dq[92]
port 248 nsew signal output
rlabel metal2 s 60922 15200 60978 16000 6 dq[93]
port 249 nsew signal output
rlabel metal2 s 61474 15200 61530 16000 6 dq[94]
port 250 nsew signal output
rlabel metal2 s 62026 15200 62082 16000 6 dq[95]
port 251 nsew signal output
rlabel metal2 s 62578 15200 62634 16000 6 dq[96]
port 252 nsew signal output
rlabel metal2 s 63130 15200 63186 16000 6 dq[97]
port 253 nsew signal output
rlabel metal2 s 63682 15200 63738 16000 6 dq[98]
port 254 nsew signal output
rlabel metal2 s 64234 15200 64290 16000 6 dq[99]
port 255 nsew signal output
rlabel metal2 s 14554 15200 14610 16000 6 dq[9]
port 256 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 latch
port 257 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 rst_n
port 258 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 sclk
port 259 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 sdi
port 260 nsew signal input
rlabel metal3 s 159200 7896 160000 8016 6 sdo
port 261 nsew signal output
rlabel metal4 s 20666 2128 20986 13648 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 60111 2128 60431 13648 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 99556 2128 99876 13648 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 139001 2128 139321 13648 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 40388 2128 40708 13648 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 79833 2128 80153 13648 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 119278 2128 119598 13648 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 158723 2128 159043 13648 6 vssd1
port 263 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 160000 16000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4676046
string GDS_FILE /home/andylithia/openmpw/Project-Reisen-Chip1_digital/openlane/cfgsr/runs/22_12_23_13_34/results/signoff/cfgsr.magic.gds
string GDS_START 118736
<< end >>

