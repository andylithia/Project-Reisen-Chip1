// This is the unpowered netlist.
module cfgsr (latch,
    rst_n,
    sclk,
    sdi,
    sdo,
    dq);
 input latch;
 input rst_n;
 input sclk;
 input sdi;
 output sdo;
 output [255:0] dq;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire \sr[0] ;
 wire \sr[100] ;
 wire \sr[101] ;
 wire \sr[102] ;
 wire \sr[103] ;
 wire \sr[104] ;
 wire \sr[105] ;
 wire \sr[106] ;
 wire \sr[107] ;
 wire \sr[108] ;
 wire \sr[109] ;
 wire \sr[10] ;
 wire \sr[110] ;
 wire \sr[111] ;
 wire \sr[112] ;
 wire \sr[113] ;
 wire \sr[114] ;
 wire \sr[115] ;
 wire \sr[116] ;
 wire \sr[117] ;
 wire \sr[118] ;
 wire \sr[119] ;
 wire \sr[11] ;
 wire \sr[120] ;
 wire \sr[121] ;
 wire \sr[122] ;
 wire \sr[123] ;
 wire \sr[124] ;
 wire \sr[125] ;
 wire \sr[126] ;
 wire \sr[127] ;
 wire \sr[128] ;
 wire \sr[129] ;
 wire \sr[12] ;
 wire \sr[130] ;
 wire \sr[131] ;
 wire \sr[132] ;
 wire \sr[133] ;
 wire \sr[134] ;
 wire \sr[135] ;
 wire \sr[136] ;
 wire \sr[137] ;
 wire \sr[138] ;
 wire \sr[139] ;
 wire \sr[13] ;
 wire \sr[140] ;
 wire \sr[141] ;
 wire \sr[142] ;
 wire \sr[143] ;
 wire \sr[144] ;
 wire \sr[145] ;
 wire \sr[146] ;
 wire \sr[147] ;
 wire \sr[148] ;
 wire \sr[149] ;
 wire \sr[14] ;
 wire \sr[150] ;
 wire \sr[151] ;
 wire \sr[152] ;
 wire \sr[153] ;
 wire \sr[154] ;
 wire \sr[155] ;
 wire \sr[156] ;
 wire \sr[157] ;
 wire \sr[158] ;
 wire \sr[159] ;
 wire \sr[15] ;
 wire \sr[160] ;
 wire \sr[161] ;
 wire \sr[162] ;
 wire \sr[163] ;
 wire \sr[164] ;
 wire \sr[165] ;
 wire \sr[166] ;
 wire \sr[167] ;
 wire \sr[168] ;
 wire \sr[169] ;
 wire \sr[16] ;
 wire \sr[170] ;
 wire \sr[171] ;
 wire \sr[172] ;
 wire \sr[173] ;
 wire \sr[174] ;
 wire \sr[175] ;
 wire \sr[176] ;
 wire \sr[177] ;
 wire \sr[178] ;
 wire \sr[179] ;
 wire \sr[17] ;
 wire \sr[180] ;
 wire \sr[181] ;
 wire \sr[182] ;
 wire \sr[183] ;
 wire \sr[184] ;
 wire \sr[185] ;
 wire \sr[186] ;
 wire \sr[187] ;
 wire \sr[188] ;
 wire \sr[189] ;
 wire \sr[18] ;
 wire \sr[190] ;
 wire \sr[191] ;
 wire \sr[192] ;
 wire \sr[193] ;
 wire \sr[194] ;
 wire \sr[195] ;
 wire \sr[196] ;
 wire \sr[197] ;
 wire \sr[198] ;
 wire \sr[199] ;
 wire \sr[19] ;
 wire \sr[1] ;
 wire \sr[200] ;
 wire \sr[201] ;
 wire \sr[202] ;
 wire \sr[203] ;
 wire \sr[204] ;
 wire \sr[205] ;
 wire \sr[206] ;
 wire \sr[207] ;
 wire \sr[208] ;
 wire \sr[209] ;
 wire \sr[20] ;
 wire \sr[210] ;
 wire \sr[211] ;
 wire \sr[212] ;
 wire \sr[213] ;
 wire \sr[214] ;
 wire \sr[215] ;
 wire \sr[216] ;
 wire \sr[217] ;
 wire \sr[218] ;
 wire \sr[219] ;
 wire \sr[21] ;
 wire \sr[220] ;
 wire \sr[221] ;
 wire \sr[222] ;
 wire \sr[223] ;
 wire \sr[224] ;
 wire \sr[225] ;
 wire \sr[226] ;
 wire \sr[227] ;
 wire \sr[228] ;
 wire \sr[229] ;
 wire \sr[22] ;
 wire \sr[230] ;
 wire \sr[231] ;
 wire \sr[232] ;
 wire \sr[233] ;
 wire \sr[234] ;
 wire \sr[235] ;
 wire \sr[236] ;
 wire \sr[237] ;
 wire \sr[238] ;
 wire \sr[239] ;
 wire \sr[23] ;
 wire \sr[240] ;
 wire \sr[241] ;
 wire \sr[242] ;
 wire \sr[243] ;
 wire \sr[244] ;
 wire \sr[245] ;
 wire \sr[246] ;
 wire \sr[247] ;
 wire \sr[248] ;
 wire \sr[249] ;
 wire \sr[24] ;
 wire \sr[250] ;
 wire \sr[251] ;
 wire \sr[252] ;
 wire \sr[253] ;
 wire \sr[254] ;
 wire \sr[25] ;
 wire \sr[26] ;
 wire \sr[27] ;
 wire \sr[28] ;
 wire \sr[29] ;
 wire \sr[2] ;
 wire \sr[30] ;
 wire \sr[31] ;
 wire \sr[32] ;
 wire \sr[33] ;
 wire \sr[34] ;
 wire \sr[35] ;
 wire \sr[36] ;
 wire \sr[37] ;
 wire \sr[38] ;
 wire \sr[39] ;
 wire \sr[3] ;
 wire \sr[40] ;
 wire \sr[41] ;
 wire \sr[42] ;
 wire \sr[43] ;
 wire \sr[44] ;
 wire \sr[45] ;
 wire \sr[46] ;
 wire \sr[47] ;
 wire \sr[48] ;
 wire \sr[49] ;
 wire \sr[4] ;
 wire \sr[50] ;
 wire \sr[51] ;
 wire \sr[52] ;
 wire \sr[53] ;
 wire \sr[54] ;
 wire \sr[55] ;
 wire \sr[56] ;
 wire \sr[57] ;
 wire \sr[58] ;
 wire \sr[59] ;
 wire \sr[5] ;
 wire \sr[60] ;
 wire \sr[61] ;
 wire \sr[62] ;
 wire \sr[63] ;
 wire \sr[64] ;
 wire \sr[65] ;
 wire \sr[66] ;
 wire \sr[67] ;
 wire \sr[68] ;
 wire \sr[69] ;
 wire \sr[6] ;
 wire \sr[70] ;
 wire \sr[71] ;
 wire \sr[72] ;
 wire \sr[73] ;
 wire \sr[74] ;
 wire \sr[75] ;
 wire \sr[76] ;
 wire \sr[77] ;
 wire \sr[78] ;
 wire \sr[79] ;
 wire \sr[7] ;
 wire \sr[80] ;
 wire \sr[81] ;
 wire \sr[82] ;
 wire \sr[83] ;
 wire \sr[84] ;
 wire \sr[85] ;
 wire \sr[86] ;
 wire \sr[87] ;
 wire \sr[88] ;
 wire \sr[89] ;
 wire \sr[8] ;
 wire \sr[90] ;
 wire \sr[91] ;
 wire \sr[92] ;
 wire \sr[93] ;
 wire \sr[94] ;
 wire \sr[95] ;
 wire \sr[96] ;
 wire \sr[97] ;
 wire \sr[98] ;
 wire \sr[99] ;
 wire \sr[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire clknet_leaf_0_sclk;
 wire clknet_leaf_1_sclk;
 wire clknet_leaf_2_sclk;
 wire clknet_leaf_3_sclk;
 wire clknet_leaf_4_sclk;
 wire clknet_leaf_5_sclk;
 wire clknet_leaf_6_sclk;
 wire clknet_leaf_7_sclk;
 wire clknet_leaf_8_sclk;
 wire clknet_leaf_9_sclk;
 wire clknet_leaf_10_sclk;
 wire clknet_0_sclk;
 wire clknet_1_0__leaf_sclk;
 wire clknet_1_1__leaf_sclk;

 sky130_fd_sc_hd__clkbuf_4 _0540_ (.A(net2),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _0541_ (.A(\sr[12] ),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _0542_ (.A(_0285_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_2 _0543_ (.A(_0284_),
    .X(_0286_));
 sky130_fd_sc_hd__and2_1 _0544_ (.A(_0286_),
    .B(\sr[13] ),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0545_ (.A(_0287_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _0546_ (.A(_0286_),
    .B(\sr[14] ),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0547_ (.A(_0288_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _0548_ (.A(_0286_),
    .B(\sr[15] ),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0549_ (.A(_0289_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _0550_ (.A(_0286_),
    .B(\sr[16] ),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0551_ (.A(_0290_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _0552_ (.A(_0286_),
    .B(\sr[17] ),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0553_ (.A(_0291_),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _0554_ (.A(_0286_),
    .B(\sr[18] ),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0555_ (.A(_0292_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _0556_ (.A(_0286_),
    .B(\sr[19] ),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0557_ (.A(_0293_),
    .X(_0064_));
 sky130_fd_sc_hd__and2_1 _0558_ (.A(_0286_),
    .B(\sr[20] ),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0559_ (.A(_0294_),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _0560_ (.A(_0286_),
    .B(\sr[21] ),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0295_),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _0562_ (.A(_0286_),
    .B(\sr[22] ),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(_0296_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_2 _0564_ (.A(_0284_),
    .X(_0297_));
 sky130_fd_sc_hd__and2_1 _0565_ (.A(_0297_),
    .B(\sr[23] ),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0566_ (.A(_0298_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _0567_ (.A(_0297_),
    .B(\sr[24] ),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0568_ (.A(_0299_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _0569_ (.A(_0297_),
    .B(\sr[25] ),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _0570_ (.A(_0300_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _0571_ (.A(_0297_),
    .B(\sr[26] ),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0572_ (.A(_0301_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _0573_ (.A(_0297_),
    .B(\sr[27] ),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _0574_ (.A(_0302_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _0575_ (.A(_0297_),
    .B(\sr[28] ),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _0576_ (.A(_0303_),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _0577_ (.A(_0297_),
    .B(\sr[29] ),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0578_ (.A(_0304_),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _0579_ (.A(_0297_),
    .B(\sr[30] ),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0580_ (.A(_0305_),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _0581_ (.A(_0297_),
    .B(\sr[31] ),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _0582_ (.A(_0306_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _0583_ (.A(_0297_),
    .B(\sr[32] ),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _0584_ (.A(_0307_),
    .X(_0077_));
 sky130_fd_sc_hd__buf_2 _0585_ (.A(_0284_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _0586_ (.A(_0308_),
    .B(\sr[33] ),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _0587_ (.A(_0309_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _0588_ (.A(_0308_),
    .B(\sr[34] ),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0589_ (.A(_0310_),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _0590_ (.A(_0308_),
    .B(\sr[35] ),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _0591_ (.A(_0311_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _0592_ (.A(_0308_),
    .B(\sr[36] ),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0593_ (.A(_0312_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _0594_ (.A(_0308_),
    .B(\sr[37] ),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0313_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _0596_ (.A(_0308_),
    .B(\sr[38] ),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0314_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _0598_ (.A(_0308_),
    .B(\sr[39] ),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _0599_ (.A(_0315_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _0600_ (.A(_0308_),
    .B(\sr[40] ),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _0601_ (.A(_0316_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _0602_ (.A(_0308_),
    .B(\sr[41] ),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(_0317_),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _0604_ (.A(_0308_),
    .B(\sr[42] ),
    .X(_0318_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0605_ (.A(_0318_),
    .X(_0087_));
 sky130_fd_sc_hd__buf_2 _0606_ (.A(_0284_),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _0607_ (.A(_0319_),
    .B(\sr[43] ),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(_0320_),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _0609_ (.A(_0319_),
    .B(\sr[44] ),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0610_ (.A(_0321_),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _0611_ (.A(_0319_),
    .B(\sr[45] ),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0322_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _0613_ (.A(_0319_),
    .B(\sr[46] ),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(_0323_),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _0615_ (.A(_0319_),
    .B(\sr[47] ),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0324_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _0617_ (.A(_0319_),
    .B(\sr[48] ),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(_0325_),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _0619_ (.A(_0319_),
    .B(\sr[49] ),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(_0326_),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0621_ (.A(_0319_),
    .B(\sr[50] ),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0327_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _0623_ (.A(_0319_),
    .B(\sr[51] ),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0328_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(_0319_),
    .B(\sr[52] ),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(_0329_),
    .X(_0097_));
 sky130_fd_sc_hd__buf_4 _0627_ (.A(net2),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_4 _0628_ (.A(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _0629_ (.A(_0331_),
    .B(\sr[53] ),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0630_ (.A(_0332_),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _0631_ (.A(_0331_),
    .B(\sr[54] ),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0333_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0633_ (.A(_0331_),
    .B(\sr[55] ),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _0634_ (.A(_0334_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _0635_ (.A(_0331_),
    .B(\sr[56] ),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0636_ (.A(_0335_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _0637_ (.A(_0331_),
    .B(\sr[57] ),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(_0336_),
    .X(_0102_));
 sky130_fd_sc_hd__and2_1 _0639_ (.A(_0331_),
    .B(\sr[58] ),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0640_ (.A(_0337_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _0641_ (.A(_0331_),
    .B(\sr[59] ),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(_0338_),
    .X(_0104_));
 sky130_fd_sc_hd__and2_1 _0643_ (.A(_0331_),
    .B(\sr[60] ),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(_0339_),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _0645_ (.A(_0331_),
    .B(\sr[61] ),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0646_ (.A(_0340_),
    .X(_0106_));
 sky130_fd_sc_hd__and2_1 _0647_ (.A(_0331_),
    .B(\sr[62] ),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0341_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_4 _0649_ (.A(_0330_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _0650_ (.A(_0342_),
    .B(\sr[63] ),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0343_),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _0652_ (.A(_0342_),
    .B(\sr[64] ),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(_0344_),
    .X(_0109_));
 sky130_fd_sc_hd__and2_1 _0654_ (.A(_0342_),
    .B(\sr[65] ),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0655_ (.A(_0345_),
    .X(_0110_));
 sky130_fd_sc_hd__and2_1 _0656_ (.A(_0342_),
    .B(\sr[66] ),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(_0346_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _0658_ (.A(_0342_),
    .B(\sr[67] ),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0659_ (.A(_0347_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(_0342_),
    .B(\sr[68] ),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _0661_ (.A(_0348_),
    .X(_0113_));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(_0342_),
    .B(\sr[69] ),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0349_),
    .X(_0114_));
 sky130_fd_sc_hd__and2_1 _0664_ (.A(_0342_),
    .B(\sr[70] ),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0665_ (.A(_0350_),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0666_ (.A(_0342_),
    .B(\sr[71] ),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0667_ (.A(_0351_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _0668_ (.A(_0342_),
    .B(\sr[72] ),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _0669_ (.A(_0352_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _0670_ (.A(_0330_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(_0353_),
    .B(\sr[73] ),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0354_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _0673_ (.A(_0353_),
    .B(\sr[74] ),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0674_ (.A(_0355_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0675_ (.A(_0353_),
    .B(\sr[75] ),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0356_),
    .X(_0120_));
 sky130_fd_sc_hd__and2_1 _0677_ (.A(_0353_),
    .B(\sr[76] ),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0357_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _0679_ (.A(_0353_),
    .B(\sr[77] ),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(_0358_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _0681_ (.A(_0353_),
    .B(\sr[78] ),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0682_ (.A(_0359_),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _0683_ (.A(_0353_),
    .B(\sr[79] ),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0684_ (.A(_0360_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _0685_ (.A(_0353_),
    .B(\sr[80] ),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0686_ (.A(_0361_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _0687_ (.A(_0353_),
    .B(\sr[81] ),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0362_),
    .X(_0126_));
 sky130_fd_sc_hd__and2_1 _0689_ (.A(_0353_),
    .B(\sr[82] ),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0363_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_2 _0691_ (.A(_0330_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _0692_ (.A(_0364_),
    .B(\sr[83] ),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0365_),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _0694_ (.A(_0364_),
    .B(\sr[84] ),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0695_ (.A(_0366_),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _0696_ (.A(_0364_),
    .B(\sr[85] ),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0367_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _0698_ (.A(_0364_),
    .B(\sr[86] ),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(_0368_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_1 _0700_ (.A(_0364_),
    .B(\sr[87] ),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0701_ (.A(_0369_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_1 _0702_ (.A(_0364_),
    .B(\sr[88] ),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0370_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _0704_ (.A(_0364_),
    .B(\sr[89] ),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0705_ (.A(_0371_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _0706_ (.A(_0364_),
    .B(\sr[90] ),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _0707_ (.A(_0372_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(_0364_),
    .B(\sr[91] ),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0373_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _0710_ (.A(_0364_),
    .B(\sr[92] ),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0711_ (.A(_0374_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_2 _0712_ (.A(_0330_),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _0713_ (.A(_0375_),
    .B(\sr[93] ),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0376_),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _0715_ (.A(_0375_),
    .B(\sr[94] ),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0377_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(_0375_),
    .B(\sr[95] ),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _0718_ (.A(_0378_),
    .X(_0140_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(_0375_),
    .B(\sr[96] ),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0379_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _0721_ (.A(_0375_),
    .B(\sr[97] ),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0380_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_1 _0723_ (.A(_0375_),
    .B(\sr[98] ),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _0724_ (.A(_0381_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _0725_ (.A(_0375_),
    .B(\sr[99] ),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _0726_ (.A(_0382_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(_0375_),
    .B(\sr[100] ),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0728_ (.A(_0383_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _0729_ (.A(_0375_),
    .B(\sr[101] ),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0730_ (.A(_0384_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_1 _0731_ (.A(_0375_),
    .B(\sr[102] ),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _0732_ (.A(_0385_),
    .X(_0147_));
 sky130_fd_sc_hd__buf_2 _0733_ (.A(_0330_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0734_ (.A(_0386_),
    .B(\sr[103] ),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0387_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _0736_ (.A(_0386_),
    .B(\sr[104] ),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0388_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _0738_ (.A(_0386_),
    .B(\sr[105] ),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0389_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _0740_ (.A(_0386_),
    .B(\sr[106] ),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0390_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _0742_ (.A(_0386_),
    .B(\sr[107] ),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0391_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_1 _0744_ (.A(_0386_),
    .B(\sr[108] ),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _0745_ (.A(_0392_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _0746_ (.A(_0386_),
    .B(\sr[109] ),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0393_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _0748_ (.A(_0386_),
    .B(\sr[110] ),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _0749_ (.A(_0394_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _0750_ (.A(_0386_),
    .B(\sr[111] ),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0395_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _0752_ (.A(_0386_),
    .B(\sr[112] ),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0396_),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_4 _0754_ (.A(_0330_),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _0755_ (.A(_0397_),
    .B(\sr[113] ),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _0756_ (.A(_0398_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _0757_ (.A(_0397_),
    .B(\sr[114] ),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0758_ (.A(_0399_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _0759_ (.A(_0397_),
    .B(\sr[115] ),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _0760_ (.A(_0400_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _0761_ (.A(_0397_),
    .B(\sr[116] ),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0762_ (.A(_0401_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _0763_ (.A(_0397_),
    .B(\sr[117] ),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _0764_ (.A(_0402_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(_0397_),
    .B(\sr[118] ),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(_0403_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _0767_ (.A(_0397_),
    .B(\sr[119] ),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(_0404_),
    .X(_0164_));
 sky130_fd_sc_hd__and2_1 _0769_ (.A(_0397_),
    .B(\sr[120] ),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0405_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _0771_ (.A(_0397_),
    .B(\sr[121] ),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0406_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(_0397_),
    .B(\sr[122] ),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0774_ (.A(_0407_),
    .X(_0167_));
 sky130_fd_sc_hd__buf_2 _0775_ (.A(_0330_),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _0776_ (.A(_0408_),
    .B(\sr[123] ),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_2 _0777_ (.A(_0409_),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _0778_ (.A(_0408_),
    .B(\sr[124] ),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _0779_ (.A(_0410_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _0780_ (.A(_0408_),
    .B(\sr[125] ),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0781_ (.A(_0411_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _0782_ (.A(_0408_),
    .B(\sr[126] ),
    .X(_0412_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0783_ (.A(_0412_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _0784_ (.A(_0408_),
    .B(\sr[127] ),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_2 _0785_ (.A(_0413_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _0786_ (.A(_0408_),
    .B(\sr[128] ),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0414_),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _0788_ (.A(_0408_),
    .B(\sr[129] ),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0789_ (.A(_0415_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _0790_ (.A(_0408_),
    .B(\sr[130] ),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0791_ (.A(_0416_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _0792_ (.A(_0408_),
    .B(\sr[131] ),
    .X(_0417_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0793_ (.A(_0417_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(_0408_),
    .B(\sr[132] ),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0795_ (.A(_0418_),
    .X(_0177_));
 sky130_fd_sc_hd__buf_2 _0796_ (.A(_0330_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _0797_ (.A(_0419_),
    .B(\sr[133] ),
    .X(_0420_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0798_ (.A(_0420_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _0799_ (.A(_0419_),
    .B(\sr[134] ),
    .X(_0421_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0800_ (.A(_0421_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _0801_ (.A(_0419_),
    .B(\sr[135] ),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0422_),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _0803_ (.A(_0419_),
    .B(\sr[136] ),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0804_ (.A(_0423_),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _0805_ (.A(_0419_),
    .B(\sr[137] ),
    .X(_0424_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0806_ (.A(_0424_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(_0419_),
    .B(\sr[138] ),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(_0425_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _0809_ (.A(_0419_),
    .B(\sr[139] ),
    .X(_0426_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0810_ (.A(_0426_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_1 _0811_ (.A(_0419_),
    .B(\sr[140] ),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_2 _0812_ (.A(_0427_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _0813_ (.A(_0419_),
    .B(\sr[141] ),
    .X(_0428_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0814_ (.A(_0428_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _0815_ (.A(_0419_),
    .B(\sr[142] ),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_2 _0816_ (.A(_0429_),
    .X(_0187_));
 sky130_fd_sc_hd__buf_2 _0817_ (.A(_0330_),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _0818_ (.A(_0430_),
    .B(\sr[143] ),
    .X(_0431_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0819_ (.A(_0431_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(_0430_),
    .B(\sr[144] ),
    .X(_0432_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0821_ (.A(_0432_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _0822_ (.A(_0430_),
    .B(\sr[145] ),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_2 _0823_ (.A(_0433_),
    .X(_0190_));
 sky130_fd_sc_hd__and2_1 _0824_ (.A(_0430_),
    .B(\sr[146] ),
    .X(_0434_));
 sky130_fd_sc_hd__buf_2 _0825_ (.A(_0434_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0826_ (.A(_0430_),
    .B(\sr[147] ),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _0827_ (.A(_0435_),
    .X(_0192_));
 sky130_fd_sc_hd__and2_1 _0828_ (.A(_0430_),
    .B(\sr[148] ),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_2 _0829_ (.A(_0436_),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _0830_ (.A(_0430_),
    .B(\sr[149] ),
    .X(_0437_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0831_ (.A(_0437_),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _0832_ (.A(_0430_),
    .B(\sr[150] ),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_2 _0833_ (.A(_0438_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_1 _0834_ (.A(_0430_),
    .B(\sr[151] ),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _0835_ (.A(_0439_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _0836_ (.A(_0430_),
    .B(\sr[152] ),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _0837_ (.A(_0440_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_4 _0838_ (.A(net2),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_2 _0839_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _0840_ (.A(_0442_),
    .B(\sr[153] ),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0841_ (.A(_0443_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _0842_ (.A(_0442_),
    .B(\sr[154] ),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _0843_ (.A(_0444_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_1 _0844_ (.A(_0442_),
    .B(\sr[155] ),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0445_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _0846_ (.A(_0442_),
    .B(\sr[156] ),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0847_ (.A(_0446_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _0848_ (.A(_0442_),
    .B(\sr[157] ),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0849_ (.A(_0447_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0850_ (.A(_0442_),
    .B(\sr[158] ),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0851_ (.A(_0448_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _0852_ (.A(_0442_),
    .B(\sr[159] ),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0853_ (.A(_0449_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _0854_ (.A(_0442_),
    .B(\sr[160] ),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0855_ (.A(_0450_),
    .X(_0205_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(_0442_),
    .B(\sr[161] ),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0857_ (.A(_0451_),
    .X(_0206_));
 sky130_fd_sc_hd__and2_1 _0858_ (.A(_0442_),
    .B(\sr[162] ),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0859_ (.A(_0452_),
    .X(_0207_));
 sky130_fd_sc_hd__buf_2 _0860_ (.A(_0441_),
    .X(_0453_));
 sky130_fd_sc_hd__and2_1 _0861_ (.A(_0453_),
    .B(\sr[163] ),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0862_ (.A(_0454_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_1 _0863_ (.A(_0453_),
    .B(\sr[164] ),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0864_ (.A(_0455_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _0865_ (.A(_0453_),
    .B(\sr[165] ),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0866_ (.A(_0456_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_1 _0867_ (.A(_0453_),
    .B(\sr[166] ),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0868_ (.A(_0457_),
    .X(_0211_));
 sky130_fd_sc_hd__and2_1 _0869_ (.A(_0453_),
    .B(\sr[167] ),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0870_ (.A(_0458_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(_0453_),
    .B(\sr[168] ),
    .X(_0459_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0872_ (.A(_0459_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _0873_ (.A(_0453_),
    .B(\sr[169] ),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0460_),
    .X(_0214_));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(_0453_),
    .B(\sr[170] ),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_2 _0876_ (.A(_0461_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0453_),
    .B(\sr[171] ),
    .X(_0462_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0878_ (.A(_0462_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(_0453_),
    .B(\sr[172] ),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_2 _0880_ (.A(_0463_),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_4 _0881_ (.A(_0441_),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _0882_ (.A(_0464_),
    .B(\sr[173] ),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0883_ (.A(_0465_),
    .X(_0218_));
 sky130_fd_sc_hd__and2_1 _0884_ (.A(_0464_),
    .B(\sr[174] ),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0885_ (.A(_0466_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _0886_ (.A(_0464_),
    .B(\sr[175] ),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0887_ (.A(_0467_),
    .X(_0220_));
 sky130_fd_sc_hd__and2_1 _0888_ (.A(_0464_),
    .B(\sr[176] ),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0468_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(_0464_),
    .B(\sr[177] ),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0891_ (.A(_0469_),
    .X(_0222_));
 sky130_fd_sc_hd__and2_1 _0892_ (.A(_0464_),
    .B(\sr[178] ),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0470_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_1 _0894_ (.A(_0464_),
    .B(\sr[179] ),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0471_),
    .X(_0224_));
 sky130_fd_sc_hd__and2_1 _0896_ (.A(_0464_),
    .B(\sr[180] ),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0472_),
    .X(_0225_));
 sky130_fd_sc_hd__and2_1 _0898_ (.A(_0464_),
    .B(\sr[181] ),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0473_),
    .X(_0226_));
 sky130_fd_sc_hd__and2_1 _0900_ (.A(_0464_),
    .B(\sr[182] ),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0474_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_4 _0902_ (.A(_0441_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _0903_ (.A(_0475_),
    .B(\sr[183] ),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _0904_ (.A(_0476_),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _0905_ (.A(_0475_),
    .B(\sr[184] ),
    .X(_0477_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0906_ (.A(_0477_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_1 _0907_ (.A(_0475_),
    .B(\sr[185] ),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _0908_ (.A(_0478_),
    .X(_0230_));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(_0475_),
    .B(\sr[186] ),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _0910_ (.A(_0479_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(_0475_),
    .B(\sr[187] ),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _0912_ (.A(_0480_),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _0913_ (.A(_0475_),
    .B(\sr[188] ),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _0914_ (.A(_0481_),
    .X(_0233_));
 sky130_fd_sc_hd__and2_1 _0915_ (.A(_0475_),
    .B(\sr[189] ),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _0916_ (.A(_0482_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(_0475_),
    .B(\sr[190] ),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _0918_ (.A(_0483_),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _0919_ (.A(_0475_),
    .B(\sr[191] ),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _0920_ (.A(_0484_),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(_0475_),
    .B(\sr[192] ),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _0922_ (.A(_0485_),
    .X(_0237_));
 sky130_fd_sc_hd__buf_2 _0923_ (.A(_0441_),
    .X(_0486_));
 sky130_fd_sc_hd__and2_1 _0924_ (.A(_0486_),
    .B(\sr[193] ),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _0925_ (.A(_0487_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_1 _0926_ (.A(_0486_),
    .B(\sr[194] ),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _0927_ (.A(_0488_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _0928_ (.A(_0486_),
    .B(\sr[195] ),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _0929_ (.A(_0489_),
    .X(_0240_));
 sky130_fd_sc_hd__and2_1 _0930_ (.A(_0486_),
    .B(\sr[196] ),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _0931_ (.A(_0490_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _0932_ (.A(_0486_),
    .B(\sr[197] ),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _0933_ (.A(_0491_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _0934_ (.A(_0486_),
    .B(\sr[198] ),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0492_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_1 _0936_ (.A(_0486_),
    .B(\sr[199] ),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(_0493_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _0938_ (.A(_0486_),
    .B(\sr[200] ),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0494_),
    .X(_0245_));
 sky130_fd_sc_hd__and2_1 _0940_ (.A(_0486_),
    .B(\sr[201] ),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _0941_ (.A(_0495_),
    .X(_0246_));
 sky130_fd_sc_hd__and2_1 _0942_ (.A(_0486_),
    .B(\sr[202] ),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0496_),
    .X(_0247_));
 sky130_fd_sc_hd__buf_2 _0944_ (.A(_0441_),
    .X(_0497_));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(_0497_),
    .B(\sr[203] ),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _0946_ (.A(_0498_),
    .X(_0248_));
 sky130_fd_sc_hd__and2_1 _0947_ (.A(_0497_),
    .B(\sr[204] ),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _0948_ (.A(_0499_),
    .X(_0249_));
 sky130_fd_sc_hd__and2_1 _0949_ (.A(_0497_),
    .B(\sr[205] ),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _0950_ (.A(_0500_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(_0497_),
    .B(\sr[206] ),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _0952_ (.A(_0501_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _0953_ (.A(_0497_),
    .B(\sr[207] ),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _0954_ (.A(_0502_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(_0497_),
    .B(\sr[208] ),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _0956_ (.A(_0503_),
    .X(_0253_));
 sky130_fd_sc_hd__and2_1 _0957_ (.A(_0497_),
    .B(\sr[209] ),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _0958_ (.A(_0504_),
    .X(_0254_));
 sky130_fd_sc_hd__and2_1 _0959_ (.A(_0497_),
    .B(\sr[210] ),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(_0505_),
    .X(_0255_));
 sky130_fd_sc_hd__and2_1 _0961_ (.A(_0497_),
    .B(\sr[211] ),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(_0506_),
    .X(_0000_));
 sky130_fd_sc_hd__and2_1 _0963_ (.A(_0497_),
    .B(\sr[212] ),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0507_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_2 _0965_ (.A(_0441_),
    .X(_0508_));
 sky130_fd_sc_hd__and2_1 _0966_ (.A(_0508_),
    .B(\sr[213] ),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _0967_ (.A(_0509_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _0968_ (.A(_0508_),
    .B(\sr[214] ),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _0969_ (.A(_0510_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _0970_ (.A(_0508_),
    .B(\sr[215] ),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _0971_ (.A(_0511_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(_0508_),
    .B(\sr[216] ),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _0973_ (.A(_0512_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _0974_ (.A(_0508_),
    .B(\sr[217] ),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _0975_ (.A(_0513_),
    .X(_0006_));
 sky130_fd_sc_hd__and2_1 _0976_ (.A(_0508_),
    .B(\sr[218] ),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0514_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _0978_ (.A(_0508_),
    .B(\sr[219] ),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _0979_ (.A(_0515_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _0980_ (.A(_0508_),
    .B(\sr[220] ),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _0981_ (.A(_0516_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _0982_ (.A(_0508_),
    .B(\sr[221] ),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0517_),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _0984_ (.A(_0508_),
    .B(\sr[222] ),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0518_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_2 _0986_ (.A(_0441_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_1 _0987_ (.A(_0519_),
    .B(\sr[223] ),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(_0520_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _0989_ (.A(_0519_),
    .B(\sr[224] ),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(_0521_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _0991_ (.A(_0519_),
    .B(\sr[225] ),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(_0522_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _0993_ (.A(_0519_),
    .B(\sr[226] ),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(_0523_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _0995_ (.A(_0519_),
    .B(\sr[227] ),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(_0524_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(_0519_),
    .B(\sr[228] ),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(_0525_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _0999_ (.A(_0519_),
    .B(\sr[229] ),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(_0526_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _1001_ (.A(_0519_),
    .B(\sr[230] ),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(_0527_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1003_ (.A(_0519_),
    .B(\sr[231] ),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(_0528_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(_0519_),
    .B(\sr[232] ),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(_0529_),
    .X(_0021_));
 sky130_fd_sc_hd__buf_2 _1007_ (.A(_0441_),
    .X(_0530_));
 sky130_fd_sc_hd__and2_1 _1008_ (.A(_0530_),
    .B(\sr[233] ),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(_0531_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _1010_ (.A(_0530_),
    .B(\sr[234] ),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(_0532_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _1012_ (.A(_0530_),
    .B(\sr[235] ),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(_0533_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _1014_ (.A(_0530_),
    .B(\sr[236] ),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(_0534_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _1016_ (.A(_0530_),
    .B(\sr[237] ),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0535_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _1018_ (.A(_0530_),
    .B(\sr[238] ),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(_0536_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _1020_ (.A(_0530_),
    .B(\sr[239] ),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(_0537_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _1022_ (.A(_0530_),
    .B(\sr[240] ),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1023_ (.A(_0538_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _1024_ (.A(_0530_),
    .B(\sr[241] ),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0539_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _1026_ (.A(_0530_),
    .B(\sr[242] ),
    .X(_0256_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1027_ (.A(_0256_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_4 _1028_ (.A(_0441_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _1029_ (.A(_0257_),
    .B(\sr[243] ),
    .X(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(_0258_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _1031_ (.A(_0257_),
    .B(\sr[244] ),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(_0259_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _1033_ (.A(_0257_),
    .B(\sr[245] ),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(_0260_),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _1035_ (.A(_0257_),
    .B(\sr[246] ),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0261_),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _1037_ (.A(_0257_),
    .B(\sr[247] ),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0262_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _1039_ (.A(_0257_),
    .B(\sr[248] ),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0263_),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _1041_ (.A(_0257_),
    .B(\sr[249] ),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _1042_ (.A(_0264_),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _1043_ (.A(_0257_),
    .B(\sr[250] ),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _1044_ (.A(_0265_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _1045_ (.A(_0257_),
    .B(\sr[251] ),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_1 _1046_ (.A(_0266_),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _1047_ (.A(_0257_),
    .B(\sr[252] ),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_1 _1048_ (.A(_0267_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_6 _1049_ (.A(net2),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _1050_ (.A(_0268_),
    .B(\sr[253] ),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0269_),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _1052_ (.A(_0268_),
    .B(\sr[254] ),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0270_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _1054_ (.A(_0268_),
    .B(net3),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0271_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _1056_ (.A(_0268_),
    .B(\sr[0] ),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_1 _1057_ (.A(_0272_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _1058_ (.A(_0268_),
    .B(\sr[1] ),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _1059_ (.A(_0273_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _1060_ (.A(_0268_),
    .B(\sr[2] ),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0274_),
    .X(_0047_));
 sky130_fd_sc_hd__and2_1 _1062_ (.A(_0268_),
    .B(\sr[3] ),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _1063_ (.A(_0275_),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _1064_ (.A(_0268_),
    .B(\sr[4] ),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0276_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _1066_ (.A(_0268_),
    .B(\sr[5] ),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _1067_ (.A(_0277_),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _1068_ (.A(_0268_),
    .B(\sr[6] ),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_1 _1069_ (.A(_0278_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _1070_ (.A(_0284_),
    .B(\sr[7] ),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_1 _1071_ (.A(_0279_),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _1072_ (.A(_0284_),
    .B(\sr[8] ),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _1073_ (.A(_0280_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _1074_ (.A(_0284_),
    .B(\sr[9] ),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(_0281_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _1076_ (.A(_0284_),
    .B(\sr[10] ),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _1077_ (.A(_0282_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _1078_ (.A(_0284_),
    .B(\sr[11] ),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _1079_ (.A(_0283_),
    .X(_0056_));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_9_sclk),
    .D(_0057_),
    .Q(\sr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_9_sclk),
    .D(_0058_),
    .Q(\sr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_leaf_9_sclk),
    .D(_0059_),
    .Q(\sr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_9_sclk),
    .D(_0060_),
    .Q(\sr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_9_sclk),
    .D(_0061_),
    .Q(\sr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_9_sclk),
    .D(_0062_),
    .Q(\sr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_0_sclk),
    .D(_0063_),
    .Q(\sr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_9_sclk),
    .D(_0064_),
    .Q(\sr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_1_sclk),
    .D(_0065_),
    .Q(\sr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_0_sclk),
    .D(_0066_),
    .Q(\sr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_9_sclk),
    .D(_0067_),
    .Q(\sr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_1_sclk),
    .D(_0068_),
    .Q(\sr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_leaf_1_sclk),
    .D(_0069_),
    .Q(\sr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_9_sclk),
    .D(_0070_),
    .Q(\sr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_1_sclk),
    .D(_0071_),
    .Q(\sr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_0_sclk),
    .D(_0072_),
    .Q(\sr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_1_sclk),
    .D(_0073_),
    .Q(\sr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1097_ (.CLK(clknet_leaf_1_sclk),
    .D(_0074_),
    .Q(\sr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_1_sclk),
    .D(_0075_),
    .Q(\sr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_1_sclk),
    .D(_0076_),
    .Q(\sr[32] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_9_sclk),
    .D(_0077_),
    .Q(\sr[33] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_leaf_9_sclk),
    .D(_0078_),
    .Q(\sr[34] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_1_sclk),
    .D(_0079_),
    .Q(\sr[35] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_1_sclk),
    .D(_0080_),
    .Q(\sr[36] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_9_sclk),
    .D(_0081_),
    .Q(\sr[37] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_0_sclk),
    .D(_0082_),
    .Q(\sr[38] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_9_sclk),
    .D(_0083_),
    .Q(\sr[39] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_1_sclk),
    .D(_0084_),
    .Q(\sr[40] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_1_sclk),
    .D(_0085_),
    .Q(\sr[41] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_1_sclk),
    .D(_0086_),
    .Q(\sr[42] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_0_sclk),
    .D(_0087_),
    .Q(\sr[43] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_1_sclk),
    .D(_0088_),
    .Q(\sr[44] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_leaf_0_sclk),
    .D(_0089_),
    .Q(\sr[45] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_0_sclk),
    .D(_0090_),
    .Q(\sr[46] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_2_sclk),
    .D(_0091_),
    .Q(\sr[47] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_0_sclk),
    .D(_0092_),
    .Q(\sr[48] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_leaf_8_sclk),
    .D(_0093_),
    .Q(\sr[49] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_leaf_0_sclk),
    .D(_0094_),
    .Q(\sr[50] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_leaf_0_sclk),
    .D(_0095_),
    .Q(\sr[51] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_leaf_0_sclk),
    .D(_0096_),
    .Q(\sr[52] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_leaf_9_sclk),
    .D(_0097_),
    .Q(\sr[53] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_leaf_0_sclk),
    .D(_0098_),
    .Q(\sr[54] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_leaf_9_sclk),
    .D(_0099_),
    .Q(\sr[55] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_leaf_0_sclk),
    .D(_0100_),
    .Q(\sr[56] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_leaf_9_sclk),
    .D(_0101_),
    .Q(\sr[57] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_leaf_1_sclk),
    .D(_0102_),
    .Q(\sr[58] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_leaf_0_sclk),
    .D(_0103_),
    .Q(\sr[59] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_leaf_1_sclk),
    .D(_0104_),
    .Q(\sr[60] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_leaf_1_sclk),
    .D(_0105_),
    .Q(\sr[61] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_leaf_0_sclk),
    .D(_0106_),
    .Q(\sr[62] ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_leaf_9_sclk),
    .D(_0107_),
    .Q(\sr[63] ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_leaf_2_sclk),
    .D(_0108_),
    .Q(\sr[64] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_leaf_9_sclk),
    .D(_0109_),
    .Q(\sr[65] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_leaf_2_sclk),
    .D(_0110_),
    .Q(\sr[66] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_leaf_1_sclk),
    .D(_0111_),
    .Q(\sr[67] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_leaf_0_sclk),
    .D(_0112_),
    .Q(\sr[68] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_leaf_9_sclk),
    .D(_0113_),
    .Q(\sr[69] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_leaf_0_sclk),
    .D(_0114_),
    .Q(\sr[70] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_leaf_9_sclk),
    .D(_0115_),
    .Q(\sr[71] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_leaf_8_sclk),
    .D(_0116_),
    .Q(\sr[72] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_leaf_0_sclk),
    .D(_0117_),
    .Q(\sr[73] ));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(clknet_leaf_1_sclk),
    .D(_0118_),
    .Q(\sr[74] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_leaf_2_sclk),
    .D(_0119_),
    .Q(\sr[75] ));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_leaf_0_sclk),
    .D(_0120_),
    .Q(\sr[76] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_leaf_0_sclk),
    .D(_0121_),
    .Q(\sr[77] ));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_leaf_9_sclk),
    .D(_0122_),
    .Q(\sr[78] ));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_leaf_8_sclk),
    .D(_0123_),
    .Q(\sr[79] ));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_leaf_8_sclk),
    .D(_0124_),
    .Q(\sr[80] ));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_leaf_8_sclk),
    .D(_0125_),
    .Q(\sr[81] ));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_leaf_2_sclk),
    .D(_0126_),
    .Q(\sr[82] ));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_leaf_2_sclk),
    .D(_0127_),
    .Q(\sr[83] ));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_leaf_10_sclk),
    .D(_0128_),
    .Q(\sr[84] ));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_leaf_2_sclk),
    .D(_0129_),
    .Q(\sr[85] ));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_leaf_2_sclk),
    .D(_0130_),
    .Q(\sr[86] ));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_leaf_0_sclk),
    .D(_0131_),
    .Q(\sr[87] ));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_leaf_0_sclk),
    .D(_0132_),
    .Q(\sr[88] ));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_leaf_2_sclk),
    .D(_0133_),
    .Q(\sr[89] ));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_leaf_2_sclk),
    .D(_0134_),
    .Q(\sr[90] ));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(clknet_leaf_2_sclk),
    .D(_0135_),
    .Q(\sr[91] ));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_leaf_10_sclk),
    .D(_0136_),
    .Q(\sr[92] ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_leaf_2_sclk),
    .D(_0137_),
    .Q(\sr[93] ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_leaf_8_sclk),
    .D(_0138_),
    .Q(\sr[94] ));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_leaf_8_sclk),
    .D(_0139_),
    .Q(\sr[95] ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_leaf_10_sclk),
    .D(_0140_),
    .Q(\sr[96] ));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_leaf_2_sclk),
    .D(_0141_),
    .Q(\sr[97] ));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_leaf_8_sclk),
    .D(_0142_),
    .Q(\sr[98] ));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_leaf_2_sclk),
    .D(_0143_),
    .Q(\sr[99] ));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_leaf_10_sclk),
    .D(_0144_),
    .Q(\sr[100] ));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_leaf_3_sclk),
    .D(_0145_),
    .Q(\sr[101] ));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_leaf_8_sclk),
    .D(_0146_),
    .Q(\sr[102] ));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_leaf_8_sclk),
    .D(_0147_),
    .Q(\sr[103] ));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_leaf_3_sclk),
    .D(_0148_),
    .Q(\sr[104] ));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_leaf_10_sclk),
    .D(_0149_),
    .Q(\sr[105] ));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_leaf_10_sclk),
    .D(_0150_),
    .Q(\sr[106] ));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_leaf_2_sclk),
    .D(_0151_),
    .Q(\sr[107] ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_leaf_5_sclk),
    .D(_0152_),
    .Q(\sr[108] ));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_leaf_8_sclk),
    .D(_0153_),
    .Q(\sr[109] ));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_leaf_8_sclk),
    .D(_0154_),
    .Q(\sr[110] ));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_leaf_2_sclk),
    .D(_0155_),
    .Q(\sr[111] ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_leaf_8_sclk),
    .D(_0156_),
    .Q(\sr[112] ));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_leaf_2_sclk),
    .D(_0157_),
    .Q(\sr[113] ));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_leaf_2_sclk),
    .D(_0158_),
    .Q(\sr[114] ));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_leaf_7_sclk),
    .D(_0159_),
    .Q(\sr[115] ));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_leaf_8_sclk),
    .D(_0160_),
    .Q(\sr[116] ));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_leaf_3_sclk),
    .D(_0161_),
    .Q(\sr[117] ));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_leaf_8_sclk),
    .D(_0162_),
    .Q(\sr[118] ));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(clknet_leaf_5_sclk),
    .D(_0163_),
    .Q(\sr[119] ));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_leaf_5_sclk),
    .D(_0164_),
    .Q(\sr[120] ));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(clknet_leaf_5_sclk),
    .D(_0165_),
    .Q(\sr[121] ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_leaf_8_sclk),
    .D(_0166_),
    .Q(\sr[122] ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_leaf_2_sclk),
    .D(_0167_),
    .Q(\sr[123] ));
 sky130_fd_sc_hd__dfxtp_2 _1191_ (.CLK(clknet_leaf_8_sclk),
    .D(_0168_),
    .Q(\sr[124] ));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_leaf_3_sclk),
    .D(_0169_),
    .Q(\sr[125] ));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_leaf_5_sclk),
    .D(_0170_),
    .Q(\sr[126] ));
 sky130_fd_sc_hd__dfxtp_2 _1194_ (.CLK(clknet_leaf_3_sclk),
    .D(_0171_),
    .Q(\sr[127] ));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_leaf_2_sclk),
    .D(_0172_),
    .Q(\sr[128] ));
 sky130_fd_sc_hd__dfxtp_2 _1196_ (.CLK(clknet_leaf_2_sclk),
    .D(_0173_),
    .Q(\sr[129] ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_leaf_3_sclk),
    .D(_0174_),
    .Q(\sr[130] ));
 sky130_fd_sc_hd__dfxtp_2 _1198_ (.CLK(clknet_leaf_4_sclk),
    .D(_0175_),
    .Q(\sr[131] ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(clknet_leaf_8_sclk),
    .D(_0176_),
    .Q(\sr[132] ));
 sky130_fd_sc_hd__dfxtp_2 _1200_ (.CLK(clknet_leaf_5_sclk),
    .D(_0177_),
    .Q(\sr[133] ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_leaf_3_sclk),
    .D(_0178_),
    .Q(\sr[134] ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_leaf_3_sclk),
    .D(_0179_),
    .Q(\sr[135] ));
 sky130_fd_sc_hd__dfxtp_2 _1203_ (.CLK(clknet_leaf_7_sclk),
    .D(_0180_),
    .Q(\sr[136] ));
 sky130_fd_sc_hd__dfxtp_2 _1204_ (.CLK(clknet_leaf_5_sclk),
    .D(_0181_),
    .Q(\sr[137] ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_leaf_8_sclk),
    .D(_0182_),
    .Q(\sr[138] ));
 sky130_fd_sc_hd__dfxtp_2 _1206_ (.CLK(clknet_leaf_3_sclk),
    .D(_0183_),
    .Q(\sr[139] ));
 sky130_fd_sc_hd__dfxtp_2 _1207_ (.CLK(clknet_leaf_3_sclk),
    .D(_0184_),
    .Q(\sr[140] ));
 sky130_fd_sc_hd__dfxtp_4 _1208_ (.CLK(clknet_leaf_8_sclk),
    .D(_0185_),
    .Q(\sr[141] ));
 sky130_fd_sc_hd__dfxtp_2 _1209_ (.CLK(clknet_leaf_3_sclk),
    .D(_0186_),
    .Q(\sr[142] ));
 sky130_fd_sc_hd__dfxtp_2 _1210_ (.CLK(clknet_leaf_3_sclk),
    .D(_0187_),
    .Q(\sr[143] ));
 sky130_fd_sc_hd__dfxtp_2 _1211_ (.CLK(clknet_leaf_8_sclk),
    .D(_0188_),
    .Q(\sr[144] ));
 sky130_fd_sc_hd__dfxtp_2 _1212_ (.CLK(clknet_leaf_3_sclk),
    .D(_0189_),
    .Q(\sr[145] ));
 sky130_fd_sc_hd__dfxtp_2 _1213_ (.CLK(clknet_leaf_2_sclk),
    .D(_0190_),
    .Q(\sr[146] ));
 sky130_fd_sc_hd__dfxtp_2 _1214_ (.CLK(clknet_leaf_2_sclk),
    .D(_0191_),
    .Q(\sr[147] ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_leaf_3_sclk),
    .D(_0192_),
    .Q(\sr[148] ));
 sky130_fd_sc_hd__dfxtp_2 _1216_ (.CLK(clknet_leaf_3_sclk),
    .D(_0193_),
    .Q(\sr[149] ));
 sky130_fd_sc_hd__dfxtp_2 _1217_ (.CLK(clknet_leaf_2_sclk),
    .D(_0194_),
    .Q(\sr[150] ));
 sky130_fd_sc_hd__dfxtp_2 _1218_ (.CLK(clknet_leaf_8_sclk),
    .D(_0195_),
    .Q(\sr[151] ));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_leaf_8_sclk),
    .D(_0196_),
    .Q(\sr[152] ));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_leaf_5_sclk),
    .D(_0197_),
    .Q(\sr[153] ));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_leaf_6_sclk),
    .D(_0198_),
    .Q(\sr[154] ));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_leaf_7_sclk),
    .D(_0199_),
    .Q(\sr[155] ));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_leaf_4_sclk),
    .D(_0200_),
    .Q(\sr[156] ));
 sky130_fd_sc_hd__dfxtp_2 _1224_ (.CLK(clknet_leaf_7_sclk),
    .D(_0201_),
    .Q(\sr[157] ));
 sky130_fd_sc_hd__dfxtp_2 _1225_ (.CLK(clknet_leaf_3_sclk),
    .D(_0202_),
    .Q(\sr[158] ));
 sky130_fd_sc_hd__dfxtp_2 _1226_ (.CLK(clknet_leaf_6_sclk),
    .D(_0203_),
    .Q(\sr[159] ));
 sky130_fd_sc_hd__dfxtp_2 _1227_ (.CLK(clknet_leaf_4_sclk),
    .D(_0204_),
    .Q(\sr[160] ));
 sky130_fd_sc_hd__dfxtp_2 _1228_ (.CLK(clknet_leaf_5_sclk),
    .D(_0205_),
    .Q(\sr[161] ));
 sky130_fd_sc_hd__dfxtp_2 _1229_ (.CLK(clknet_leaf_7_sclk),
    .D(_0206_),
    .Q(\sr[162] ));
 sky130_fd_sc_hd__dfxtp_2 _1230_ (.CLK(clknet_leaf_4_sclk),
    .D(_0207_),
    .Q(\sr[163] ));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_leaf_7_sclk),
    .D(_0208_),
    .Q(\sr[164] ));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_leaf_5_sclk),
    .D(_0209_),
    .Q(\sr[165] ));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_leaf_4_sclk),
    .D(_0210_),
    .Q(\sr[166] ));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_leaf_4_sclk),
    .D(_0211_),
    .Q(\sr[167] ));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_leaf_6_sclk),
    .D(_0212_),
    .Q(\sr[168] ));
 sky130_fd_sc_hd__dfxtp_2 _1236_ (.CLK(clknet_leaf_5_sclk),
    .D(_0213_),
    .Q(\sr[169] ));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_leaf_6_sclk),
    .D(_0214_),
    .Q(\sr[170] ));
 sky130_fd_sc_hd__dfxtp_2 _1238_ (.CLK(clknet_leaf_7_sclk),
    .D(_0215_),
    .Q(\sr[171] ));
 sky130_fd_sc_hd__dfxtp_2 _1239_ (.CLK(clknet_leaf_7_sclk),
    .D(_0216_),
    .Q(\sr[172] ));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_leaf_7_sclk),
    .D(_0217_),
    .Q(\sr[173] ));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_leaf_6_sclk),
    .D(_0218_),
    .Q(\sr[174] ));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_leaf_5_sclk),
    .D(_0219_),
    .Q(\sr[175] ));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_leaf_5_sclk),
    .D(_0220_),
    .Q(\sr[176] ));
 sky130_fd_sc_hd__dfxtp_2 _1244_ (.CLK(clknet_leaf_5_sclk),
    .D(_0221_),
    .Q(\sr[177] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_leaf_3_sclk),
    .D(_0222_),
    .Q(\sr[178] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_leaf_4_sclk),
    .D(_0223_),
    .Q(\sr[179] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_leaf_6_sclk),
    .D(_0224_),
    .Q(\sr[180] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_leaf_4_sclk),
    .D(_0225_),
    .Q(\sr[181] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_leaf_5_sclk),
    .D(_0226_),
    .Q(\sr[182] ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_leaf_7_sclk),
    .D(_0227_),
    .Q(\sr[183] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_leaf_6_sclk),
    .D(_0228_),
    .Q(\sr[184] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_leaf_7_sclk),
    .D(_0229_),
    .Q(\sr[185] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_leaf_5_sclk),
    .D(_0230_),
    .Q(\sr[186] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_leaf_7_sclk),
    .D(_0231_),
    .Q(\sr[187] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_leaf_7_sclk),
    .D(_0232_),
    .Q(\sr[188] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_leaf_6_sclk),
    .D(_0233_),
    .Q(\sr[189] ));
 sky130_fd_sc_hd__dfxtp_2 _1257_ (.CLK(clknet_leaf_4_sclk),
    .D(_0234_),
    .Q(\sr[190] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_leaf_6_sclk),
    .D(_0235_),
    .Q(\sr[191] ));
 sky130_fd_sc_hd__dfxtp_2 _1259_ (.CLK(clknet_leaf_7_sclk),
    .D(_0236_),
    .Q(\sr[192] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_leaf_3_sclk),
    .D(_0237_),
    .Q(\sr[193] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_leaf_6_sclk),
    .D(_0238_),
    .Q(\sr[194] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_leaf_7_sclk),
    .D(_0239_),
    .Q(\sr[195] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_leaf_4_sclk),
    .D(_0240_),
    .Q(\sr[196] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_leaf_7_sclk),
    .D(_0241_),
    .Q(\sr[197] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_leaf_4_sclk),
    .D(_0242_),
    .Q(\sr[198] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_leaf_4_sclk),
    .D(_0243_),
    .Q(\sr[199] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_leaf_6_sclk),
    .D(_0244_),
    .Q(\sr[200] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_leaf_4_sclk),
    .D(_0245_),
    .Q(\sr[201] ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_leaf_4_sclk),
    .D(_0246_),
    .Q(\sr[202] ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_leaf_4_sclk),
    .D(_0247_),
    .Q(\sr[203] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_leaf_4_sclk),
    .D(_0248_),
    .Q(\sr[204] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_leaf_3_sclk),
    .D(_0249_),
    .Q(\sr[205] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_leaf_3_sclk),
    .D(_0250_),
    .Q(\sr[206] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_leaf_5_sclk),
    .D(_0251_),
    .Q(\sr[207] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_leaf_6_sclk),
    .D(_0252_),
    .Q(\sr[208] ));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_leaf_6_sclk),
    .D(_0253_),
    .Q(\sr[209] ));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_leaf_6_sclk),
    .D(_0254_),
    .Q(\sr[210] ));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_leaf_6_sclk),
    .D(_0255_),
    .Q(\sr[211] ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_leaf_4_sclk),
    .D(_0000_),
    .Q(\sr[212] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_leaf_5_sclk),
    .D(_0001_),
    .Q(\sr[213] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_leaf_7_sclk),
    .D(_0002_),
    .Q(\sr[214] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_leaf_4_sclk),
    .D(_0003_),
    .Q(\sr[215] ));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_leaf_7_sclk),
    .D(_0004_),
    .Q(\sr[216] ));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_leaf_6_sclk),
    .D(_0005_),
    .Q(\sr[217] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_leaf_5_sclk),
    .D(_0006_),
    .Q(\sr[218] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_leaf_6_sclk),
    .D(_0007_),
    .Q(\sr[219] ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_leaf_5_sclk),
    .D(_0008_),
    .Q(\sr[220] ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_leaf_6_sclk),
    .D(_0009_),
    .Q(\sr[221] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_leaf_6_sclk),
    .D(_0010_),
    .Q(\sr[222] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_leaf_6_sclk),
    .D(_0011_),
    .Q(\sr[223] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_leaf_6_sclk),
    .D(_0012_),
    .Q(\sr[224] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_leaf_4_sclk),
    .D(_0013_),
    .Q(\sr[225] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_leaf_3_sclk),
    .D(_0014_),
    .Q(\sr[226] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_leaf_7_sclk),
    .D(_0015_),
    .Q(\sr[227] ));
 sky130_fd_sc_hd__dfxtp_2 _1295_ (.CLK(clknet_leaf_6_sclk),
    .D(_0016_),
    .Q(\sr[228] ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_leaf_4_sclk),
    .D(_0017_),
    .Q(\sr[229] ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_leaf_4_sclk),
    .D(_0018_),
    .Q(\sr[230] ));
 sky130_fd_sc_hd__dfxtp_2 _1298_ (.CLK(clknet_leaf_4_sclk),
    .D(_0019_),
    .Q(\sr[231] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_leaf_3_sclk),
    .D(_0020_),
    .Q(\sr[232] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_leaf_4_sclk),
    .D(_0021_),
    .Q(\sr[233] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_leaf_7_sclk),
    .D(_0022_),
    .Q(\sr[234] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_leaf_4_sclk),
    .D(_0023_),
    .Q(\sr[235] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_leaf_6_sclk),
    .D(_0024_),
    .Q(\sr[236] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_leaf_7_sclk),
    .D(_0025_),
    .Q(\sr[237] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_leaf_5_sclk),
    .D(_0026_),
    .Q(\sr[238] ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_leaf_6_sclk),
    .D(_0027_),
    .Q(\sr[239] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_leaf_6_sclk),
    .D(_0028_),
    .Q(\sr[240] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_leaf_4_sclk),
    .D(_0029_),
    .Q(\sr[241] ));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_leaf_7_sclk),
    .D(_0030_),
    .Q(\sr[242] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_leaf_7_sclk),
    .D(_0031_),
    .Q(\sr[243] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_leaf_3_sclk),
    .D(_0032_),
    .Q(\sr[244] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_leaf_7_sclk),
    .D(_0033_),
    .Q(\sr[245] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_leaf_5_sclk),
    .D(_0034_),
    .Q(\sr[246] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_leaf_5_sclk),
    .D(_0035_),
    .Q(\sr[247] ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_leaf_3_sclk),
    .D(_0036_),
    .Q(\sr[248] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_leaf_2_sclk),
    .D(_0037_),
    .Q(\sr[249] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_leaf_5_sclk),
    .D(_0038_),
    .Q(\sr[250] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_leaf_7_sclk),
    .D(_0039_),
    .Q(\sr[251] ));
 sky130_fd_sc_hd__dfxtp_2 _1319_ (.CLK(clknet_leaf_8_sclk),
    .D(_0040_),
    .Q(\sr[252] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_leaf_3_sclk),
    .D(_0041_),
    .Q(\sr[253] ));
 sky130_fd_sc_hd__dfxtp_2 _1321_ (.CLK(clknet_leaf_8_sclk),
    .D(_0042_),
    .Q(\sr[254] ));
 sky130_fd_sc_hd__dfxtp_2 _1322_ (.CLK(clknet_leaf_5_sclk),
    .D(_0043_),
    .Q(net260));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(net262),
    .D(\sr[0] ),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(net261),
    .D(\sr[1] ),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(net263),
    .D(\sr[2] ),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(net261),
    .D(\sr[3] ),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_1 _1327_ (.CLK(net261),
    .D(\sr[4] ),
    .Q(net204));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(net261),
    .D(\sr[5] ),
    .Q(net215));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(net261),
    .D(\sr[6] ),
    .Q(net226));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(net265),
    .D(\sr[7] ),
    .Q(net237));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(net265),
    .D(\sr[8] ),
    .Q(net248));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(net263),
    .D(\sr[9] ),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_1 _1333_ (.CLK(net265),
    .D(\sr[10] ),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1334_ (.CLK(net264),
    .D(\sr[11] ),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1335_ (.CLK(net263),
    .D(\sr[12] ),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1336_ (.CLK(net263),
    .D(\sr[13] ),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _1337_ (.CLK(net264),
    .D(\sr[14] ),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _1338_ (.CLK(net262),
    .D(\sr[15] ),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _1339_ (.CLK(net263),
    .D(\sr[16] ),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _1340_ (.CLK(net261),
    .D(\sr[17] ),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _1341_ (.CLK(net262),
    .D(\sr[18] ),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _1342_ (.CLK(net264),
    .D(\sr[19] ),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _1343_ (.CLK(net262),
    .D(\sr[20] ),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _1344_ (.CLK(net265),
    .D(\sr[21] ),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _1345_ (.CLK(net266),
    .D(\sr[22] ),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _1346_ (.CLK(net263),
    .D(\sr[23] ),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _1347_ (.CLK(net264),
    .D(\sr[24] ),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_1 _1348_ (.CLK(net265),
    .D(\sr[25] ),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_1 _1349_ (.CLK(net262),
    .D(\sr[26] ),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_1 _1350_ (.CLK(net262),
    .D(\sr[27] ),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _1351_ (.CLK(net261),
    .D(\sr[28] ),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_1 _1352_ (.CLK(net265),
    .D(\sr[29] ),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_1 _1353_ (.CLK(net271),
    .D(\sr[30] ),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_1 _1354_ (.CLK(net264),
    .D(\sr[31] ),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _1355_ (.CLK(net271),
    .D(\sr[32] ),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 _1356_ (.CLK(net266),
    .D(\sr[33] ),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_1 _1357_ (.CLK(net266),
    .D(\sr[34] ),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _1358_ (.CLK(net261),
    .D(\sr[35] ),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_1 _1359_ (.CLK(net261),
    .D(\sr[36] ),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_1 _1360_ (.CLK(net268),
    .D(\sr[37] ),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_1 _1361_ (.CLK(net261),
    .D(\sr[38] ),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_1 _1362_ (.CLK(net262),
    .D(\sr[39] ),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_1 _1363_ (.CLK(net268),
    .D(\sr[40] ),
    .Q(net194));
 sky130_fd_sc_hd__dfxtp_1 _1364_ (.CLK(net262),
    .D(\sr[41] ),
    .Q(net195));
 sky130_fd_sc_hd__dfxtp_1 _1365_ (.CLK(net265),
    .D(\sr[42] ),
    .Q(net196));
 sky130_fd_sc_hd__dfxtp_1 _1366_ (.CLK(net271),
    .D(\sr[43] ),
    .Q(net197));
 sky130_fd_sc_hd__dfxtp_1 _1367_ (.CLK(net269),
    .D(\sr[44] ),
    .Q(net198));
 sky130_fd_sc_hd__dfxtp_1 _1368_ (.CLK(net264),
    .D(\sr[45] ),
    .Q(net199));
 sky130_fd_sc_hd__dfxtp_1 _1369_ (.CLK(net266),
    .D(\sr[46] ),
    .Q(net200));
 sky130_fd_sc_hd__dfxtp_1 _1370_ (.CLK(net269),
    .D(\sr[47] ),
    .Q(net201));
 sky130_fd_sc_hd__dfxtp_1 _1371_ (.CLK(net264),
    .D(\sr[48] ),
    .Q(net202));
 sky130_fd_sc_hd__dfxtp_1 _1372_ (.CLK(net262),
    .D(\sr[49] ),
    .Q(net203));
 sky130_fd_sc_hd__dfxtp_1 _1373_ (.CLK(net266),
    .D(\sr[50] ),
    .Q(net205));
 sky130_fd_sc_hd__dfxtp_1 _1374_ (.CLK(net264),
    .D(\sr[51] ),
    .Q(net206));
 sky130_fd_sc_hd__dfxtp_1 _1375_ (.CLK(net264),
    .D(\sr[52] ),
    .Q(net207));
 sky130_fd_sc_hd__dfxtp_1 _1376_ (.CLK(net266),
    .D(\sr[53] ),
    .Q(net208));
 sky130_fd_sc_hd__dfxtp_1 _1377_ (.CLK(net266),
    .D(\sr[54] ),
    .Q(net209));
 sky130_fd_sc_hd__dfxtp_1 _1378_ (.CLK(net272),
    .D(\sr[55] ),
    .Q(net210));
 sky130_fd_sc_hd__dfxtp_1 _1379_ (.CLK(net266),
    .D(\sr[56] ),
    .Q(net211));
 sky130_fd_sc_hd__dfxtp_1 _1380_ (.CLK(net266),
    .D(\sr[57] ),
    .Q(net212));
 sky130_fd_sc_hd__dfxtp_1 _1381_ (.CLK(net262),
    .D(\sr[58] ),
    .Q(net213));
 sky130_fd_sc_hd__dfxtp_1 _1382_ (.CLK(net266),
    .D(\sr[59] ),
    .Q(net214));
 sky130_fd_sc_hd__dfxtp_1 _1383_ (.CLK(net265),
    .D(\sr[60] ),
    .Q(net216));
 sky130_fd_sc_hd__dfxtp_1 _1384_ (.CLK(net267),
    .D(\sr[61] ),
    .Q(net217));
 sky130_fd_sc_hd__dfxtp_1 _1385_ (.CLK(net271),
    .D(\sr[62] ),
    .Q(net218));
 sky130_fd_sc_hd__dfxtp_1 _1386_ (.CLK(net267),
    .D(\sr[63] ),
    .Q(net219));
 sky130_fd_sc_hd__dfxtp_1 _1387_ (.CLK(net269),
    .D(\sr[64] ),
    .Q(net220));
 sky130_fd_sc_hd__dfxtp_1 _1388_ (.CLK(net267),
    .D(\sr[65] ),
    .Q(net221));
 sky130_fd_sc_hd__dfxtp_1 _1389_ (.CLK(net267),
    .D(\sr[66] ),
    .Q(net222));
 sky130_fd_sc_hd__dfxtp_1 _1390_ (.CLK(net272),
    .D(\sr[67] ),
    .Q(net223));
 sky130_fd_sc_hd__dfxtp_1 _1391_ (.CLK(net263),
    .D(\sr[68] ),
    .Q(net224));
 sky130_fd_sc_hd__dfxtp_1 _1392_ (.CLK(net264),
    .D(\sr[69] ),
    .Q(net225));
 sky130_fd_sc_hd__dfxtp_1 _1393_ (.CLK(net271),
    .D(\sr[70] ),
    .Q(net227));
 sky130_fd_sc_hd__dfxtp_1 _1394_ (.CLK(net277),
    .D(\sr[71] ),
    .Q(net228));
 sky130_fd_sc_hd__dfxtp_1 _1395_ (.CLK(net272),
    .D(\sr[72] ),
    .Q(net229));
 sky130_fd_sc_hd__dfxtp_1 _1396_ (.CLK(net269),
    .D(\sr[73] ),
    .Q(net230));
 sky130_fd_sc_hd__dfxtp_1 _1397_ (.CLK(net274),
    .D(\sr[74] ),
    .Q(net231));
 sky130_fd_sc_hd__dfxtp_1 _1398_ (.CLK(net267),
    .D(\sr[75] ),
    .Q(net232));
 sky130_fd_sc_hd__dfxtp_1 _1399_ (.CLK(net267),
    .D(\sr[76] ),
    .Q(net233));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(net269),
    .D(\sr[77] ),
    .Q(net234));
 sky130_fd_sc_hd__dfxtp_1 _1401_ (.CLK(net271),
    .D(\sr[78] ),
    .Q(net235));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(net275),
    .D(\sr[79] ),
    .Q(net236));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(net274),
    .D(\sr[80] ),
    .Q(net238));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(net274),
    .D(\sr[81] ),
    .Q(net239));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(net269),
    .D(\sr[82] ),
    .Q(net240));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(net269),
    .D(\sr[83] ),
    .Q(net241));
 sky130_fd_sc_hd__dfxtp_1 _1407_ (.CLK(net271),
    .D(\sr[84] ),
    .Q(net242));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(net267),
    .D(\sr[85] ),
    .Q(net243));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(net270),
    .D(\sr[86] ),
    .Q(net244));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(net272),
    .D(\sr[87] ),
    .Q(net245));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(net270),
    .D(\sr[88] ),
    .Q(net246));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(net269),
    .D(\sr[89] ),
    .Q(net247));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(net270),
    .D(\sr[90] ),
    .Q(net249));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(net269),
    .D(\sr[91] ),
    .Q(net250));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(net269),
    .D(\sr[92] ),
    .Q(net251));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(net270),
    .D(\sr[93] ),
    .Q(net252));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(net270),
    .D(\sr[94] ),
    .Q(net253));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(net273),
    .D(\sr[95] ),
    .Q(net254));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(net270),
    .D(\sr[96] ),
    .Q(net255));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(net272),
    .D(\sr[97] ),
    .Q(net256));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(net272),
    .D(\sr[98] ),
    .Q(net257));
 sky130_fd_sc_hd__dfxtp_1 _1422_ (.CLK(net273),
    .D(\sr[99] ),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_1 _1423_ (.CLK(net273),
    .D(\sr[100] ),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_1 _1424_ (.CLK(net277),
    .D(\sr[101] ),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _1425_ (.CLK(net275),
    .D(\sr[102] ),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _1426_ (.CLK(net272),
    .D(\sr[103] ),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _1427_ (.CLK(net275),
    .D(\sr[104] ),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(net274),
    .D(\sr[105] ),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(net274),
    .D(\sr[106] ),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(net279),
    .D(\sr[107] ),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(net278),
    .D(\sr[108] ),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(net274),
    .D(\sr[109] ),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(net275),
    .D(\sr[110] ),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1434_ (.CLK(net278),
    .D(\sr[111] ),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1435_ (.CLK(net278),
    .D(\sr[112] ),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(net279),
    .D(\sr[113] ),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(net275),
    .D(\sr[114] ),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(net275),
    .D(\sr[115] ),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(net278),
    .D(\sr[116] ),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(net275),
    .D(\sr[117] ),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(net279),
    .D(\sr[118] ),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(net275),
    .D(\sr[119] ),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(net274),
    .D(\sr[120] ),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(net280),
    .D(\sr[121] ),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(net278),
    .D(\sr[122] ),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(net279),
    .D(\sr[123] ),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(net274),
    .D(\sr[124] ),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(net275),
    .D(\sr[125] ),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(net280),
    .D(\sr[126] ),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(net274),
    .D(\sr[127] ),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(net276),
    .D(\sr[128] ),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(net274),
    .D(\sr[129] ),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(net276),
    .D(\sr[130] ),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(net270),
    .D(\sr[131] ),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(net279),
    .D(\sr[132] ),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1456_ (.CLK(net276),
    .D(\sr[133] ),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(net278),
    .D(\sr[134] ),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(net278),
    .D(\sr[135] ),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(net279),
    .D(\sr[136] ),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(net272),
    .D(\sr[137] ),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(net279),
    .D(\sr[138] ),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(net276),
    .D(\sr[139] ),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(net276),
    .D(\sr[140] ),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(net272),
    .D(\sr[141] ),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(net278),
    .D(\sr[142] ),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(net273),
    .D(\sr[143] ),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(net276),
    .D(\sr[144] ),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(net279),
    .D(\sr[145] ),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(net273),
    .D(\sr[146] ),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(net273),
    .D(\sr[147] ),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(net282),
    .D(\sr[148] ),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _1472_ (.CLK(net276),
    .D(\sr[149] ),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _1473_ (.CLK(net272),
    .D(\sr[150] ),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _1474_ (.CLK(net273),
    .D(\sr[151] ),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _1475_ (.CLK(net280),
    .D(\sr[152] ),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_2 _1476_ (.CLK(net287),
    .D(\sr[153] ),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_2 _1477_ (.CLK(net289),
    .D(\sr[154] ),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_2 _1478_ (.CLK(net288),
    .D(\sr[155] ),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _1479_ (.CLK(net287),
    .D(\sr[156] ),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _1480_ (.CLK(net282),
    .D(\sr[157] ),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _1481_ (.CLK(net280),
    .D(\sr[158] ),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _1482_ (.CLK(net278),
    .D(\sr[159] ),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _1483_ (.CLK(net276),
    .D(\sr[160] ),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _1484_ (.CLK(net278),
    .D(\sr[161] ),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _1485_ (.CLK(net283),
    .D(\sr[162] ),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _1486_ (.CLK(net280),
    .D(\sr[163] ),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _1487_ (.CLK(net284),
    .D(\sr[164] ),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _1488_ (.CLK(net289),
    .D(\sr[165] ),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _1489_ (.CLK(net281),
    .D(\sr[166] ),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _1490_ (.CLK(net284),
    .D(\sr[167] ),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _1491_ (.CLK(net284),
    .D(\sr[168] ),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _1492_ (.CLK(net280),
    .D(\sr[169] ),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _1493_ (.CLK(net283),
    .D(\sr[170] ),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _1494_ (.CLK(net275),
    .D(\sr[171] ),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _1495_ (.CLK(net279),
    .D(\sr[172] ),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _1496_ (.CLK(net282),
    .D(\sr[173] ),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _1497_ (.CLK(net283),
    .D(\sr[174] ),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _1498_ (.CLK(net282),
    .D(\sr[175] ),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _1499_ (.CLK(net281),
    .D(\sr[176] ),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _1500_ (.CLK(net281),
    .D(\sr[177] ),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_2 _1501_ (.CLK(net290),
    .D(\sr[178] ),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _1502_ (.CLK(net290),
    .D(\sr[179] ),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _1503_ (.CLK(net285),
    .D(\sr[180] ),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _1504_ (.CLK(net288),
    .D(\sr[181] ),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _1505_ (.CLK(net288),
    .D(\sr[182] ),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _1506_ (.CLK(net289),
    .D(\sr[183] ),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _1507_ (.CLK(net282),
    .D(\sr[184] ),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _1508_ (.CLK(net284),
    .D(\sr[185] ),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _1509_ (.CLK(net281),
    .D(\sr[186] ),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _1510_ (.CLK(net281),
    .D(\sr[187] ),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _1511_ (.CLK(net285),
    .D(\sr[188] ),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _1512_ (.CLK(net281),
    .D(\sr[189] ),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _1513_ (.CLK(net282),
    .D(\sr[190] ),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _1514_ (.CLK(net289),
    .D(\sr[191] ),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _1515_ (.CLK(net282),
    .D(\sr[192] ),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _1516_ (.CLK(net289),
    .D(\sr[193] ),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _1517_ (.CLK(net290),
    .D(\sr[194] ),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _1518_ (.CLK(net288),
    .D(\sr[195] ),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _1519_ (.CLK(net290),
    .D(\sr[196] ),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _1520_ (.CLK(net288),
    .D(\sr[197] ),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _1521_ (.CLK(net289),
    .D(\sr[198] ),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_1 _1522_ (.CLK(net285),
    .D(\sr[199] ),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_1 _1523_ (.CLK(net285),
    .D(\sr[200] ),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _1524_ (.CLK(net285),
    .D(\sr[201] ),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _1525_ (.CLK(net287),
    .D(\sr[202] ),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _1526_ (.CLK(net288),
    .D(\sr[203] ),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _1527_ (.CLK(net288),
    .D(\sr[204] ),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _1528_ (.CLK(net290),
    .D(\sr[205] ),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _1529_ (.CLK(net289),
    .D(\sr[206] ),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _1530_ (.CLK(net289),
    .D(\sr[207] ),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _1531_ (.CLK(net287),
    .D(\sr[208] ),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _1532_ (.CLK(net283),
    .D(\sr[209] ),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(net288),
    .D(\sr[210] ),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _1534_ (.CLK(net287),
    .D(\sr[211] ),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _1535_ (.CLK(net287),
    .D(\sr[212] ),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _1536_ (.CLK(net284),
    .D(\sr[213] ),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _1537_ (.CLK(net290),
    .D(\sr[214] ),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(net287),
    .D(\sr[215] ),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(net287),
    .D(\sr[216] ),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _1540_ (.CLK(net289),
    .D(\sr[217] ),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _1541_ (.CLK(net291),
    .D(\sr[218] ),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(net285),
    .D(\sr[219] ),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _1543_ (.CLK(net285),
    .D(\sr[220] ),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(net284),
    .D(\sr[221] ),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(net283),
    .D(\sr[222] ),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _1546_ (.CLK(net283),
    .D(\sr[223] ),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _1547_ (.CLK(net283),
    .D(\sr[224] ),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(net281),
    .D(\sr[225] ),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _1549_ (.CLK(net281),
    .D(\sr[226] ),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _1550_ (.CLK(net283),
    .D(\sr[227] ),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _1551_ (.CLK(net282),
    .D(\sr[228] ),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _1552_ (.CLK(net284),
    .D(\sr[229] ),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(net283),
    .D(\sr[230] ),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _1554_ (.CLK(net281),
    .D(\sr[231] ),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _1555_ (.CLK(net285),
    .D(\sr[232] ),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _1556_ (.CLK(net281),
    .D(\sr[233] ),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _1557_ (.CLK(net287),
    .D(\sr[234] ),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(net284),
    .D(\sr[235] ),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(net288),
    .D(\sr[236] ),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(net283),
    .D(\sr[237] ),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(net285),
    .D(\sr[238] ),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(net292),
    .D(\sr[239] ),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(net286),
    .D(\sr[240] ),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(net289),
    .D(\sr[241] ),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _1565_ (.CLK(net290),
    .D(\sr[242] ),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(net286),
    .D(\sr[243] ),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(net285),
    .D(\sr[244] ),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _1568_ (.CLK(net282),
    .D(\sr[245] ),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _1569_ (.CLK(net284),
    .D(\sr[246] ),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _1570_ (.CLK(net288),
    .D(\sr[247] ),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _1571_ (.CLK(net286),
    .D(\sr[248] ),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_1 _1572_ (.CLK(net287),
    .D(\sr[249] ),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_1 _1573_ (.CLK(net286),
    .D(\sr[250] ),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(net286),
    .D(\sr[251] ),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(net290),
    .D(\sr[252] ),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_2 _1576_ (.CLK(net282),
    .D(\sr[253] ),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(net286),
    .D(\sr[254] ),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(net291),
    .D(net260),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(clknet_leaf_1_sclk),
    .D(_0044_),
    .Q(\sr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(clknet_leaf_1_sclk),
    .D(_0045_),
    .Q(\sr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(clknet_leaf_1_sclk),
    .D(_0046_),
    .Q(\sr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(clknet_leaf_0_sclk),
    .D(_0047_),
    .Q(\sr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(clknet_leaf_0_sclk),
    .D(_0048_),
    .Q(\sr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(clknet_leaf_1_sclk),
    .D(_0049_),
    .Q(\sr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(clknet_leaf_0_sclk),
    .D(_0050_),
    .Q(\sr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(clknet_leaf_9_sclk),
    .D(_0051_),
    .Q(\sr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(clknet_leaf_9_sclk),
    .D(_0052_),
    .Q(\sr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(clknet_leaf_9_sclk),
    .D(_0053_),
    .Q(\sr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(clknet_leaf_9_sclk),
    .D(_0054_),
    .Q(\sr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(clknet_leaf_1_sclk),
    .D(_0055_),
    .Q(\sr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(clknet_leaf_1_sclk),
    .D(_0056_),
    .Q(\sr[12] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(latch),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(sdi),
    .X(net3));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(dq[0]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(dq[100]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(dq[101]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(dq[102]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(dq[103]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(dq[104]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dq[105]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dq[106]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dq[107]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dq[108]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dq[109]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dq[10]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dq[110]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dq[111]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dq[112]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dq[113]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dq[114]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dq[115]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dq[116]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dq[117]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dq[118]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dq[119]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dq[11]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dq[120]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dq[121]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dq[122]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dq[123]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dq[124]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(dq[125]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dq[126]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dq[127]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(dq[128]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(dq[129]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dq[12]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(dq[130]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(dq[131]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dq[132]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(dq[133]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(dq[134]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(dq[135]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(dq[136]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(dq[137]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(dq[138]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(dq[139]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(dq[13]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(dq[140]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(dq[141]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(dq[142]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(dq[143]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(dq[144]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(dq[145]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(dq[146]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(dq[147]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(dq[148]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(dq[149]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(dq[14]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(dq[150]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(dq[151]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(dq[152]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(dq[153]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(dq[154]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(dq[155]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(dq[156]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(dq[157]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(dq[158]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(dq[159]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(dq[15]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(dq[160]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(dq[161]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(dq[162]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(dq[163]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(dq[164]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(dq[165]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(dq[166]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(dq[167]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(dq[168]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(dq[169]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(dq[16]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(dq[170]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(dq[171]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(dq[172]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(dq[173]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(dq[174]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(dq[175]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(dq[176]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(dq[177]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(dq[178]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(dq[179]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(dq[17]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(dq[180]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(dq[181]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(dq[182]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(dq[183]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(dq[184]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(dq[185]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(dq[186]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(dq[187]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(dq[188]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(dq[189]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dq[18]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(dq[190]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(dq[191]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(dq[192]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(dq[193]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(dq[194]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(dq[195]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(dq[196]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(dq[197]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(dq[198]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(dq[199]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(dq[19]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(dq[1]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(dq[200]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(dq[201]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(dq[202]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(dq[203]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(dq[204]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(dq[205]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(dq[206]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(dq[207]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(dq[208]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(dq[209]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(dq[20]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(dq[210]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(dq[211]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(dq[212]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(dq[213]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(dq[214]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(dq[215]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(dq[216]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(dq[217]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(dq[218]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(dq[219]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(dq[21]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(dq[220]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(dq[221]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(dq[222]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(dq[223]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(dq[224]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(dq[225]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(dq[226]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(dq[227]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(dq[228]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(dq[229]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(dq[22]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(dq[230]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(dq[231]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(dq[232]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(dq[233]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(dq[234]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(dq[235]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(dq[236]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(dq[237]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(dq[238]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(dq[239]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(dq[23]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(dq[240]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(dq[241]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(dq[242]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(dq[243]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(dq[244]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(dq[245]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(dq[246]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(dq[247]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(dq[248]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(dq[249]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(dq[24]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(dq[250]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(dq[251]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(dq[252]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(dq[253]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(dq[254]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(dq[255]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(dq[25]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(dq[26]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(dq[27]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(dq[28]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(dq[29]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(dq[2]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(dq[30]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(dq[31]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(dq[32]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(dq[33]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(dq[34]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(dq[35]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(dq[36]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(dq[37]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(dq[38]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(dq[39]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(dq[3]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(dq[40]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(dq[41]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(dq[42]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(dq[43]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(dq[44]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(dq[45]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(dq[46]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(dq[47]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(dq[48]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(dq[49]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(dq[4]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(dq[50]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(dq[51]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(dq[52]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(dq[53]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(dq[54]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(dq[55]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(dq[56]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(dq[57]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(dq[58]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(dq[59]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(dq[5]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(dq[60]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(dq[61]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(dq[62]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(dq[63]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(dq[64]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(dq[65]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(dq[66]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(dq[67]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(dq[68]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(dq[69]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(dq[6]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(dq[70]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(dq[71]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(dq[72]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(dq[73]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(dq[74]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(dq[75]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(dq[76]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(dq[77]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(dq[78]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(dq[79]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(dq[7]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(dq[80]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(dq[81]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(dq[82]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(dq[83]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(dq[84]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(dq[85]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(dq[86]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(dq[87]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(dq[88]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(dq[89]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(dq[8]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(dq[90]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(dq[91]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(dq[92]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(dq[93]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(dq[94]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(dq[95]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(dq[96]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(dq[97]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(dq[98]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(dq[99]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(dq[9]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(sdo));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(net268),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net268),
    .X(net263));
 sky130_fd_sc_hd__buf_2 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(net268),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(net1),
    .X(net268));
 sky130_fd_sc_hd__buf_2 fanout269 (.A(net271),
    .X(net269));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_2 fanout271 (.A(net277),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 fanout273 (.A(net277),
    .X(net273));
 sky130_fd_sc_hd__buf_2 fanout274 (.A(net276),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_2 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net1),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 fanout280 (.A(net292),
    .X(net280));
 sky130_fd_sc_hd__buf_2 fanout281 (.A(net292),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(net292),
    .X(net282));
 sky130_fd_sc_hd__buf_2 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net292),
    .X(net284));
 sky130_fd_sc_hd__buf_2 fanout285 (.A(net292),
    .X(net285));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout286 (.A(net292),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(net291),
    .X(net287));
 sky130_fd_sc_hd__buf_2 fanout288 (.A(net291),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net1),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_sclk (.A(clknet_1_1__leaf_sclk),
    .X(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_sclk (.A(clknet_1_1__leaf_sclk),
    .X(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_sclk (.A(clknet_1_1__leaf_sclk),
    .X(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_sclk (.A(clknet_1_1__leaf_sclk),
    .X(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_sclk (.A(clknet_1_1__leaf_sclk),
    .X(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_sclk (.A(clknet_1_0__leaf_sclk),
    .X(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_sclk (.A(sclk),
    .X(clknet_0_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_sclk (.A(clknet_0_sclk),
    .X(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_sclk (.A(clknet_0_sclk),
    .X(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__D (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__D (.DIODE(_0031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__D (.DIODE(_0032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__D (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__D (.DIODE(_0148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__D (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__D (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__D (.DIODE(_0162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__D (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__D (.DIODE(_0167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__D (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__D (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__D (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__D (.DIODE(_0173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__D (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__D (.DIODE(_0178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__D (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__D (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__D (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__D (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__D (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__D (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__D (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__D (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__D (.DIODE(_0190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__D (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__D (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__D (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__D (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__D (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__D (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__D (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__D (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__D (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__D (.DIODE(_0213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__D (.DIODE(_0214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__D (.DIODE(_0215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__D (.DIODE(_0216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__D (.DIODE(_0217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__D (.DIODE(_0222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__D (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__D (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__D (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__D (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__D (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__D (.DIODE(_0243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__B (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0552__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__A (.DIODE(_0286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__A (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__A (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A (.DIODE(_0375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0930__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0951__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A (.DIODE(_0508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(latch));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_sclk_A (.DIODE(sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(sdi));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__D (.DIODE(\sr[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__B (.DIODE(\sr[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__D (.DIODE(\sr[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__B (.DIODE(\sr[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__D (.DIODE(\sr[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__B (.DIODE(\sr[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__D (.DIODE(\sr[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__B (.DIODE(\sr[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__D (.DIODE(\sr[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__B (.DIODE(\sr[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__D (.DIODE(\sr[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__B (.DIODE(\sr[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__D (.DIODE(\sr[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__B (.DIODE(\sr[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__D (.DIODE(\sr[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__B (.DIODE(\sr[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1334__D (.DIODE(\sr[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__B (.DIODE(\sr[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__D (.DIODE(\sr[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__B (.DIODE(\sr[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__D (.DIODE(\sr[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__B (.DIODE(\sr[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__D (.DIODE(\sr[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B (.DIODE(\sr[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__D (.DIODE(\sr[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__B (.DIODE(\sr[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__D (.DIODE(\sr[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B (.DIODE(\sr[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__D (.DIODE(\sr[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__B (.DIODE(\sr[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__D (.DIODE(\sr[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(\sr[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__D (.DIODE(\sr[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__B (.DIODE(\sr[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__D (.DIODE(\sr[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__B (.DIODE(\sr[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__D (.DIODE(\sr[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__B (.DIODE(\sr[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__D (.DIODE(\sr[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__B (.DIODE(\sr[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__D (.DIODE(\sr[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__B (.DIODE(\sr[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__D (.DIODE(\sr[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__B (.DIODE(\sr[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__D (.DIODE(\sr[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__B (.DIODE(\sr[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__D (.DIODE(\sr[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__B (.DIODE(\sr[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1460__D (.DIODE(\sr[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__B (.DIODE(\sr[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__D (.DIODE(\sr[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__B (.DIODE(\sr[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__D (.DIODE(\sr[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__B (.DIODE(\sr[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__D (.DIODE(\sr[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__B (.DIODE(\sr[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__D (.DIODE(\sr[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__B (.DIODE(\sr[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__D (.DIODE(\sr[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__B (.DIODE(\sr[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__D (.DIODE(\sr[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__B (.DIODE(\sr[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__D (.DIODE(\sr[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__B (.DIODE(\sr[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__D (.DIODE(\sr[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__B (.DIODE(\sr[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__D (.DIODE(\sr[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__B (.DIODE(\sr[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__D (.DIODE(\sr[147] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__B (.DIODE(\sr[147] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__D (.DIODE(\sr[148] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__B (.DIODE(\sr[148] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__D (.DIODE(\sr[149] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__B (.DIODE(\sr[149] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1337__D (.DIODE(\sr[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__B (.DIODE(\sr[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__D (.DIODE(\sr[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__B (.DIODE(\sr[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__D (.DIODE(\sr[151] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__B (.DIODE(\sr[151] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__D (.DIODE(\sr[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__B (.DIODE(\sr[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__D (.DIODE(\sr[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__B (.DIODE(\sr[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__D (.DIODE(\sr[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__B (.DIODE(\sr[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__D (.DIODE(\sr[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B (.DIODE(\sr[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__D (.DIODE(\sr[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__B (.DIODE(\sr[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__D (.DIODE(\sr[160] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__B (.DIODE(\sr[160] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__D (.DIODE(\sr[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__B (.DIODE(\sr[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__D (.DIODE(\sr[162] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B (.DIODE(\sr[162] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__D (.DIODE(\sr[163] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__B (.DIODE(\sr[163] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__D (.DIODE(\sr[164] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B (.DIODE(\sr[164] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__D (.DIODE(\sr[166] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__B (.DIODE(\sr[166] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__D (.DIODE(\sr[167] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__B (.DIODE(\sr[167] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__D (.DIODE(\sr[168] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B (.DIODE(\sr[168] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__D (.DIODE(\sr[169] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__B (.DIODE(\sr[169] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__D (.DIODE(\sr[170] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__B (.DIODE(\sr[170] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__D (.DIODE(\sr[171] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__B (.DIODE(\sr[171] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__D (.DIODE(\sr[172] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__B (.DIODE(\sr[172] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__D (.DIODE(\sr[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__B (.DIODE(\sr[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__D (.DIODE(\sr[180] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__B (.DIODE(\sr[180] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__D (.DIODE(\sr[181] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__B (.DIODE(\sr[181] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__D (.DIODE(\sr[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__B (.DIODE(\sr[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__D (.DIODE(\sr[183] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__B (.DIODE(\sr[183] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__D (.DIODE(\sr[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__B (.DIODE(\sr[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__D (.DIODE(\sr[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__B (.DIODE(\sr[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__D (.DIODE(\sr[190] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__B (.DIODE(\sr[190] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__D (.DIODE(\sr[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__B (.DIODE(\sr[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__D (.DIODE(\sr[199] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__B (.DIODE(\sr[199] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__D (.DIODE(\sr[202] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__B (.DIODE(\sr[202] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__D (.DIODE(\sr[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__B (.DIODE(\sr[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__D (.DIODE(\sr[209] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__B (.DIODE(\sr[209] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__D (.DIODE(\sr[213] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__B (.DIODE(\sr[213] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__D (.DIODE(\sr[219] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__B (.DIODE(\sr[219] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__D (.DIODE(\sr[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__B (.DIODE(\sr[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__D (.DIODE(\sr[220] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__B (.DIODE(\sr[220] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__D (.DIODE(\sr[221] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__B (.DIODE(\sr[221] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__D (.DIODE(\sr[222] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__B (.DIODE(\sr[222] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__D (.DIODE(\sr[223] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__B (.DIODE(\sr[223] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__D (.DIODE(\sr[224] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (.DIODE(\sr[224] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__D (.DIODE(\sr[225] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (.DIODE(\sr[225] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__D (.DIODE(\sr[226] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__B (.DIODE(\sr[226] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__D (.DIODE(\sr[227] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (.DIODE(\sr[227] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__D (.DIODE(\sr[228] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__B (.DIODE(\sr[228] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__D (.DIODE(\sr[229] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__B (.DIODE(\sr[229] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__D (.DIODE(\sr[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__B (.DIODE(\sr[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__D (.DIODE(\sr[230] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (.DIODE(\sr[230] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__D (.DIODE(\sr[231] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__B (.DIODE(\sr[231] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__D (.DIODE(\sr[232] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__B (.DIODE(\sr[232] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__D (.DIODE(\sr[233] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__B (.DIODE(\sr[233] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__D (.DIODE(\sr[234] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__B (.DIODE(\sr[234] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__D (.DIODE(\sr[235] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B (.DIODE(\sr[235] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__D (.DIODE(\sr[237] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__B (.DIODE(\sr[237] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__D (.DIODE(\sr[239] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__B (.DIODE(\sr[239] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__D (.DIODE(\sr[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__B (.DIODE(\sr[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__D (.DIODE(\sr[240] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__B (.DIODE(\sr[240] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__D (.DIODE(\sr[242] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__B (.DIODE(\sr[242] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__D (.DIODE(\sr[244] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B (.DIODE(\sr[244] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__D (.DIODE(\sr[247] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B (.DIODE(\sr[247] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__D (.DIODE(\sr[248] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B (.DIODE(\sr[248] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__D (.DIODE(\sr[249] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__B (.DIODE(\sr[249] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__D (.DIODE(\sr[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__B (.DIODE(\sr[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__D (.DIODE(\sr[250] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B (.DIODE(\sr[250] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__D (.DIODE(\sr[251] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B (.DIODE(\sr[251] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__D (.DIODE(\sr[252] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__B (.DIODE(\sr[252] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__D (.DIODE(\sr[254] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__B (.DIODE(\sr[254] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1348__D (.DIODE(\sr[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__B (.DIODE(\sr[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__D (.DIODE(\sr[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__B (.DIODE(\sr[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__D (.DIODE(\sr[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__B (.DIODE(\sr[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__D (.DIODE(\sr[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__B (.DIODE(\sr[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__D (.DIODE(\sr[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__B (.DIODE(\sr[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__D (.DIODE(\sr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__B (.DIODE(\sr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__D (.DIODE(\sr[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__B (.DIODE(\sr[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__D (.DIODE(\sr[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__B (.DIODE(\sr[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__D (.DIODE(\sr[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__B (.DIODE(\sr[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__D (.DIODE(\sr[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__B (.DIODE(\sr[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__D (.DIODE(\sr[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__B (.DIODE(\sr[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__D (.DIODE(\sr[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__B (.DIODE(\sr[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__D (.DIODE(\sr[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__B (.DIODE(\sr[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__D (.DIODE(\sr[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__B (.DIODE(\sr[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__D (.DIODE(\sr[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__B (.DIODE(\sr[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__D (.DIODE(\sr[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__B (.DIODE(\sr[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__D (.DIODE(\sr[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__B (.DIODE(\sr[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__D (.DIODE(\sr[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__B (.DIODE(\sr[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__D (.DIODE(\sr[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__B (.DIODE(\sr[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__D (.DIODE(\sr[68] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__B (.DIODE(\sr[68] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__D (.DIODE(\sr[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__B (.DIODE(\sr[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__D (.DIODE(\sr[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B (.DIODE(\sr[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__D (.DIODE(\sr[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B (.DIODE(\sr[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__D (.DIODE(\sr[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B (.DIODE(\sr[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__D (.DIODE(\sr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__B (.DIODE(\sr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__D (.DIODE(\sr[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__B (.DIODE(\sr[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__D (.DIODE(\sr[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__B (.DIODE(\sr[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__D (.DIODE(\sr[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__B (.DIODE(\sr[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__D (.DIODE(\sr[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B (.DIODE(\sr[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__D (.DIODE(\sr[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__B (.DIODE(\sr[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_output9_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_output12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_output13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_output231_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_output236_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_output237_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_output238_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_output239_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_output248_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__D (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__CLK (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__CLK (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__CLK (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__CLK (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__CLK (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__CLK (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__CLK (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__CLK (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__CLK (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__CLK (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__CLK (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__CLK (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__CLK (.DIODE(clknet_leaf_0_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__CLK (.DIODE(clknet_leaf_1_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1316__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__CLK (.DIODE(clknet_leaf_2_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__CLK (.DIODE(clknet_leaf_3_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1279__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1298__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1282__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1292__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__CLK (.DIODE(clknet_leaf_4_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1220__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__CLK (.DIODE(clknet_leaf_5_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1295__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__CLK (.DIODE(clknet_leaf_6_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1294__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__CLK (.DIODE(clknet_leaf_7_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__CLK (.DIODE(clknet_leaf_8_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__CLK (.DIODE(clknet_leaf_9_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__CLK (.DIODE(clknet_leaf_10_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_sclk_A (.DIODE(clknet_1_0__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_sclk_A (.DIODE(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_sclk_A (.DIODE(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_sclk_A (.DIODE(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_sclk_A (.DIODE(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_sclk_A (.DIODE(clknet_1_1__leaf_sclk));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1454 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1476 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1517 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1545 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1632 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1644 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1659 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1678 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1691 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1698 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1448 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1472 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1515 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1529 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1538 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1551 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1571 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1594 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1618 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1639 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1650 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1675 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1695 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1702 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1374 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1472 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1484 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1545 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1576 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1598 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1644 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1670 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1702 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1394 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1517 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1572 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1592 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1662 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1669 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1673 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1686 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1700 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1706 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1307 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1424 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1430 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1471 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1488 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1532 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1552 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1587 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1643 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1659 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1667 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1702 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1416 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1424 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1434 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1452 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1458 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1464 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1624 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1631 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1639 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1646 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1672 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1690 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1704 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1327 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1424 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1430 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1471 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1492 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1498 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1543 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1639 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1650 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1656 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1669 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1702 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1443 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1491 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1503 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1507 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1514 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1584 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1672 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1690 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1704 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1480 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1510 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1546 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1566 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1575 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1615 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1643 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1668 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1494 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1512 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1559 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1592 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1637 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1646 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1666 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1700 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1706 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1367 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1471 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1489 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1518 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1545 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1644 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1654 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1688 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1697 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1351 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1448 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1458 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1472 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1503 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1559 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1587 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1621 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1639 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1660 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1669 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1678 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1696 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1263 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1471 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1503 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1523 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1529 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1546 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1566 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1588 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1608 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1623 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1631 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1648 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1666 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1710 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1482 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1492 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1498 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1504 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1517 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1562 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1582 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1650 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1676 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1685 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1694 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1431 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1451 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1508 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1519 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1558 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1643 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1387 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1451 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1482 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1526 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1530 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1536 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1563 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1583 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1604 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1608 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1626 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1646 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1680 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1696 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1433 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1475 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1542 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1643 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1697 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1415 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1433 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1499 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1560 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1611 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1634 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1641 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1680 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1688 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1696 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1391 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1415 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1477 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1499 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1535 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1543 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1643 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1702 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1471 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1499 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1527 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1545 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1573 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1659 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1667 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1709 ();
endmodule

