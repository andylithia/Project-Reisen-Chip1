magic
tech sky130A
magscale 1 2
timestamp 1671331890
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 4 49 845 248
rect 0 0 196 49
rect 204 48 388 49
rect 396 48 580 49
rect 588 48 772 49
rect 780 48 933 49
rect 205 0 388 48
rect 397 0 580 48
rect 589 0 772 48
rect 781 0 933 48
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 278 368 308 592
rect 368 368 398 592
rect 470 368 500 592
rect 560 368 590 592
rect 662 368 692 592
rect 752 368 782 592
<< nmoslvt >>
rect 87 74 117 222
rect 173 74 206 222
rect 279 74 309 222
rect 365 74 398 222
rect 471 74 501 222
rect 557 74 590 222
rect 663 74 693 222
rect 749 74 782 222
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 210 173 222
rect 117 176 128 210
rect 162 176 173 210
rect 117 120 173 176
rect 117 86 128 120
rect 162 86 173 120
rect 117 74 173 86
rect 206 210 279 222
rect 206 176 234 210
rect 268 176 279 210
rect 206 120 279 176
rect 206 86 234 120
rect 268 86 279 120
rect 206 74 279 86
rect 309 210 365 222
rect 309 176 320 210
rect 354 176 365 210
rect 309 120 365 176
rect 309 86 320 120
rect 354 86 365 120
rect 309 74 365 86
rect 398 210 471 222
rect 398 176 426 210
rect 460 176 471 210
rect 398 120 471 176
rect 398 86 426 120
rect 460 86 471 120
rect 398 74 471 86
rect 501 210 557 222
rect 501 176 512 210
rect 546 176 557 210
rect 501 120 557 176
rect 501 86 512 120
rect 546 86 557 120
rect 501 74 557 86
rect 590 210 663 222
rect 590 176 618 210
rect 652 176 663 210
rect 590 120 663 176
rect 590 86 618 120
rect 652 86 663 120
rect 590 74 663 86
rect 693 210 749 222
rect 693 176 704 210
rect 738 176 749 210
rect 693 120 749 176
rect 693 86 704 120
rect 738 86 749 120
rect 693 74 749 86
rect 782 74 812 222
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 510 176 546
rect 116 476 129 510
rect 163 476 176 510
rect 116 440 176 476
rect 116 406 129 440
rect 163 406 176 440
rect 116 368 176 406
rect 206 580 278 592
rect 206 546 231 580
rect 265 546 278 580
rect 206 497 278 546
rect 206 463 231 497
rect 265 463 278 497
rect 206 414 278 463
rect 206 380 231 414
rect 265 380 278 414
rect 206 368 278 380
rect 308 580 368 592
rect 308 546 321 580
rect 355 546 368 580
rect 308 510 368 546
rect 308 476 321 510
rect 355 476 368 510
rect 308 440 368 476
rect 308 406 321 440
rect 355 406 368 440
rect 308 368 368 406
rect 398 580 470 592
rect 398 546 423 580
rect 457 546 470 580
rect 398 497 470 546
rect 398 463 423 497
rect 457 463 470 497
rect 398 414 470 463
rect 398 380 423 414
rect 457 380 470 414
rect 398 368 470 380
rect 500 580 560 592
rect 500 546 513 580
rect 547 546 560 580
rect 500 510 560 546
rect 500 476 513 510
rect 547 476 560 510
rect 500 440 560 476
rect 500 406 513 440
rect 547 406 560 440
rect 500 368 560 406
rect 590 580 662 592
rect 590 546 615 580
rect 649 546 662 580
rect 590 497 662 546
rect 590 463 615 497
rect 649 463 662 497
rect 590 414 662 463
rect 590 380 615 414
rect 649 380 662 414
rect 590 368 662 380
rect 692 580 752 592
rect 692 546 705 580
rect 739 546 752 580
rect 692 510 752 546
rect 692 476 705 510
rect 739 476 752 510
rect 692 440 752 476
rect 692 406 705 440
rect 739 406 752 440
rect 692 368 752 406
rect 782 368 832 592
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 176 162 210
rect 128 86 162 120
rect 234 176 268 210
rect 234 86 268 120
rect 320 176 354 210
rect 320 86 354 120
rect 426 176 460 210
rect 426 86 460 120
rect 512 176 546 210
rect 512 86 546 120
rect 618 176 652 210
rect 618 86 652 120
rect 704 176 738 210
rect 704 86 738 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 476 163 510
rect 129 406 163 440
rect 231 546 265 580
rect 231 463 265 497
rect 231 380 265 414
rect 321 546 355 580
rect 321 476 355 510
rect 321 406 355 440
rect 423 546 457 580
rect 423 463 457 497
rect 423 380 457 414
rect 513 546 547 580
rect 513 476 547 510
rect 513 406 547 440
rect 615 546 649 580
rect 615 463 649 497
rect 615 380 649 414
rect 705 546 739 580
rect 705 476 739 510
rect 705 406 739 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 278 592 308 618
rect 368 592 398 618
rect 470 592 500 618
rect 560 592 590 618
rect 662 592 692 618
rect 752 592 782 618
rect 869 372 927 388
rect 86 353 116 368
rect 176 353 206 368
rect 278 353 308 368
rect 368 353 398 368
rect 470 353 500 368
rect 560 353 590 368
rect 662 353 692 368
rect 752 353 782 368
rect 869 353 879 372
rect 83 334 879 353
rect 917 334 927 372
rect 83 314 927 334
rect 83 252 899 272
rect 83 240 851 252
rect 87 222 117 240
rect 173 222 206 240
rect 279 222 309 240
rect 365 222 398 240
rect 471 222 501 240
rect 557 222 590 240
rect 663 222 693 240
rect 749 222 782 240
rect 841 214 851 240
rect 889 214 899 252
rect 841 198 899 214
rect 87 48 117 74
rect 173 48 206 74
rect 279 48 309 74
rect 365 48 398 74
rect 471 48 501 74
rect 557 48 590 74
rect 663 48 693 74
rect 749 48 782 74
<< polycont >>
rect 879 334 917 372
rect 851 214 889 252
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 864 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 497 73 546
rect 23 476 39 497
rect 23 442 34 476
rect 68 442 73 463
rect 23 414 73 442
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 163 596
rect 113 555 129 580
rect 113 521 124 555
rect 158 521 163 546
rect 113 510 163 521
rect 113 476 129 510
rect 113 440 163 476
rect 113 406 129 440
rect 113 364 163 406
rect 215 580 265 596
rect 215 546 231 580
rect 215 497 265 546
rect 215 476 231 497
rect 215 442 226 476
rect 260 442 265 463
rect 215 414 265 442
rect 215 380 231 414
rect 215 364 265 380
rect 305 580 355 596
rect 305 555 321 580
rect 305 521 316 555
rect 350 521 355 546
rect 305 510 355 521
rect 305 476 321 510
rect 305 440 355 476
rect 305 406 321 440
rect 305 364 355 406
rect 407 580 457 596
rect 407 546 423 580
rect 407 497 457 546
rect 407 476 423 497
rect 407 442 418 476
rect 452 442 457 463
rect 407 414 457 442
rect 407 380 423 414
rect 407 364 457 380
rect 497 580 547 596
rect 497 555 513 580
rect 497 521 508 555
rect 542 521 547 546
rect 497 510 547 521
rect 497 476 513 510
rect 497 440 547 476
rect 497 406 513 440
rect 497 364 547 406
rect 599 580 649 596
rect 599 546 615 580
rect 599 497 649 546
rect 599 476 615 497
rect 599 442 610 476
rect 644 442 649 463
rect 599 414 649 442
rect 599 380 615 414
rect 599 364 649 380
rect 689 580 739 596
rect 689 555 705 580
rect 689 521 700 555
rect 734 521 739 546
rect 689 510 739 521
rect 689 476 705 510
rect 689 440 739 476
rect 689 406 705 440
rect 689 364 739 406
rect 863 334 879 372
rect 917 334 933 372
rect 26 216 76 226
rect 26 182 37 216
rect 71 210 76 216
rect 26 176 42 182
rect 26 120 76 176
rect 26 86 42 120
rect 26 70 76 86
rect 112 210 162 226
rect 112 176 128 210
rect 112 126 162 176
rect 112 92 123 126
rect 157 120 162 126
rect 112 86 128 92
rect 112 70 162 86
rect 218 216 268 226
rect 218 182 229 216
rect 263 210 268 216
rect 218 176 234 182
rect 218 120 268 176
rect 218 86 234 120
rect 218 70 268 86
rect 304 210 354 226
rect 304 176 320 210
rect 304 126 354 176
rect 304 92 315 126
rect 349 120 354 126
rect 304 86 320 92
rect 304 70 354 86
rect 410 216 460 226
rect 410 182 421 216
rect 455 210 460 216
rect 410 176 426 182
rect 410 120 460 176
rect 410 86 426 120
rect 410 70 460 86
rect 496 210 546 226
rect 496 176 512 210
rect 496 126 546 176
rect 496 92 507 126
rect 541 120 546 126
rect 496 86 512 92
rect 496 70 546 86
rect 602 216 652 226
rect 602 182 613 216
rect 647 210 652 216
rect 602 176 618 182
rect 602 120 652 176
rect 602 86 618 120
rect 602 70 652 86
rect 688 210 738 226
rect 835 214 851 252
rect 889 214 905 252
rect 688 176 704 210
rect 688 126 738 176
rect 688 92 699 126
rect 733 120 738 126
rect 688 86 704 92
rect 688 70 738 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 935 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 34 463 39 476
rect 39 463 68 476
rect 34 442 68 463
rect 124 546 129 555
rect 129 546 158 555
rect 124 521 158 546
rect 226 463 231 476
rect 231 463 260 476
rect 226 442 260 463
rect 316 546 321 555
rect 321 546 350 555
rect 316 521 350 546
rect 418 463 423 476
rect 423 463 452 476
rect 418 442 452 463
rect 508 546 513 555
rect 513 546 542 555
rect 508 521 542 546
rect 610 463 615 476
rect 615 463 644 476
rect 610 442 644 463
rect 700 546 705 555
rect 705 546 734 555
rect 700 521 734 546
rect 37 210 71 216
rect 37 182 42 210
rect 42 182 71 210
rect 123 120 157 126
rect 123 92 128 120
rect 128 92 157 120
rect 229 210 263 216
rect 229 182 234 210
rect 234 182 263 210
rect 315 120 349 126
rect 315 92 320 120
rect 320 92 349 120
rect 421 210 455 216
rect 421 182 426 210
rect 426 182 455 210
rect 507 120 541 126
rect 507 92 512 120
rect 512 92 541 120
rect 613 210 647 216
rect 613 182 618 210
rect 618 182 647 210
rect 699 120 733 126
rect 699 92 704 120
rect 704 92 733 120
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 864 683
rect 0 617 864 649
rect 23 555 746 561
rect 23 521 124 555
rect 158 521 316 555
rect 350 521 508 555
rect 542 521 700 555
rect 734 521 746 555
rect 23 515 746 521
rect 22 476 659 482
rect 22 442 34 476
rect 68 442 226 476
rect 260 442 418 476
rect 452 442 610 476
rect 644 442 659 476
rect 22 436 659 442
rect 609 222 659 436
rect 25 216 659 222
rect 25 182 37 216
rect 71 182 229 216
rect 263 182 421 216
rect 455 182 613 216
rect 647 182 659 216
rect 25 176 659 182
rect 699 132 746 515
rect 25 126 746 132
rect 25 92 123 126
rect 157 92 315 126
rect 349 92 507 126
rect 541 92 699 126
rect 733 92 746 126
rect 25 86 746 92
rect 0 17 935 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 935 17
rect 0 -49 935 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_8
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 1 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 2 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 3 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
<< end >>
