magic
tech sky130A
magscale 1 2
timestamp 1671648335
<< error_s >>
rect 3640 4874 3698 4880
rect 3832 4874 3890 4880
rect 4024 4874 4082 4880
rect 4216 4874 4274 4880
rect 3640 4840 3652 4874
rect 3832 4840 3844 4874
rect 4024 4840 4036 4874
rect 4216 4840 4228 4874
rect 3640 4834 3698 4840
rect 3832 4834 3890 4840
rect 4024 4834 4082 4840
rect 4216 4834 4274 4840
rect 3544 4346 3602 4352
rect 3736 4346 3794 4352
rect 3928 4346 3986 4352
rect 4120 4346 4178 4352
rect 3544 4312 3556 4346
rect 3736 4312 3748 4346
rect 3928 4312 3940 4346
rect 4120 4312 4132 4346
rect 3544 4306 3602 4312
rect 3736 4306 3794 4312
rect 3928 4306 3986 4312
rect 4120 4306 4178 4312
rect 3640 3986 3698 3992
rect 3832 3986 3890 3992
rect 4024 3986 4082 3992
rect 4216 3986 4274 3992
rect 3640 3952 3652 3986
rect 3832 3952 3844 3986
rect 4024 3952 4036 3986
rect 4216 3952 4228 3986
rect 3640 3946 3698 3952
rect 3832 3946 3890 3952
rect 4024 3946 4082 3952
rect 4216 3946 4274 3952
rect 3544 3676 3602 3682
rect 3736 3676 3794 3682
rect 3928 3676 3986 3682
rect 4120 3676 4178 3682
rect 3544 3642 3556 3676
rect 3736 3642 3748 3676
rect 3928 3642 3940 3676
rect 4120 3642 4132 3676
rect 3544 3636 3602 3642
rect 3736 3636 3794 3642
rect 3928 3636 3986 3642
rect 4120 3636 4178 3642
rect 4062 1800 4100 1818
rect 4062 1750 4072 1768
rect 4934 1670 4972 1688
rect 4962 1620 4972 1638
<< dnwell >>
rect 3475 682 5555 2994
<< nwell >>
rect 3395 2788 5635 3074
rect 3395 888 3681 2788
rect 3935 1696 5095 2534
rect 5349 888 5635 2788
rect 3395 602 5635 888
<< pwell >>
rect 3935 1076 5095 1696
<< nmos >>
rect 4131 1286 4191 1486
rect 4249 1286 4309 1486
rect 4367 1286 4427 1486
rect 4485 1286 4545 1486
rect 4603 1286 4663 1486
rect 4721 1286 4781 1486
rect 4839 1286 4899 1486
<< pmos >>
rect 4131 1915 4191 2315
rect 4249 1915 4309 2315
rect 4367 1915 4427 2315
rect 4485 1915 4545 2315
rect 4603 1915 4663 2315
rect 4721 1915 4781 2315
rect 4839 1915 4899 2315
<< ndiff >>
rect 4073 1474 4131 1486
rect 4073 1298 4085 1474
rect 4119 1298 4131 1474
rect 4073 1286 4131 1298
rect 4191 1474 4249 1486
rect 4191 1298 4203 1474
rect 4237 1298 4249 1474
rect 4191 1286 4249 1298
rect 4309 1474 4367 1486
rect 4309 1298 4321 1474
rect 4355 1298 4367 1474
rect 4309 1286 4367 1298
rect 4427 1474 4485 1486
rect 4427 1298 4439 1474
rect 4473 1298 4485 1474
rect 4427 1286 4485 1298
rect 4545 1474 4603 1486
rect 4545 1298 4557 1474
rect 4591 1298 4603 1474
rect 4545 1286 4603 1298
rect 4663 1474 4721 1486
rect 4663 1298 4675 1474
rect 4709 1298 4721 1474
rect 4663 1286 4721 1298
rect 4781 1474 4839 1486
rect 4781 1298 4793 1474
rect 4827 1298 4839 1474
rect 4781 1286 4839 1298
rect 4899 1474 4957 1486
rect 4899 1298 4911 1474
rect 4945 1298 4957 1474
rect 4899 1286 4957 1298
<< pdiff >>
rect 4073 2303 4131 2315
rect 4073 1927 4085 2303
rect 4119 1927 4131 2303
rect 4073 1915 4131 1927
rect 4191 2303 4249 2315
rect 4191 1927 4203 2303
rect 4237 1927 4249 2303
rect 4191 1915 4249 1927
rect 4309 2303 4367 2315
rect 4309 1927 4321 2303
rect 4355 1927 4367 2303
rect 4309 1915 4367 1927
rect 4427 2303 4485 2315
rect 4427 1927 4439 2303
rect 4473 1927 4485 2303
rect 4427 1915 4485 1927
rect 4545 2303 4603 2315
rect 4545 1927 4557 2303
rect 4591 1927 4603 2303
rect 4545 1915 4603 1927
rect 4663 2303 4721 2315
rect 4663 1927 4675 2303
rect 4709 1927 4721 2303
rect 4663 1915 4721 1927
rect 4781 2303 4839 2315
rect 4781 1927 4793 2303
rect 4827 1927 4839 2303
rect 4781 1915 4839 1927
rect 4899 2303 4957 2315
rect 4899 1927 4911 2303
rect 4945 1927 4957 2303
rect 4899 1915 4957 1927
<< ndiffc >>
rect 4085 1298 4119 1474
rect 4203 1298 4237 1474
rect 4321 1298 4355 1474
rect 4439 1298 4473 1474
rect 4557 1298 4591 1474
rect 4675 1298 4709 1474
rect 4793 1298 4827 1474
rect 4911 1298 4945 1474
<< pdiffc >>
rect 4085 1927 4119 2303
rect 4203 1927 4237 2303
rect 4321 1927 4355 2303
rect 4439 1927 4473 2303
rect 4557 1927 4591 2303
rect 4675 1927 4709 2303
rect 4793 1927 4827 2303
rect 4911 1927 4945 2303
<< psubdiff >>
rect 3971 1626 4067 1660
rect 4972 1626 5059 1660
rect 3971 1564 4005 1626
rect 5025 1564 5059 1626
rect 3971 1146 4005 1208
rect 5025 1146 5059 1208
rect 3971 1112 4067 1146
rect 4963 1112 5059 1146
<< nsubdiff >>
rect 3432 3017 5598 3037
rect 3432 2983 3512 3017
rect 5518 2983 5598 3017
rect 3432 2963 5598 2983
rect 3432 2957 3506 2963
rect 3432 719 3452 2957
rect 3486 719 3506 2957
rect 5524 2957 5598 2963
rect 3971 2464 4067 2498
rect 4963 2464 5059 2498
rect 3971 2402 4005 2464
rect 5025 2402 5059 2464
rect 3971 1766 4005 1828
rect 5025 1766 5059 1828
rect 3971 1732 4067 1766
rect 4963 1732 5059 1766
rect 3432 713 3506 719
rect 5524 719 5544 2957
rect 5578 719 5598 2957
rect 5524 713 5598 719
rect 3432 693 5598 713
rect 3432 659 3512 693
rect 5518 659 5598 693
rect 3432 639 5598 659
<< psubdiffcont >>
rect 4067 1626 4972 1660
rect 3971 1208 4005 1564
rect 5025 1208 5059 1564
rect 4067 1112 4963 1146
<< nsubdiffcont >>
rect 3512 2983 5518 3017
rect 3452 719 3486 2957
rect 4067 2464 4963 2498
rect 3971 1828 4005 2402
rect 5025 1828 5059 2402
rect 4067 1732 4963 1766
rect 5544 719 5578 2957
rect 3512 659 5518 693
<< poly >>
rect 4128 2396 4194 2412
rect 4128 2362 4144 2396
rect 4178 2362 4194 2396
rect 4128 2346 4194 2362
rect 4246 2396 4312 2412
rect 4246 2362 4262 2396
rect 4296 2362 4312 2396
rect 4246 2346 4312 2362
rect 4364 2396 4430 2412
rect 4364 2362 4380 2396
rect 4414 2362 4430 2396
rect 4364 2346 4430 2362
rect 4482 2396 4548 2412
rect 4482 2362 4498 2396
rect 4532 2362 4548 2396
rect 4482 2346 4548 2362
rect 4600 2396 4666 2412
rect 4600 2362 4616 2396
rect 4650 2362 4666 2396
rect 4600 2346 4666 2362
rect 4718 2396 4784 2412
rect 4718 2362 4734 2396
rect 4768 2362 4784 2396
rect 4718 2346 4784 2362
rect 4836 2396 4902 2412
rect 4836 2362 4852 2396
rect 4886 2362 4902 2396
rect 4836 2346 4902 2362
rect 4131 2315 4191 2346
rect 4249 2315 4309 2346
rect 4367 2315 4427 2346
rect 4485 2315 4545 2346
rect 4603 2315 4663 2346
rect 4721 2315 4781 2346
rect 4839 2315 4899 2346
rect 4131 1884 4191 1915
rect 4249 1884 4309 1915
rect 4367 1884 4427 1915
rect 4485 1884 4545 1915
rect 4603 1884 4663 1915
rect 4721 1884 4781 1915
rect 4839 1884 4899 1915
rect 4128 1818 4194 1884
rect 4246 1818 4312 1884
rect 4364 1818 4430 1884
rect 4482 1818 4548 1884
rect 4600 1818 4666 1884
rect 4718 1818 4784 1884
rect 4836 1818 4902 1884
rect 4128 1508 4194 1574
rect 4246 1508 4312 1574
rect 4364 1508 4430 1574
rect 4482 1508 4548 1574
rect 4600 1508 4666 1574
rect 4718 1508 4784 1574
rect 4836 1508 4902 1574
rect 4131 1486 4191 1508
rect 4249 1486 4309 1508
rect 4367 1486 4427 1508
rect 4485 1486 4545 1508
rect 4603 1486 4663 1508
rect 4721 1486 4781 1508
rect 4839 1486 4899 1508
rect 4131 1264 4191 1286
rect 4249 1264 4309 1286
rect 4367 1264 4427 1286
rect 4485 1264 4545 1286
rect 4603 1264 4663 1286
rect 4721 1264 4781 1286
rect 4839 1264 4899 1286
rect 4128 1248 4194 1264
rect 4128 1214 4144 1248
rect 4178 1214 4194 1248
rect 4128 1198 4194 1214
rect 4246 1248 4312 1264
rect 4246 1214 4262 1248
rect 4296 1214 4312 1248
rect 4246 1198 4312 1214
rect 4364 1248 4430 1264
rect 4364 1214 4380 1248
rect 4414 1214 4430 1248
rect 4364 1198 4430 1214
rect 4482 1248 4548 1264
rect 4482 1214 4498 1248
rect 4532 1214 4548 1248
rect 4482 1198 4548 1214
rect 4600 1248 4666 1264
rect 4600 1214 4616 1248
rect 4650 1214 4666 1248
rect 4600 1198 4666 1214
rect 4718 1248 4784 1264
rect 4718 1214 4734 1248
rect 4768 1214 4784 1248
rect 4718 1198 4784 1214
rect 4836 1248 4902 1264
rect 4836 1214 4852 1248
rect 4886 1214 4902 1248
rect 4836 1198 4902 1214
<< polycont >>
rect 4144 2362 4178 2396
rect 4262 2362 4296 2396
rect 4380 2362 4414 2396
rect 4498 2362 4532 2396
rect 4616 2362 4650 2396
rect 4734 2362 4768 2396
rect 4852 2362 4886 2396
rect 4144 1214 4178 1248
rect 4262 1214 4296 1248
rect 4380 1214 4414 1248
rect 4498 1214 4532 1248
rect 4616 1214 4650 1248
rect 4734 1214 4768 1248
rect 4852 1214 4886 1248
<< locali >>
rect 3452 2983 3512 3017
rect 5518 2983 5578 3017
rect 3452 2957 3486 2983
rect 5544 2957 5578 2983
rect 3971 2521 5060 2534
rect 3971 2480 4006 2521
rect 5025 2480 5060 2521
rect 3971 2464 4067 2480
rect 4963 2464 5060 2480
rect 3971 2402 4005 2464
rect 5025 2402 5059 2464
rect 4128 2362 4144 2396
rect 4178 2362 4194 2396
rect 4246 2362 4262 2396
rect 4296 2362 4312 2396
rect 4364 2362 4380 2396
rect 4414 2362 4430 2396
rect 4482 2362 4498 2396
rect 4532 2362 4548 2396
rect 4600 2362 4616 2396
rect 4650 2362 4666 2396
rect 4718 2362 4734 2396
rect 4768 2362 4784 2396
rect 4836 2362 4852 2396
rect 4886 2362 4902 2396
rect 4085 2303 4119 2319
rect 4085 1911 4119 1927
rect 4203 2303 4237 2319
rect 4203 1911 4237 1927
rect 4321 2303 4355 2319
rect 4321 1911 4355 1927
rect 4439 2303 4473 2319
rect 4439 1911 4473 1927
rect 4557 2303 4591 2319
rect 4557 1911 4591 1927
rect 4675 2303 4709 2319
rect 4675 1911 4709 1927
rect 4793 2303 4827 2319
rect 4793 1911 4827 1927
rect 4911 2303 4945 2319
rect 4911 1911 4945 1927
rect 3971 1766 4005 1828
rect 5025 1766 5059 1828
rect 3971 1732 4067 1766
rect 4963 1732 5059 1766
rect 3971 1626 4067 1660
rect 4972 1626 5059 1660
rect 3971 1564 4005 1626
rect 5025 1564 5059 1626
rect 4085 1474 4119 1490
rect 4085 1282 4119 1298
rect 4203 1474 4237 1490
rect 4203 1282 4237 1298
rect 4321 1474 4355 1490
rect 4321 1282 4355 1298
rect 4439 1474 4473 1490
rect 4439 1282 4473 1298
rect 4557 1474 4591 1490
rect 4557 1282 4591 1298
rect 4675 1474 4709 1490
rect 4675 1282 4709 1298
rect 4793 1474 4827 1490
rect 4793 1282 4827 1298
rect 4911 1474 4945 1490
rect 4911 1282 4945 1298
rect 4128 1214 4144 1248
rect 4178 1214 4194 1248
rect 4246 1214 4262 1248
rect 4296 1214 4312 1248
rect 4364 1214 4380 1248
rect 4414 1214 4430 1248
rect 4482 1214 4498 1248
rect 4532 1214 4548 1248
rect 4600 1214 4616 1248
rect 4650 1214 4666 1248
rect 4718 1214 4734 1248
rect 4768 1214 4784 1248
rect 4836 1214 4852 1248
rect 4886 1214 4902 1248
rect 3971 1146 4005 1208
rect 5025 1146 5059 1208
rect 3971 1130 4067 1146
rect 4963 1130 5059 1146
rect 3971 1112 4012 1130
rect 5012 1112 5059 1130
rect 3992 1090 4012 1112
rect 5012 1090 5032 1112
rect 3992 1070 5032 1090
rect 3452 693 3486 719
rect 5544 693 5578 719
rect 3452 659 3512 693
rect 5518 659 5578 693
<< viali >>
rect 4006 2498 5025 2521
rect 4006 2480 4067 2498
rect 4067 2480 4963 2498
rect 4963 2480 5025 2498
rect 4144 2362 4178 2396
rect 4262 2362 4296 2396
rect 4380 2362 4414 2396
rect 4498 2362 4532 2396
rect 4616 2362 4650 2396
rect 4734 2362 4768 2396
rect 4852 2362 4886 2396
rect 4085 1927 4119 2303
rect 4203 1927 4237 2303
rect 4321 1927 4355 2303
rect 4439 1927 4473 2303
rect 4557 1927 4591 2303
rect 4675 1927 4709 2303
rect 4793 1927 4827 2303
rect 4911 1927 4945 2303
rect 4085 1298 4119 1474
rect 4203 1298 4237 1474
rect 4321 1298 4355 1474
rect 4439 1298 4473 1474
rect 4557 1298 4591 1474
rect 4675 1298 4709 1474
rect 4793 1298 4827 1474
rect 4911 1298 4945 1474
rect 4144 1214 4178 1248
rect 4262 1214 4296 1248
rect 4380 1214 4414 1248
rect 4498 1214 4532 1248
rect 4616 1214 4650 1248
rect 4734 1214 4768 1248
rect 4852 1214 4886 1248
rect 4012 1112 4067 1130
rect 4067 1112 4963 1130
rect 4963 1112 5012 1130
rect 4012 1090 5012 1112
<< metal1 >>
rect 3971 2464 4005 2534
rect 4477 2521 5060 2534
rect 5025 2480 5060 2521
rect 4477 2464 5060 2480
rect 4132 2396 4898 2402
rect 4132 2362 4144 2396
rect 4178 2362 4262 2396
rect 4296 2362 4380 2396
rect 4414 2362 4498 2396
rect 4532 2362 4616 2396
rect 4650 2362 4734 2396
rect 4768 2362 4852 2396
rect 4886 2362 4898 2396
rect 4132 2356 4898 2362
rect 4079 2303 4125 2315
rect 4079 1927 4085 2303
rect 4119 1927 4125 2303
rect 4079 1800 4125 1927
rect 4197 2303 4243 2315
rect 4197 1927 4203 2303
rect 4237 1927 4243 2303
rect 4062 1740 4072 1800
rect 4132 1740 4142 1800
rect 4079 1474 4125 1740
rect 4197 1670 4243 1927
rect 4315 2303 4361 2315
rect 4315 1927 4321 2303
rect 4355 1927 4361 2303
rect 4315 1800 4361 1927
rect 4433 2303 4479 2315
rect 4433 1927 4439 2303
rect 4473 1927 4479 2303
rect 4302 1740 4312 1800
rect 4372 1740 4382 1800
rect 4172 1610 4182 1670
rect 4242 1610 4252 1670
rect 4079 1298 4085 1474
rect 4119 1298 4125 1474
rect 4079 1286 4125 1298
rect 4197 1474 4243 1610
rect 4197 1298 4203 1474
rect 4237 1298 4243 1474
rect 4197 1286 4243 1298
rect 4315 1474 4361 1740
rect 4433 1670 4479 1927
rect 4551 2303 4597 2315
rect 4551 1927 4557 2303
rect 4591 1927 4597 2303
rect 4551 1800 4597 1927
rect 4669 2303 4715 2315
rect 4669 1927 4675 2303
rect 4709 1927 4715 2303
rect 4532 1740 4542 1800
rect 4602 1740 4612 1800
rect 4422 1610 4432 1670
rect 4492 1610 4502 1670
rect 4315 1298 4321 1474
rect 4355 1298 4361 1474
rect 4315 1286 4361 1298
rect 4433 1474 4479 1610
rect 4433 1298 4439 1474
rect 4473 1298 4479 1474
rect 4433 1286 4479 1298
rect 4551 1474 4597 1740
rect 4669 1670 4715 1927
rect 4787 2303 4833 2315
rect 4787 1927 4793 2303
rect 4827 1927 4833 2303
rect 4787 1800 4833 1927
rect 4905 2303 4951 2315
rect 4905 1927 4911 2303
rect 4945 1927 4951 2303
rect 4772 1740 4782 1800
rect 4842 1740 4852 1800
rect 4652 1610 4662 1670
rect 4722 1610 4732 1670
rect 4551 1298 4557 1474
rect 4591 1298 4597 1474
rect 4551 1286 4597 1298
rect 4669 1474 4715 1610
rect 4669 1298 4675 1474
rect 4709 1298 4715 1474
rect 4669 1286 4715 1298
rect 4787 1474 4833 1740
rect 4905 1670 4951 1927
rect 4892 1610 4902 1670
rect 4962 1610 4972 1670
rect 4787 1298 4793 1474
rect 4827 1298 4833 1474
rect 4787 1286 4833 1298
rect 4905 1474 4951 1610
rect 4905 1298 4911 1474
rect 4945 1298 4951 1474
rect 4905 1286 4951 1298
rect 4132 1248 4898 1254
rect 4132 1214 4144 1248
rect 4178 1214 4262 1248
rect 4296 1214 4380 1248
rect 4414 1214 4498 1248
rect 4532 1214 4616 1248
rect 4650 1214 4734 1248
rect 4768 1214 4852 1248
rect 4886 1214 4898 1248
rect 4132 1208 4898 1214
rect 3992 1070 4012 1150
rect 4492 1130 5032 1150
rect 5012 1090 5032 1130
rect 4492 1070 5032 1090
<< via1 >>
rect 4005 2521 4477 2534
rect 4005 2480 4006 2521
rect 4006 2480 4477 2521
rect 4005 2464 4477 2480
rect 4072 1740 4132 1800
rect 4312 1740 4372 1800
rect 4182 1610 4242 1670
rect 4542 1740 4602 1800
rect 4432 1610 4492 1670
rect 4782 1740 4842 1800
rect 4662 1610 4722 1670
rect 4902 1610 4962 1670
rect 4012 1130 4492 1150
rect 4012 1090 4492 1130
rect 4012 1070 4492 1090
<< metal2 >>
rect 3971 2464 4005 2534
rect 4477 2464 4515 2534
rect 4062 1790 4072 1800
rect 4062 1740 4072 1750
rect 4132 1790 4142 1800
rect 4302 1790 4312 1800
rect 4132 1750 4312 1790
rect 4132 1740 4142 1750
rect 4302 1740 4312 1750
rect 4372 1790 4382 1800
rect 4532 1790 4542 1800
rect 4372 1750 4542 1790
rect 4372 1740 4382 1750
rect 4532 1740 4542 1750
rect 4602 1790 4612 1800
rect 4772 1790 4782 1800
rect 4602 1750 4782 1790
rect 4602 1740 4612 1750
rect 4772 1740 4782 1750
rect 4842 1740 4852 1800
rect 4172 1610 4182 1670
rect 4242 1660 4252 1670
rect 4422 1660 4432 1670
rect 4242 1620 4432 1660
rect 4242 1610 4252 1620
rect 4422 1610 4432 1620
rect 4492 1660 4502 1670
rect 4652 1660 4662 1670
rect 4492 1620 4662 1660
rect 4492 1610 4502 1620
rect 4652 1610 4662 1620
rect 4722 1660 4732 1670
rect 4892 1660 4902 1670
rect 4722 1620 4902 1660
rect 4722 1610 4732 1620
rect 4892 1610 4902 1620
rect 4962 1660 4972 1670
rect 4962 1610 4972 1620
rect 3992 1070 4012 1150
rect 4492 1070 4512 1150
<< via2 >>
rect 4005 2469 4477 2529
rect 4012 1080 4492 1140
<< metal3 >>
rect 4662 3440 4902 8540
rect 5122 3430 5362 8530
rect 4052 2534 4172 3130
rect 3971 2529 4515 2534
rect 3971 2469 4005 2529
rect 4477 2469 4515 2529
rect 3971 2464 4515 2469
rect 3992 1140 4512 1150
rect 3992 1080 4012 1140
rect 4492 1080 4512 1140
rect 3992 1070 4512 1080
rect 4022 530 4142 1070
use cmota_1_flat_1  cmota_1_flat_1_0
timestamp 1671334909
transform 1 0 -2776 0 1 3180
box -164 -3800 5363 2800
use sky130_fd_pr__nfet_01v8_NMSMYT  sky130_fd_pr__nfet_01v8_NMSMYT_0
timestamp 1671209795
transform 1 0 3909 0 1 3814
box -551 -310 551 310
use sky130_fd_pr__pfet_01v8_U4PWGH  sky130_fd_pr__pfet_01v8_U4PWGH_0
timestamp 1671209795
transform 1 0 3909 0 1 4593
box -551 -419 551 419
<< end >>
