* NGSPICE file created from unitcell.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2_2 A B VGND VPWR X a_118_74# VNB VPB a_31_74#
X0 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.072e+11p pd=2.04e+06u as=5.217e+11p ps=4.37e+06u w=740000u l=150000u
X1 a_118_74# A a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u w=740000u l=150000u
X2 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 ad=9.96e+11p pd=8.34e+06u as=3.36e+11p ps=2.84e+06u w=1.12e+06u l=150000u
X3 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND B a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR B a_31_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X6 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_31_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 X VGND 0.09fF
C1 VPWR VGND 0.06fF
C2 VPWR X 0.12fF
C3 B VGND 0.01fF
C4 B X 0.00fF
C5 A VGND 0.01fF
C6 A X 0.00fF
C7 B VPWR 0.01fF
C8 VPB VGND 0.02fF
C9 A VPWR 0.04fF
C10 VPB X 0.01fF
C11 A B 0.11fF
C12 VPB VPWR 0.07fF
C13 a_118_74# VGND 0.00fF
C14 VPB B 0.02fF
C15 VPB A 0.02fF
C16 a_118_74# X 0.00fF
C17 a_31_74# VGND 0.12fF
C18 a_31_74# X 0.11fF
C19 a_118_74# VPWR 0.00fF
C20 a_118_74# B 0.00fF
C21 a_31_74# VPWR 0.21fF
C22 a_31_74# B 0.19fF
C23 a_31_74# A 0.03fF
C24 a_31_74# VPB 0.03fF
C25 a_31_74# a_118_74# 0.00fF
C26 VGND VNB 0.34fF
C27 X VNB 0.06fF
C28 VPWR VNB 0.37fF
C29 B VNB 0.09fF
C30 A VNB 0.18fF
C31 VPB VNB 0.62fF
C32 a_31_74# VNB 0.28fF
.ends

.subckt sky130_fd_sc_hs__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=3.24e+06 area=6.417e+11
C0 VPWR VGND 0.02fF
C1 DIODE VGND 0.08fF
C2 DIODE VPWR 0.08fF
C3 VPB VGND 0.01fF
C4 VPB VPWR 0.02fF
C5 VPB DIODE 0.05fF
C6 VGND VNB 0.15fF
C7 VPWR VNB 0.14fF
C8 DIODE VNB 0.24fF
C9 VPB VNB 0.30fF
.ends

.subckt sky130_fd_sc_hs__nand2_2 A B VGND VPWR Y VNB VPB a_27_74#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=1.008e+12p pd=8.52e+06u as=6.72e+11p ps=5.68e+06u w=1.12e+06u l=150000u
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=2.442e+11p pd=2.14e+06u as=6.438e+11p ps=6.18e+06u w=740000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=2.442e+11p pd=2.14e+06u as=0p ps=0u w=740000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
C0 A VPWR 0.01fF
C1 B VPWR 0.01fF
C2 VPB VPWR 0.07fF
C3 B A 0.09fF
C4 VPB A 0.03fF
C5 VPB B 0.03fF
C6 a_27_74# VPWR 0.03fF
C7 a_27_74# A 0.01fF
C8 VGND VPWR 0.05fF
C9 a_27_74# B 0.07fF
C10 a_27_74# VPB 0.01fF
C11 Y VPWR 0.34fF
C12 VGND A 0.01fF
C13 VGND B 0.01fF
C14 Y A 0.12fF
C15 Y B 0.10fF
C16 VGND VPB 0.02fF
C17 Y VPB 0.01fF
C18 VGND a_27_74# 0.24fF
C19 Y a_27_74# 0.13fF
C20 Y VGND 0.01fF
C21 VGND VNB 0.31fF
C22 Y VNB 0.09fF
C23 VPWR VNB 0.36fF
C24 A VNB 0.21fF
C25 B VNB 0.23fF
C26 VPB VNB 0.62fF
C27 a_27_74# VNB 0.09fF
.ends

.subckt cellselect sky130_fd_sc_hs__nand2_2_0/a_27_74# YAND YNAND sky130_fd_sc_hs__and2_2_0/a_118_74#
+ sky130_fd_sc_hs__and2_2_0/a_31_74# S2 S1 VHI VLO
Xsky130_fd_sc_hs__and2_2_0 S2 S1 VLO VHI YAND sky130_fd_sc_hs__and2_2_0/a_118_74#
+ VLO VHI sky130_fd_sc_hs__and2_2_0/a_31_74# sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__diode_2_0 S1 VLO VHI VHI VLO sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__diode_2_1 S2 VLO VHI VHI VLO sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nand2_2_0 S1 S2 VLO VHI YNAND VLO VHI sky130_fd_sc_hs__nand2_2_0/a_27_74#
+ sky130_fd_sc_hs__nand2_2
C0 YAND sky130_fd_sc_hs__and2_2_0/a_31_74# 0.01fF
C1 S1 YNAND 0.07fF
C2 S2 YNAND 0.02fF
C3 S2 S1 1.10fF
C4 sky130_fd_sc_hs__nand2_2_0/a_27_74# YNAND 0.00fF
C5 VHI YNAND 0.03fF
C6 sky130_fd_sc_hs__nand2_2_0/a_27_74# S1 0.01fF
C7 sky130_fd_sc_hs__nand2_2_0/a_27_74# S2 0.00fF
C8 VHI S1 0.25fF
C9 VHI S2 0.36fF
C10 VHI sky130_fd_sc_hs__nand2_2_0/a_27_74# -0.00fF
C11 sky130_fd_sc_hs__and2_2_0/a_118_74# YNAND 0.00fF
C12 sky130_fd_sc_hs__and2_2_0/a_31_74# YNAND 0.00fF
C13 sky130_fd_sc_hs__and2_2_0/a_118_74# S1 0.00fF
C14 sky130_fd_sc_hs__and2_2_0/a_118_74# S2 0.00fF
C15 sky130_fd_sc_hs__and2_2_0/a_31_74# S1 0.02fF
C16 YAND YNAND 0.00fF
C17 sky130_fd_sc_hs__and2_2_0/a_31_74# S2 0.08fF
C18 YAND S1 0.10fF
C19 YAND S2 0.03fF
C20 sky130_fd_sc_hs__and2_2_0/a_118_74# sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.00fF
C21 sky130_fd_sc_hs__and2_2_0/a_118_74# VHI 0.00fF
C22 sky130_fd_sc_hs__and2_2_0/a_31_74# sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.00fF
C23 sky130_fd_sc_hs__and2_2_0/a_31_74# VHI 0.01fF
C24 YAND sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.02fF
C25 YAND VHI 0.03fF
C26 YNAND VLO 0.16fF
C27 S1 VLO 0.88fF
C28 S2 VLO 0.52fF
C29 sky130_fd_sc_hs__nand2_2_0/a_27_74# VLO 0.16fF
C30 VHI VLO 2.98fF
C31 YAND VLO 0.05fF
C32 sky130_fd_sc_hs__and2_2_0/a_118_74# VLO 0.00fF
C33 sky130_fd_sc_hs__and2_2_0/a_31_74# VLO 0.28fF
.ends

.subckt QCS_unit1_flat_dnw G NSUB SD VSUB w_1806_n394# VSUBS
X0 SD G SD VSUB sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
C0 w_1806_n394# VSUB 0.24fF
C1 SD NSUB 0.05fF
C2 G NSUB 0.13fF
C3 G SD 0.12fF
C4 VSUB NSUB 1.34fF
C5 VSUB SD 0.47fF
C6 VSUB G 0.20fF
C7 w_1806_n394# NSUB 5.85fF
C8 w_1806_n394# SD 0.02fF
C9 w_1806_n394# G 0.07fF
C10 SD VSUBS -0.01fF
C11 G VSUBS 0.02fF
C12 VSUB VSUBS 0.10fF
C13 NSUB VSUBS 15.61fF
.ends

.subckt imirror2 OUT a_5468_1540# a_4094_1540# a_4493_207# VLO VHI a_5868_1637# IN
+ a_4036_1637#
X0 VHI a_4493_207# a_4493_207# VHI sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X1 a_4493_207# VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=4.35e+12p ps=3.174e+07u w=5e+06u l=2e+06u
X2 VLO VLO OUT VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X3 a_5868_1637# a_5468_1540# OUT VHI sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X4 OUT OUT VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X5 VLO IN a_4493_207# VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X6 a_4493_207# a_4094_1540# a_4036_1637# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X7 OUT a_4493_207# VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
C0 VHI a_4094_1540# 0.99fF
C1 OUT a_4036_1637# 0.03fF
C2 VHI a_4036_1637# 0.68fF
C3 a_5468_1540# a_4094_1540# 0.00fF
C4 a_5468_1540# a_4036_1637# 0.01fF
C5 IN a_4493_207# 0.46fF
C6 a_5868_1637# a_4493_207# 0.22fF
C7 VHI OUT 1.31fF
C8 a_5468_1540# OUT 0.53fF
C9 a_5468_1540# VHI 0.99fF
C10 a_4094_1540# a_4493_207# 0.44fF
C11 a_4036_1637# a_4493_207# 0.63fF
C12 a_4094_1540# IN 0.17fF
C13 a_4036_1637# IN 0.03fF
C14 a_4094_1540# a_5868_1637# 0.01fF
C15 OUT a_4493_207# 0.88fF
C16 OUT IN 0.22fF
C17 VHI a_4493_207# 3.25fF
C18 a_5468_1540# a_4493_207# 0.22fF
C19 VHI IN 0.19fF
C20 OUT a_5868_1637# 0.47fF
C21 VHI a_5868_1637# 0.45fF
C22 a_5468_1540# a_5868_1637# 0.15fF
C23 a_4036_1637# a_4094_1540# 0.15fF
C24 OUT a_4094_1540# 0.10fF
C25 OUT VLO 3.20fF
C26 VHI VLO 18.78fF
C27 IN VLO 2.36fF
C28 a_5868_1637# VLO 0.34fF
C29 a_4036_1637# VLO 0.34fF
C30 a_5468_1540# VLO 0.34fF
C31 a_4493_207# VLO 1.55fF
C32 a_4094_1540# VLO 0.34fF
.ends

.subckt gated_iref_fix imirror2_0/a_5468_1540# imirror2_0/a_4094_1540# SBAR a_1444_106#
+ imirror2_0/OUT imirror2_0/a_5868_1637# VSUB imirror2_0/VHI imirror2_0/a_4493_207#
+ imirror2_0/a_4036_1637# a_1712_150# S imirror2_0/IN
Ximirror2_0 imirror2_0/OUT imirror2_0/a_5468_1540# imirror2_0/a_4094_1540# imirror2_0/a_4493_207#
+ VSUB imirror2_0/VHI imirror2_0/a_5868_1637# imirror2_0/IN imirror2_0/a_4036_1637#
+ imirror2
X0 imirror2_0/OUT a_1444_106# VSUB sky130_fd_pr__res_xhigh_po w=350000u l=1.49e+06u
X1 VSUB SBAR a_1712_150# VSUB sky130_fd_pr__nfet_01v8 ad=5.95e+12p pd=4.302e+07u as=1.65e+12p ps=1.132e+07u w=2.5e+06u l=150000u
X2 VSUB a_1712_150# sky130_fd_pr__cap_mim_m3_1 l=6.2e+06u w=2.76e+07u
X3 a_1712_150# VSUB sky130_fd_pr__cap_mim_m3_2 l=6.2e+06u w=2.76e+07u
X4 a_1712_150# S a_1444_106# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.6e+12p ps=1.128e+07u w=2.5e+06u l=150000u
X5 VSUB VSUB a_1444_106# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X6 a_1712_150# SBAR VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X7 a_1444_106# S a_1712_150# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
C0 imirror2_0/IN imirror2_0/a_4493_207# 0.12fF
C1 a_1712_150# imirror2_0/a_4493_207# 0.29fF
C2 imirror2_0/IN imirror2_0/VHI 0.00fF
C3 imirror2_0/OUT imirror2_0/a_4493_207# 0.00fF
C4 imirror2_0/VHI a_1712_150# 0.88fF
C5 imirror2_0/IN a_1712_150# 0.12fF
C6 imirror2_0/IN a_1444_106# 0.00fF
C7 imirror2_0/IN SBAR 0.01fF
C8 imirror2_0/IN S 0.01fF
C9 imirror2_0/VHI imirror2_0/OUT 0.03fF
C10 imirror2_0/IN imirror2_0/OUT 0.07fF
C11 a_1444_106# a_1712_150# 0.93fF
C12 SBAR a_1712_150# 0.25fF
C13 SBAR a_1444_106# 0.07fF
C14 S a_1712_150# 0.27fF
C15 S a_1444_106# 0.03fF
C16 S SBAR 0.71fF
C17 imirror2_0/OUT a_1712_150# 1.57fF
C18 imirror2_0/OUT a_1444_106# 0.33fF
C19 imirror2_0/OUT SBAR 0.14fF
C20 imirror2_0/OUT S 0.13fF
C21 a_1712_150# imirror2_0/a_5868_1637# 0.33fF
C22 a_1712_150# imirror2_0/a_5468_1540# 0.33fF
C23 imirror2_0/OUT imirror2_0/a_5868_1637# 0.00fF
C24 imirror2_0/OUT imirror2_0/a_5468_1540# 0.00fF
C25 a_1712_150# VSUB 39.40fF
C26 a_1444_106# VSUB 1.29fF
C27 SBAR VSUB 0.76fF
C28 S VSUB 0.77fF
C29 imirror2_0/OUT VSUB 4.89fF
C30 imirror2_0/VHI VSUB 19.26fF
C31 imirror2_0/IN VSUB 4.59fF
C32 imirror2_0/a_5868_1637# VSUB 0.44fF
C33 imirror2_0/a_4036_1637# VSUB 0.34fF
C34 imirror2_0/a_5468_1540# VSUB 0.49fF
C35 imirror2_0/a_4493_207# VSUB 1.64fF
C36 imirror2_0/a_4094_1540# VSUB 0.34fF
.ends

.subckt sky130_fd_pr__res_high_po_0p69_G8QCSG a_48_n518# a_n186_n518# a_n316_n648#
X0 a_n186_n518# a_48_n518# a_n316_n648# sky130_fd_pr__res_high_po w=690000u l=5.83e+06u
C0 a_n186_n518# a_48_n518# 0.18fF
C1 a_48_n518# a_n316_n648# 0.52fF
C2 a_n186_n518# a_n316_n648# 0.52fF
.ends

.subckt cmota_gb_rp VREF COM VIP VIN DP li_5300_n960# VLO a_2217_285# DN VOP VHI a_2925_285#
+ VMN
Xsky130_fd_pr__res_high_po_0p69_G8QCSG_0 li_5300_n960# VMN VLO sky130_fd_pr__res_high_po_0p69_G8QCSG
X0 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=4.93e+13p pd=3.4986e+08u as=1.16e+13p ps=8.232e+07u w=1e+07u l=300000u
X1 VHI DN DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.174e+07u w=1e+07u l=300000u
X2 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+13p ps=8.232e+07u w=1e+07u l=300000u
X3 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.264e+07u as=1.3225e+13p ps=9.21e+07u w=2.5e+06u l=150000u
X4 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X5 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.264e+07u as=0p ps=0u w=2.5e+06u l=150000u
X6 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X7 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X8 VHI VHI VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X9 a_2925_285# DN VHI VHI sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=300000u
X10 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X11 li_5300_n960# VOP sky130_fd_pr__cap_mim_m3_2 l=1.32e+07u w=3.7e+06u
X12 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X13 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X14 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X15 COM VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.8e+13p ps=2.69525e+08u w=2.5e+06u l=150000u
X16 VLO VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.116e+07u w=1e+07u l=300000u
X17 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X18 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X19 VHI DN DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.174e+07u w=1e+07u l=300000u
X20 VHI DP DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X21 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X22 VLO VREF COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X23 VMN VHI VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X24 DN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X25 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X26 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X27 VLO VREF COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X28 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X29 DN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X30 DP DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X31 DN DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X32 DP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X33 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X34 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X35 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X36 VHI DN DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X37 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X38 VMN VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=5.8e+12p pd=4.116e+07u as=0p ps=0u w=1e+07u l=300000u
X39 VLO VMN VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X40 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X41 VOP VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X42 VHI DP DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X43 VLO VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X44 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X45 VLO VLO COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X46 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X47 VHI DP a_2217_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=300000u
X48 VHI DP DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X49 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X50 COM VREF VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X51 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X52 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X53 COM VREF VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X54 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X55 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X56 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X57 DP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X58 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X59 a_2217_285# DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X60 VMN VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X61 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X62 VLO VMN VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X63 VOP VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X64 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X65 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X66 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X67 VOP li_5300_n960# sky130_fd_pr__cap_mim_m3_1 l=1.32e+07u w=3.7e+06u
X68 VHI DN a_2925_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X69 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
C0 VIP COM 0.71fF
C1 VIN COM 0.71fF
C2 VIN VIP 0.11fF
C3 VOP COM 0.05fF
C4 VOP VIP 0.01fF
C5 a_2925_285# COM 0.01fF
C6 a_2925_285# VIP 0.00fF
C7 a_2925_285# VOP 0.05fF
C8 COM VREF 2.35fF
C9 VIP VREF 0.36fF
C10 VIN VREF 0.36fF
C11 COM VMN 0.33fF
C12 VOP VREF 0.03fF
C13 a_2925_285# VREF 0.00fF
C14 VIP VMN 0.14fF
C15 VIN VMN 0.15fF
C16 COM DN 6.05fF
C17 VOP li_5300_n960# 9.33fF
C18 VIP DN 0.05fF
C19 VOP VMN 0.72fF
C20 a_2925_285# VMN 0.01fF
C21 VIN DN 0.53fF
C22 COM a_2217_285# 0.01fF
C23 VOP DN 0.06fF
C24 a_2925_285# DN 0.13fF
C25 COM VHI 0.10fF
C26 VIN a_2217_285# 0.00fF
C27 VIP VHI 0.10fF
C28 COM DP 6.02fF
C29 VOP a_2217_285# 0.01fF
C30 a_2925_285# a_2217_285# 0.02fF
C31 VIP DP 0.53fF
C32 VIN VHI 0.11fF
C33 VOP VHI 18.23fF
C34 VIN DP 0.04fF
C35 a_2925_285# VHI 4.31fF
C36 VOP DP 0.97fF
C37 VMN VREF 0.10fF
C38 a_2925_285# DP 0.17fF
C39 DN VREF 0.14fF
C40 VMN li_5300_n960# 1.12fF
C41 a_2217_285# VREF 0.00fF
C42 DN VMN 1.12fF
C43 VHI VREF 0.04fF
C44 a_2217_285# VMN 0.06fF
C45 DP VREF 0.14fF
C46 VHI li_5300_n960# 2.02fF
C47 a_2217_285# DN 0.17fF
C48 VHI VMN 17.75fF
C49 DP li_5300_n960# 0.48fF
C50 DP VMN 0.34fF
C51 VHI DN 16.22fF
C52 DP DN 1.21fF
C53 VHI a_2217_285# 4.31fF
C54 DP a_2217_285# 0.13fF
C55 DP VHI 16.22fF
C56 VREF VLO 7.20fF
C57 COM VLO 6.11fF
C58 VIP VLO 0.78fF
C59 VIN VLO 0.79fF
C60 VOP VLO 9.34fF
C61 a_2925_285# VLO -0.04fF
C62 a_2217_285# VLO -0.04fF
C63 DP VLO 1.36fF
C64 DN VLO 1.42fF
C65 VHI VLO 35.14fF
C66 li_5300_n960# VLO 3.02fF
C67 VMN VLO 13.45fF
.ends

.subckt cmota_gb_rp_gp cmota_gb_rp_0/DP cmota_gb_rp_0/DN cmota_gb_rp_0/COM gated_iref_fix_0/imirror2_0/a_4094_1540#
+ gated_iref_fix_0/imirror2_0/a_5468_1540# VREF gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_0/VMN
+ gated_iref_fix_0/imirror2_0/a_5868_1637# VIP cmota_gb_rp_0/li_5300_n960# SBAR VIN
+ gated_iref_fix_0/imirror2_0/a_4036_1637# S VOP VHI gated_iref_fix_0/a_1444_106#
+ cmota_gb_rp_0/a_2217_285# gated_iref_fix_0/imirror2_0/a_4493_207# VREF_GATED cmota_gb_rp_0/a_2925_285#
+ VLO
Xgated_iref_fix_0 gated_iref_fix_0/imirror2_0/a_5468_1540# gated_iref_fix_0/imirror2_0/a_4094_1540#
+ SBAR gated_iref_fix_0/a_1444_106# gated_iref_fix_0/imirror2_0/OUT gated_iref_fix_0/imirror2_0/a_5868_1637#
+ VLO VHI gated_iref_fix_0/imirror2_0/a_4493_207# gated_iref_fix_0/imirror2_0/a_4036_1637#
+ VREF_GATED S VREF gated_iref_fix
Xcmota_gb_rp_0 VREF_GATED cmota_gb_rp_0/COM VIP VIN cmota_gb_rp_0/DP cmota_gb_rp_0/li_5300_n960#
+ VLO cmota_gb_rp_0/a_2217_285# cmota_gb_rp_0/DN VOP VHI cmota_gb_rp_0/a_2925_285#
+ cmota_gb_rp_0/VMN cmota_gb_rp
X0 VLO VHI sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=1.3e+07u
X1 VHI VLO sky130_fd_pr__cap_mim_m3_1 l=3.1e+07u w=1.3e+07u
C0 SBAR gated_iref_fix_0/a_1444_106# 0.00fF
C1 S SBAR 0.10fF
C2 VREF gated_iref_fix_0/a_1444_106# 0.00fF
C3 gated_iref_fix_0/imirror2_0/a_5468_1540# VREF_GATED -0.31fF
C4 gated_iref_fix_0/imirror2_0/a_4493_207# VREF_GATED -0.29fF
C5 VREF SBAR 0.02fF
C6 VREF S 0.03fF
C7 gated_iref_fix_0/imirror2_0/a_5468_1540# VHI 0.00fF
C8 gated_iref_fix_0/imirror2_0/a_4493_207# VHI 0.19fF
C9 cmota_gb_rp_0/VMN VREF_GATED 1.54fF
C10 cmota_gb_rp_0/VMN cmota_gb_rp_0/COM -0.00fF
C11 gated_iref_fix_0/imirror2_0/a_4094_1540# VHI 0.01fF
C12 VREF_GATED gated_iref_fix_0/a_1444_106# 0.00fF
C13 cmota_gb_rp_0/VMN VIN -0.00fF
C14 cmota_gb_rp_0/VMN VHI 0.15fF
C15 VREF_GATED SBAR 0.02fF
C16 cmota_gb_rp_0/VMN VOP 0.00fF
C17 VHI gated_iref_fix_0/a_1444_106# 0.00fF
C18 VREF_GATED S 0.00fF
C19 gated_iref_fix_0/imirror2_0/OUT SBAR 0.00fF
C20 VHI cmota_gb_rp_0/li_5300_n960# 0.03fF
C21 cmota_gb_rp_0/li_5300_n960# VOP 0.00fF
C22 gated_iref_fix_0/imirror2_0/OUT S 0.00fF
C23 VHI SBAR 0.00fF
C24 VHI S 0.00fF
C25 VREF_GATED VREF -0.04fF
C26 gated_iref_fix_0/imirror2_0/OUT VREF 0.00fF
C27 VHI gated_iref_fix_0/imirror2_0/a_4036_1637# 0.07fF
C28 VHI VREF 0.16fF
C29 VREF_GATED cmota_gb_rp_0/COM 0.17fF
C30 gated_iref_fix_0/imirror2_0/a_5868_1637# VREF_GATED -0.07fF
C31 gated_iref_fix_0/imirror2_0/OUT VREF_GATED -0.37fF
C32 VREF_GATED VIN 0.00fF
C33 VHI VREF_GATED 3.68fF
C34 VIN cmota_gb_rp_0/COM -0.00fF
C35 VHI gated_iref_fix_0/imirror2_0/a_5868_1637# 0.03fF
C36 VIN VIP 0.00fF
C37 VHI gated_iref_fix_0/imirror2_0/OUT 0.17fF
C38 VHI VOP 0.11fF
C39 VHI cmota_gb_rp_0/a_2925_285# 0.04fF
C40 VREF_GATED cmota_gb_rp_0/DN 0.40fF
C41 VHI cmota_gb_rp_0/a_2217_285# 0.04fF
C42 VHI cmota_gb_rp_0/DP 0.81fF
C43 cmota_gb_rp_0/DP VOP -0.00fF
C44 VHI cmota_gb_rp_0/DN 0.89fF
C45 cmota_gb_rp_0/COM VLO 6.15fF
C46 VIP VLO 0.78fF
C47 VIN VLO 0.79fF
C48 VOP VLO 9.31fF
C49 cmota_gb_rp_0/a_2925_285# VLO -0.04fF
C50 cmota_gb_rp_0/a_2217_285# VLO -0.04fF
C51 cmota_gb_rp_0/DP VLO 1.36fF
C52 cmota_gb_rp_0/DN VLO 1.55fF
C53 cmota_gb_rp_0/li_5300_n960# VLO 2.88fF
C54 cmota_gb_rp_0/VMN VLO 14.06fF
C55 VREF_GATED VLO 52.16fF
C56 gated_iref_fix_0/a_1444_106# VLO 1.29fF
C57 SBAR VLO 0.76fF
C58 S VLO 0.78fF
C59 gated_iref_fix_0/imirror2_0/OUT VLO 6.43fF
C60 VHI VLO 134.20fF
C61 VREF VLO 6.75fF
C62 gated_iref_fix_0/imirror2_0/a_5868_1637# VLO 0.48fF
C63 gated_iref_fix_0/imirror2_0/a_4036_1637# VLO 0.88fF
C64 gated_iref_fix_0/imirror2_0/a_5468_1540# VLO 0.63fF
C65 gated_iref_fix_0/imirror2_0/a_4493_207# VLO 4.55fF
C66 gated_iref_fix_0/imirror2_0/a_4094_1540# VLO 0.94fF
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_EP3CBP a_48_n582# a_n118_150# a_n118_n582#
+ a_48_150# a_n248_n712#
X0 a_48_n582# a_48_150# a_n248_n712# sky130_fd_pr__res_xhigh_po_0p35 l=1.5e+06u
X1 a_n118_n582# a_n118_150# a_n248_n712# sky130_fd_pr__res_xhigh_po_0p35 l=1.5e+06u
C0 a_48_n582# a_48_150# 0.02fF
C1 a_48_n582# a_n118_n582# 0.29fF
C2 a_n118_150# a_48_150# 0.29fF
C3 a_n118_150# a_n118_n582# 0.02fF
C4 a_48_n582# a_n248_n712# 0.47fF
C5 a_48_150# a_n248_n712# 0.47fF
C6 a_n118_n582# a_n248_n712# 0.51fF
C7 a_n118_150# a_n248_n712# 0.51fF
.ends

.subckt unitcell VMID VSD VHI VTW ROWSEL VREF A B COLSEL VMID_1 VSD_1 QCS_GATE VLO
Xcellselect_0 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# cellselect_0/YAND cellselect_0/YNAND
+ cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74#
+ COLSEL ROWSEL VHI VLO cellselect
Xcellselect_1 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# cellselect_1/YAND cellselect_1/YNAND
+ cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74#
+ COLSEL ROWSEL VHI VLO cellselect
XQCS_unit1_flat_dnw_0 QCS_GATE VHI VSD_1 A w_20886_n3514# VLO QCS_unit1_flat_dnw
Xcmota_gb_rp_gp_1 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP cmota_gb_rp_gp_1/cmota_gb_rp_0/DN
+ cmota_gb_rp_gp_1/cmota_gb_rp_0/COM cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4094_1540#
+ cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# VREF cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT
+ cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637#
+ cmota_gb_rp_gp_1/VIP cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# cellselect_1/YNAND
+ cmota_gb_rp_gp_1/VIN cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4036_1637# cellselect_1/YAND
+ QCS_GATE VHI cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2217_285#
+ cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_1/VREF_GATED
+ cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2925_285# VLO cmota_gb_rp_gp
Xcmota_gb_rp_gp_2 cmota_gb_rp_gp_2/cmota_gb_rp_0/DP cmota_gb_rp_gp_2/cmota_gb_rp_0/DN
+ cmota_gb_rp_gp_2/cmota_gb_rp_0/COM cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4094_1540#
+ cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# VREF cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT
+ cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637#
+ VMID_1 cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# cellselect_0/YNAND A cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4036_1637#
+ cellselect_0/YAND B VHI cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2217_285#
+ cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_2/VREF_GATED
+ cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2925_285# VLO cmota_gb_rp_gp
Xsky130_fd_pr__res_xhigh_po_0p35_EP3CBP_0 QCS_GATE cmota_gb_rp_gp_1/VIN QCS_GATE VMID_1
+ VLO sky130_fd_pr__res_xhigh_po_0p35_EP3CBP
X0 VLO VMID_1 sky130_fd_pr__cap_mim_m3_1 l=1.16e+07u w=7.8e+06u
X1 VLO VMID_1 sky130_fd_pr__cap_mim_m3_1 l=4.6e+06u w=6.5e+06u
X2 VHI VMID_1 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.8e+06u
X3 VSD VSD_1 VLO sky130_fd_pr__res_xhigh_po_0p35 l=2e+06u
X4 VMID_1 VLO sky130_fd_pr__cap_mim_m3_2 l=4.6e+06u w=6.5e+06u
X5 VLO VSD_1 sky130_fd_pr__cap_mim_m3_1 l=1.01e+07u w=7.8e+06u
X6 VMID VMID_1 VLO sky130_fd_pr__res_xhigh_po_0p35 l=2e+06u
X7 VMID_1 VHI sky130_fd_pr__cap_mim_m3_2 l=1.77e+07u w=2.2e+06u
C0 VREF VMID_1 0.61fF
C1 VSD_1 VMID 0.06fF
C2 cellselect_1/YAND cmota_gb_rp_gp_1/VREF_GATED 0.03fF
C3 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# ROWSEL 0.00fF
C4 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# VMID_1 1.95fF
C5 cmota_gb_rp_gp_2/VREF_GATED cmota_gb_rp_gp_2/cmota_gb_rp_0/COM -0.00fF
C6 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# COLSEL 0.01fF
C7 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# -0.00fF
C8 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# -0.00fF
C9 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_2/VREF_GATED -0.10fF
C10 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# VREF 0.01fF
C11 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# cmota_gb_rp_gp_1/VREF_GATED -0.01fF
C12 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# 0.13fF
C13 VHI cmota_gb_rp_gp_1/VREF_GATED 0.05fF
C14 VHI cmota_gb_rp_gp_2/cmota_gb_rp_0/DP 0.00fF
C15 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_1/VREF_GATED 0.01fF
C16 VMID VSD 15.30fF
C17 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# -0.00fF
C18 ROWSEL cmota_gb_rp_gp_1/VREF_GATED 0.04fF
C19 cmota_gb_rp_gp_2/VREF_GATED B 0.00fF
C20 cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# VMID_1 1.14fF
C21 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN VHI 0.02fF
C22 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cellselect_0/YNAND 0.01fF
C23 COLSEL cmota_gb_rp_gp_1/VREF_GATED 2.49fF
C24 cmota_gb_rp_gp_1/VREF_GATED cmota_gb_rp_gp_1/VIN 0.02fF
C25 VREF cmota_gb_rp_gp_1/VREF_GATED 0.10fF
C26 VMID_1 VTW 0.49fF
C27 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# 0.11fF
C28 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN COLSEL 0.01fF
C29 w_20886_n3514# VMID_1 0.44fF
C30 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/VIN 0.33fF
C31 ROWSEL VMID 8.06fF
C32 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C33 VHI cmota_gb_rp_gp_1/VIP -0.02fF
C34 COLSEL VMID 0.29fF
C35 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# -0.08fF
C36 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# -0.03fF
C37 VREF VMID 4.69fF
C38 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# cmota_gb_rp_gp_1/VREF_GATED 0.01fF
C39 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_1/VREF_GATED -0.00fF
C40 QCS_GATE cmota_gb_rp_gp_1/cmota_gb_rp_0/COM 0.00fF
C41 cmota_gb_rp_gp_1/VIN cmota_gb_rp_gp_1/VIP 0.32fF
C42 A cmota_gb_rp_gp_2/cmota_gb_rp_0/COM 0.50fF
C43 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN cmota_gb_rp_gp_2/cmota_gb_rp_0/COM 0.02fF
C44 cellselect_0/YAND cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.00fF
C45 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# cmota_gb_rp_gp_1/VREF_GATED 0.00fF
C46 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.02fF
C47 cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2925_285# cmota_gb_rp_gp_1/VIN 0.00fF
C48 cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2925_285# VMID_1 0.00fF
C49 B A 2.20fF
C50 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C51 cellselect_1/YAND cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT -0.01fF
C52 ROWSEL cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.00fF
C53 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN w_20886_n3514# 0.00fF
C54 VHI cmota_gb_rp_gp_1/cmota_gb_rp_0/DP 0.01fF
C55 cellselect_1/YAND cellselect_1/YNAND 0.05fF
C56 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.01fF
C57 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# cmota_gb_rp_gp_1/VREF_GATED -0.03fF
C58 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# -0.00fF
C59 VHI cmota_gb_rp_gp_1/cmota_gb_rp_0/DN 0.00fF
C60 VREF cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.01fF
C61 VMID VTW 2.37fF
C62 cellselect_1/YNAND cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.00fF
C63 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT -0.09fF
C64 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4094_1540# 0.00fF
C65 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP cmota_gb_rp_gp_1/VIN 0.06fF
C66 cmota_gb_rp_gp_2/cmota_gb_rp_0/DP VMID_1 0.03fF
C67 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT VHI -0.11fF
C68 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C69 cmota_gb_rp_gp_1/cmota_gb_rp_0/DN cmota_gb_rp_gp_1/VIN 0.01fF
C70 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN VMID_1 0.06fF
C71 cellselect_1/YNAND VHI 0.03fF
C72 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT ROWSEL 0.01fF
C73 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# cellselect_1/YNAND 0.00fF
C74 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cellselect_0/YAND -0.00fF
C75 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4094_1540# 0.00fF
C76 cellselect_1/YNAND ROWSEL 0.00fF
C77 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT COLSEL 0.84fF
C78 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT -0.11fF
C79 VREF cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C80 VMID_1 VMID 0.63fF
C81 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4036_1637# 0.00fF
C82 cellselect_1/YNAND COLSEL 0.17fF
C83 ROWSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.01fF
C84 cellselect_0/YNAND cmota_gb_rp_gp_2/VREF_GATED 0.05fF
C85 VREF cellselect_1/YNAND 0.04fF
C86 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.88fF
C87 VREF cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C88 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# -0.00fF
C89 VHI B 4.50fF
C90 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# cmota_gb_rp_gp_2/VREF_GATED 0.01fF
C91 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.00fF
C92 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT -0.00fF
C93 cellselect_1/YNAND cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# -0.00fF
C94 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# cmota_gb_rp_gp_2/VREF_GATED -0.03fF
C95 COLSEL B 4.52fF
C96 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/VREF_GATED -0.00fF
C97 QCS_GATE A 0.17fF
C98 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# 0.00fF
C99 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# B 0.03fF
C100 VSD_1 QCS_GATE 0.19fF
C101 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# cellselect_0/YNAND -0.00fF
C102 cmota_gb_rp_gp_2/VREF_GATED A 0.78fF
C103 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN cmota_gb_rp_gp_2/VREF_GATED 0.01fF
C104 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP VMID_1 0.00fF
C105 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/VIP -0.06fF
C106 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.00fF
C107 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT -0.03fF
C108 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# cmota_gb_rp_gp_2/VREF_GATED 0.00fF
C109 cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# B 0.13fF
C110 cmota_gb_rp_gp_1/VIN cmota_gb_rp_gp_1/cmota_gb_rp_0/COM 0.10fF
C111 VMID_1 cmota_gb_rp_gp_2/cmota_gb_rp_0/COM 0.29fF
C112 VHI QCS_GATE 1.86fF
C113 cellselect_0/YAND cmota_gb_rp_gp_2/VREF_GATED 0.03fF
C114 VHI cmota_gb_rp_gp_2/VREF_GATED 0.03fF
C115 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT 0.00fF
C116 cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2925_285# cmota_gb_rp_gp_1/VIP -0.00fF
C117 QCS_GATE cmota_gb_rp_gp_1/VIN 0.26fF
C118 B VMID_1 0.80fF
C119 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/cmota_gb_rp_0/DP -0.00fF
C120 ROWSEL cmota_gb_rp_gp_2/VREF_GATED 0.04fF
C121 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN A 0.33fF
C122 COLSEL cmota_gb_rp_gp_2/VREF_GATED 2.76fF
C123 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# QCS_GATE 0.76fF
C124 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_1/VREF_GATED -0.14fF
C125 VSD_1 A 0.27fF
C126 cellselect_0/YAND cellselect_0/YNAND 0.07fF
C127 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# -0.00fF
C128 VREF cmota_gb_rp_gp_2/VREF_GATED 0.10fF
C129 cellselect_1/YNAND cmota_gb_rp_gp_1/VREF_GATED 0.05fF
C130 VHI cellselect_0/YNAND 0.02fF
C131 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP cmota_gb_rp_gp_1/VIP -0.09fF
C132 cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2217_285# A 0.00fF
C133 ROWSEL cellselect_0/YNAND 0.00fF
C134 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# cellselect_0/YAND 0.02fF
C135 cmota_gb_rp_gp_1/cmota_gb_rp_0/DN cmota_gb_rp_gp_1/VIP -0.01fF
C136 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# -0.09fF
C137 COLSEL cellselect_0/YNAND 0.14fF
C138 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# VHI 0.00fF
C139 QCS_GATE cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# 0.02fF
C140 VREF cellselect_0/YNAND 0.04fF
C141 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# ROWSEL 0.00fF
C142 VHI cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# -0.01fF
C143 cmota_gb_rp_gp_2/cmota_gb_rp_0/DN A 0.04fF
C144 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# COLSEL 0.01fF
C145 w_20886_n3514# QCS_GATE 0.24fF
C146 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# VREF 0.01fF
C147 VSD_1 VSD 0.49fF
C148 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN cmota_gb_rp_gp_2/cmota_gb_rp_0/DN 0.00fF
C149 COLSEL cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# 0.22fF
C150 VHI cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4036_1637# 0.00fF
C151 VHI A 6.64fF
C152 VHI cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN 0.02fF
C153 VHI VSD_1 1.59fF
C154 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# cellselect_0/YAND 0.00fF
C155 COLSEL A 6.71fF
C156 cmota_gb_rp_gp_1/VIN A 0.00fF
C157 QCS_GATE VMID_1 1.30fF
C158 ROWSEL VSD_1 0.05fF
C159 VHI cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4094_1540# 0.00fF
C160 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# VHI 0.00fF
C161 COLSEL cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN 0.01fF
C162 cellselect_1/YAND cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.00fF
C163 cmota_gb_rp_gp_1/VIN cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN 0.00fF
C164 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# ROWSEL 0.00fF
C165 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# A 0.02fF
C166 VREF VSD_1 0.13fF
C167 cmota_gb_rp_gp_2/VREF_GATED VMID_1 0.87fF
C168 COLSEL cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4094_1540# 0.00fF
C169 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# COLSEL 0.00fF
C170 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# -0.00fF
C171 cellselect_1/YAND VHI 0.04fF
C172 VREF cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# 0.00fF
C173 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# cellselect_1/YAND 0.01fF
C174 cellselect_1/YAND ROWSEL 0.25fF
C175 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN cmota_gb_rp_gp_1/cmota_gb_rp_0/COM -0.00fF
C176 VHI cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.03fF
C177 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_2/VREF_GATED 0.01fF
C178 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.00fF
C179 ROWSEL VSD 2.52fF
C180 cellselect_1/YAND COLSEL 0.63fF
C181 VHI cellselect_0/YAND 0.03fF
C182 ROWSEL cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.00fF
C183 cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# A 1.53fF
C184 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT cellselect_1/YNAND 0.01fF
C185 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# VHI -0.00fF
C186 cellselect_1/YAND VREF 0.09fF
C187 COLSEL VSD 0.17fF
C188 ROWSEL cellselect_0/YAND 0.17fF
C189 COLSEL cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.01fF
C190 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_2/VREF_GATED -0.00fF
C191 VREF VSD 4.80fF
C192 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# VHI 0.02fF
C193 VREF cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# 0.01fF
C194 COLSEL cellselect_0/YAND 0.64fF
C195 ROWSEL VHI 0.90fF
C196 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# COLSEL 0.11fF
C197 cmota_gb_rp_gp_1/VIP cmota_gb_rp_gp_1/cmota_gb_rp_0/COM -0.05fF
C198 w_20886_n3514# A 0.21fF
C199 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# ROWSEL 0.00fF
C200 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN QCS_GATE 0.32fF
C201 VREF cellselect_0/YAND 0.10fF
C202 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# cellselect_0/YNAND 0.00fF
C203 COLSEL VHI 11.34fF
C204 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# COLSEL 0.01fF
C205 VHI cmota_gb_rp_gp_1/VIN 0.05fF
C206 w_20886_n3514# cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN 0.00fF
C207 VSD_1 VTW 0.57fF
C208 VREF VHI 0.91fF
C209 cellselect_1/YAND cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.02fF
C210 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# VREF 0.01fF
C211 w_20886_n3514# VSD_1 0.31fF
C212 COLSEL ROWSEL 2.68fF
C213 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# cmota_gb_rp_gp_2/VREF_GATED -0.01fF
C214 VREF ROWSEL 8.01fF
C215 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# VHI 0.91fF
C216 VREF COLSEL 1.05fF
C217 QCS_GATE cmota_gb_rp_gp_1/VIP 0.00fF
C218 A VMID_1 1.63fF
C219 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# -0.00fF
C220 cellselect_1/YAND cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# 0.00fF
C221 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# VHI 0.01fF
C222 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN VMID_1 0.16fF
C223 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# VHI -0.01fF
C224 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# cmota_gb_rp_gp_1/VIN 0.26fF
C225 VSD_1 VMID_1 2.31fF
C226 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# ROWSEL 0.00fF
C227 VSD VTW 4.61fF
C228 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# -0.00fF
C229 VHI cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# 0.87fF
C230 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# COLSEL 0.02fF
C231 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# COLSEL 0.13fF
C232 cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2925_285# A 0.00fF
C233 VREF cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# 0.01fF
C234 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# VHI 0.00fF
C235 VHI VTW 0.14fF
C236 w_20886_n3514# VHI 0.34fF
C237 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# ROWSEL 0.00fF
C238 cmota_gb_rp_gp_1/VIN cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# 0.02fF
C239 ROWSEL VTW 0.47fF
C240 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# COLSEL 0.00fF
C241 VMID_1 VSD 0.39fF
C242 COLSEL VTW 0.33fF
C243 VREF cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# 0.00fF
C244 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP QCS_GATE 0.01fF
C245 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# 0.02fF
C246 cmota_gb_rp_gp_2/cmota_gb_rp_0/DN VMID_1 0.00fF
C247 cmota_gb_rp_gp_2/cmota_gb_rp_0/DP A 0.12fF
C248 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# VHI -0.01fF
C249 VREF VTW 7.49fF
C250 w_20886_n3514# cmota_gb_rp_gp_1/VIN 0.01fF
C251 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN A 0.00fF
C252 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN cmota_gb_rp_gp_2/cmota_gb_rp_0/DP 0.02fF
C253 VHI VMID_1 10.40fF
C254 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# COLSEL 0.25fF
C255 ROWSEL VMID_1 0.24fF
C256 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# cellselect_0/YAND 0.01fF
C257 cellselect_0/YNAND cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# 0.00fF
C258 cmota_gb_rp_gp_1/VIN VMID_1 0.24fF
C259 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# VHI 0.01fF
C260 VTW VLO 17.46fF
C261 VSD VLO 24.39fF
C262 VMID VLO 13.04fF
C263 cmota_gb_rp_gp_2/cmota_gb_rp_0/COM VLO 6.14fF
C264 VMID_1 VLO 28.79fF
C265 A VLO 71.20fF
C266 B VLO 77.54fF
C267 cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2925_285# VLO -0.04fF
C268 cmota_gb_rp_gp_2/cmota_gb_rp_0/a_2217_285# VLO -0.04fF
C269 cmota_gb_rp_gp_2/cmota_gb_rp_0/DP VLO 1.36fF
C270 cmota_gb_rp_gp_2/cmota_gb_rp_0/DN VLO 1.42fF
C271 cmota_gb_rp_gp_2/cmota_gb_rp_0/li_5300_n960# VLO 2.89fF
C272 cmota_gb_rp_gp_2/cmota_gb_rp_0/VMN VLO 13.49fF
C273 cmota_gb_rp_gp_2/VREF_GATED VLO 44.14fF
C274 cmota_gb_rp_gp_2/gated_iref_fix_0/a_1444_106# VLO 1.22fF
C275 cellselect_0/YNAND VLO 0.90fF
C276 cellselect_0/YAND VLO 1.04fF
C277 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/OUT VLO 4.23fF
C278 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5868_1637# VLO 0.34fF
C279 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4036_1637# VLO 0.34fF
C280 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_5468_1540# VLO 0.34fF
C281 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4493_207# VLO 1.55fF
C282 cmota_gb_rp_gp_2/gated_iref_fix_0/imirror2_0/a_4094_1540# VLO 0.34fF
C283 cmota_gb_rp_gp_1/cmota_gb_rp_0/COM VLO 6.11fF
C284 cmota_gb_rp_gp_1/VIP VLO 0.78fF
C285 cmota_gb_rp_gp_1/VIN VLO 2.40fF
C286 QCS_GATE VLO 11.22fF
C287 cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2925_285# VLO -0.04fF
C288 cmota_gb_rp_gp_1/cmota_gb_rp_0/a_2217_285# VLO -0.04fF
C289 cmota_gb_rp_gp_1/cmota_gb_rp_0/DP VLO 1.36fF
C290 cmota_gb_rp_gp_1/cmota_gb_rp_0/DN VLO 1.42fF
C291 cmota_gb_rp_gp_1/cmota_gb_rp_0/li_5300_n960# VLO 2.89fF
C292 cmota_gb_rp_gp_1/cmota_gb_rp_0/VMN VLO 13.26fF
C293 cmota_gb_rp_gp_1/VREF_GATED VLO 44.11fF
C294 cmota_gb_rp_gp_1/gated_iref_fix_0/a_1444_106# VLO 1.22fF
C295 cellselect_1/YNAND VLO 0.88fF
C296 cellselect_1/YAND VLO 0.95fF
C297 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/OUT VLO 4.22fF
C298 VHI VLO 284.28fF
C299 VREF VLO 25.59fF
C300 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5868_1637# VLO 0.34fF
C301 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4036_1637# VLO 0.34fF
C302 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_5468_1540# VLO 0.34fF
C303 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4493_207# VLO 1.55fF
C304 cmota_gb_rp_gp_1/gated_iref_fix_0/imirror2_0/a_4094_1540# VLO 0.34fF
C305 VSD_1 VLO 12.49fF
C306 w_20886_n3514# VLO 0.20fF
C307 ROWSEL VLO 21.24fF
C308 COLSEL VLO 35.41fF
C309 cellselect_1/sky130_fd_sc_hs__nand2_2_0/a_27_74# VLO 0.12fF
C310 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_118_74# VLO 0.00fF
C311 cellselect_1/sky130_fd_sc_hs__and2_2_0/a_31_74# VLO 0.32fF
C312 cellselect_0/sky130_fd_sc_hs__nand2_2_0/a_27_74# VLO 0.12fF
C313 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_118_74# VLO 0.00fF
C314 cellselect_0/sky130_fd_sc_hs__and2_2_0/a_31_74# VLO 0.32fF
.ends

