* NGSPICE file created from largecap1.ext - technology: sky130A

X0 A B VLO sky130_fd_pr__res_xhigh_po_0p35 l=1e+08u
X1 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X2 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X3 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X4 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X5 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X6 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X7 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X8 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X9 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X10 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X11 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X12 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X13 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X14 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X15 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X16 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X17 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X18 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X19 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X20 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X21 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X22 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X23 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X24 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X25 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X26 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X27 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X28 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X29 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X30 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X31 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X32 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X33 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X34 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X35 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X36 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X37 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X38 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X39 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X40 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X41 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X42 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X43 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X44 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X45 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X46 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X47 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X48 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X49 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X50 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X51 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X52 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X53 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X54 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X55 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X56 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X57 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X58 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X59 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X60 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X61 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X62 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X63 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X64 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X65 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X66 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X67 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X68 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X69 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X70 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X71 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X72 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X73 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X74 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X75 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X76 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X77 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X78 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X79 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X80 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X81 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X82 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X83 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X84 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X85 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X86 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X87 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X88 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X89 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X90 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X91 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X92 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X93 A B sky130_fd_pr__cap_mim_m3_1 l=9.86e+07u w=4.16e+07u
X94 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X95 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
X96 B A sky130_fd_pr__cap_mim_m3_2 l=9.86e+07u w=4.16e+07u
C0 A B 30956.81fF
C1 A 0 392.52fF $ **FLOATING
C2 B 0 3661.24fF $ **FLOATING
