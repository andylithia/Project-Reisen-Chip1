magic
tech sky130A
timestamp 1671334348
<< xpolycontact >>
rect -59 -159 -24 57
rect 24 -159 59 57
<< xpolyres >>
rect -59 124 59 159
rect -59 57 -24 124
rect 24 57 59 124
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 0.5 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 8.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
