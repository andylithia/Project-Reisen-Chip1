magic
tech sky130A
magscale 1 2
timestamp 1672463705
<< error_p >>
rect 19 322 77 328
rect 19 288 31 322
rect 19 282 77 288
rect -77 -288 -19 -282
rect -77 -322 -65 -288
rect -77 -328 -19 -322
<< pwell >>
rect -263 -460 263 460
<< nmos >>
rect -63 -250 -33 250
rect 33 -250 63 250
<< ndiff >>
rect -125 238 -63 250
rect -125 -238 -113 238
rect -79 -238 -63 238
rect -125 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 125 250
rect 63 -238 79 238
rect 113 -238 125 238
rect 63 -250 125 -238
<< ndiffc >>
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
<< psubdiff >>
rect -227 390 227 424
rect -227 -390 -193 390
rect 193 -390 227 390
rect -227 -424 227 -390
<< poly >>
rect 15 322 81 338
rect 15 288 31 322
rect 65 288 81 322
rect -63 250 -33 276
rect 15 272 81 288
rect 33 250 63 272
rect -63 -272 -33 -250
rect -81 -288 -15 -272
rect 33 -276 63 -250
rect -81 -322 -65 -288
rect -31 -322 -15 -288
rect -81 -338 -15 -322
<< polycont >>
rect 31 288 65 322
rect -65 -322 -31 -288
<< locali >>
rect 15 288 31 322
rect 65 288 81 322
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
rect -81 -322 -65 -288
rect -31 -322 -15 -288
<< viali >>
rect 31 288 65 322
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect -65 -322 -31 -288
<< metal1 >>
rect 19 322 77 328
rect 19 288 31 322
rect 65 288 77 322
rect 19 282 77 288
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
rect -77 -288 -19 -282
rect -77 -322 -65 -288
rect -31 -322 -19 -288
rect -77 -328 -19 -322
<< properties >>
string FIXED_BBOX -210 -407 210 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
