magic
tech sky130A
magscale 1 2
timestamp 1671395052
<< metal1 >>
rect 380 -1000 820 22680
<< metal2 >>
rect 260 21964 440 22004
rect 400 21290 440 21964
rect 260 21250 440 21290
rect 400 20576 440 21250
rect 260 20536 440 20576
rect 400 19862 440 20536
rect 260 19822 440 19862
rect 400 19148 440 19822
rect 260 19108 440 19148
rect 400 18434 440 19108
rect 260 18394 440 18434
rect 400 17720 440 18394
rect 260 17680 440 17720
rect 400 17006 440 17680
rect 260 16966 440 17006
rect 400 16292 440 16966
rect 260 16252 440 16292
rect 400 15578 440 16252
rect 260 15538 440 15578
rect 400 14864 440 15538
rect 260 14824 440 14864
rect 400 14150 440 14824
rect 260 14110 440 14150
rect 400 13436 440 14110
rect 260 13396 440 13436
rect 400 12722 440 13396
rect 260 12682 440 12722
rect 400 12008 440 12682
rect 260 11968 440 12008
rect 400 11294 440 11968
rect 260 11254 440 11294
rect 400 10580 440 11254
rect 260 10540 440 10580
rect 400 9866 440 10540
rect 260 9826 440 9866
rect 400 9152 440 9826
rect 260 9112 440 9152
rect 400 8438 440 9112
rect 260 8398 440 8438
rect 400 7724 440 8398
rect 260 7684 440 7724
rect 400 7010 440 7684
rect 260 6970 440 7010
rect 400 6296 440 6970
rect 260 6256 440 6296
rect 400 5582 440 6256
rect 260 5542 440 5582
rect 400 4868 440 5542
rect 260 4828 440 4868
rect 400 4154 440 4828
rect 260 4114 440 4154
rect 400 3440 440 4114
rect 260 3400 440 3440
rect 400 2726 440 3400
rect 260 2686 440 2726
rect 400 2012 440 2686
rect 260 1972 440 2012
rect 400 1298 440 1972
rect 260 1258 440 1298
rect 400 584 440 1258
rect 260 544 440 584
rect 400 -130 440 544
rect 260 -170 440 -130
rect 400 -840 440 -170
rect 250 -880 440 -840
rect 400 -1060 440 -880
rect 470 21970 960 22010
rect 470 21296 510 21970
rect 470 21256 960 21296
rect 470 20582 510 21256
rect 470 20542 960 20582
rect 470 19868 510 20542
rect 470 19828 960 19868
rect 470 19154 510 19828
rect 470 19114 960 19154
rect 470 18440 510 19114
rect 470 18400 960 18440
rect 470 17726 510 18400
rect 470 17686 960 17726
rect 470 17012 510 17686
rect 470 16972 960 17012
rect 470 16298 510 16972
rect 470 16258 960 16298
rect 470 15584 510 16258
rect 470 15544 960 15584
rect 470 14870 510 15544
rect 470 14830 960 14870
rect 470 14156 510 14830
rect 470 14116 960 14156
rect 470 13442 510 14116
rect 470 13402 960 13442
rect 470 12728 510 13402
rect 470 12688 960 12728
rect 470 12014 510 12688
rect 470 11974 960 12014
rect 470 11300 510 11974
rect 470 11260 970 11300
rect 470 -1060 510 11260
rect 540 10540 950 10580
rect 540 9870 580 10540
rect 540 9830 940 9870
rect 540 9150 580 9830
rect 540 9110 950 9150
rect 540 8440 580 9110
rect 540 8400 950 8440
rect 540 7730 580 8400
rect 540 7690 970 7730
rect 540 7010 580 7690
rect 540 6970 960 7010
rect 540 6290 580 6970
rect 540 6250 950 6290
rect 540 5580 580 6250
rect 540 5540 960 5580
rect 540 -1060 580 5540
rect 610 4830 940 4870
rect 610 4150 650 4830
rect 610 4110 950 4150
rect 610 3440 650 4110
rect 610 3400 940 3440
rect 610 2730 650 3400
rect 610 2690 930 2730
rect 610 -1060 650 2690
rect 680 1970 960 2010
rect 680 1300 720 1970
rect 680 1260 950 1300
rect 680 -1060 720 1260
rect 750 540 940 580
rect 750 -1060 790 540
rect 820 -160 940 -120
rect 820 -1060 860 -160
rect 940 -1060 980 -840
<< metal3 >>
rect 460 -1080 760 23570
<< metal4 >>
rect -1200 22800 2400 23400
rect -1200 -740 -600 22800
rect 1800 -760 2400 22800
use tcap_50f  tcap_50f_0
timestamp 1671378086
transform 1 0 853 0 1 -947
box -233 -53 2220 767
use tcap_100f  tcap_100f_0
timestamp 1671378102
transform 1 0 853 0 1 -233
box -233 -53 3790 767
use tcap_200f  tcap_200f_0
timestamp 1671378131
transform 1 0 853 0 1 5479
box -269 -53 6920 767
use tcap_200f  tcap_200f_3
timestamp 1671378131
transform 1 0 853 0 1 481
box -269 -53 6920 767
use tcap_200f  tcap_200f_4
timestamp 1671378131
transform 1 0 853 0 1 1195
box -269 -53 6920 767
use tcap_200f  tcap_200f_5
timestamp 1671378131
transform 1 0 853 0 1 1909
box -269 -53 6920 767
use tcap_200f  tcap_200f_6
timestamp 1671378131
transform 1 0 853 0 1 2623
box -269 -53 6920 767
use tcap_200f  tcap_200f_7
timestamp 1671378131
transform 1 0 853 0 1 3337
box -269 -53 6920 767
use tcap_200f  tcap_200f_8
timestamp 1671378131
transform 1 0 853 0 1 4051
box -269 -53 6920 767
use tcap_200f  tcap_200f_9
timestamp 1671378131
transform 1 0 853 0 1 4765
box -269 -53 6920 767
use tcap_200f  tcap_200f_10
timestamp 1671378131
transform 1 0 853 0 1 6907
box -269 -53 6920 767
use tcap_200f  tcap_200f_11
timestamp 1671378131
transform 1 0 853 0 1 6193
box -269 -53 6920 767
use tcap_200f  tcap_200f_12
timestamp 1671378131
transform 1 0 853 0 1 8335
box -269 -53 6920 767
use tcap_200f  tcap_200f_13
timestamp 1671378131
transform 1 0 853 0 1 7621
box -269 -53 6920 767
use tcap_200f  tcap_200f_14
timestamp 1671378131
transform 1 0 853 0 1 9049
box -269 -53 6920 767
use tcap_200f  tcap_200f_15
timestamp 1671378131
transform 1 0 853 0 1 16903
box -269 -53 6920 767
use tcap_200f  tcap_200f_16
timestamp 1671378131
transform 1 0 853 0 1 9763
box -269 -53 6920 767
use tcap_200f  tcap_200f_17
timestamp 1671378131
transform 1 0 853 0 1 10477
box -269 -53 6920 767
use tcap_200f  tcap_200f_18
timestamp 1671378131
transform 1 0 853 0 1 11191
box -269 -53 6920 767
use tcap_200f  tcap_200f_19
timestamp 1671378131
transform 1 0 853 0 1 11905
box -269 -53 6920 767
use tcap_200f  tcap_200f_20
timestamp 1671378131
transform 1 0 853 0 1 12619
box -269 -53 6920 767
use tcap_200f  tcap_200f_21
timestamp 1671378131
transform 1 0 853 0 1 13333
box -269 -53 6920 767
use tcap_200f  tcap_200f_22
timestamp 1671378131
transform 1 0 853 0 1 14047
box -269 -53 6920 767
use tcap_200f  tcap_200f_23
timestamp 1671378131
transform 1 0 853 0 1 14761
box -269 -53 6920 767
use tcap_200f  tcap_200f_24
timestamp 1671378131
transform 1 0 853 0 1 15475
box -269 -53 6920 767
use tcap_200f  tcap_200f_25
timestamp 1671378131
transform 1 0 853 0 1 16189
box -269 -53 6920 767
use tcap_200f  tcap_200f_26
timestamp 1671378131
transform 1 0 853 0 1 18331
box -269 -53 6920 767
use tcap_200f  tcap_200f_27
timestamp 1671378131
transform 1 0 853 0 1 17617
box -269 -53 6920 767
use tcap_200f  tcap_200f_28
timestamp 1671378131
transform 1 0 853 0 1 19759
box -269 -53 6920 767
use tcap_200f  tcap_200f_29
timestamp 1671378131
transform 1 0 853 0 1 19045
box -269 -53 6920 767
use tcap_200f  tcap_200f_30
timestamp 1671378131
transform 1 0 853 0 1 21187
box -269 -53 6920 767
use tcap_200f  tcap_200f_31
timestamp 1671378131
transform 1 0 853 0 1 20473
box -269 -53 6920 767
use tcap_200f  tcap_200f_32
timestamp 1671378131
transform 1 0 853 0 1 21901
box -269 -53 6920 767
use tcap_200f  tcap_200f_33
timestamp 1671378131
transform -1 0 351 0 1 21901
box -269 -53 6920 767
use tcap_200f  tcap_200f_34
timestamp 1671378131
transform -1 0 351 0 1 21187
box -269 -53 6920 767
use tcap_200f  tcap_200f_35
timestamp 1671378131
transform -1 0 351 0 1 20473
box -269 -53 6920 767
use tcap_200f  tcap_200f_36
timestamp 1671378131
transform -1 0 351 0 1 19759
box -269 -53 6920 767
use tcap_200f  tcap_200f_37
timestamp 1671378131
transform -1 0 351 0 1 19045
box -269 -53 6920 767
use tcap_200f  tcap_200f_38
timestamp 1671378131
transform -1 0 351 0 1 18331
box -269 -53 6920 767
use tcap_200f  tcap_200f_39
timestamp 1671378131
transform -1 0 351 0 1 17617
box -269 -53 6920 767
use tcap_200f  tcap_200f_40
timestamp 1671378131
transform -1 0 351 0 1 16903
box -269 -53 6920 767
use tcap_200f  tcap_200f_41
timestamp 1671378131
transform -1 0 351 0 1 16189
box -269 -53 6920 767
use tcap_200f  tcap_200f_42
timestamp 1671378131
transform -1 0 351 0 1 15475
box -269 -53 6920 767
use tcap_200f  tcap_200f_43
timestamp 1671378131
transform -1 0 351 0 1 14761
box -269 -53 6920 767
use tcap_200f  tcap_200f_44
timestamp 1671378131
transform -1 0 351 0 1 14047
box -269 -53 6920 767
use tcap_200f  tcap_200f_45
timestamp 1671378131
transform -1 0 351 0 1 13333
box -269 -53 6920 767
use tcap_200f  tcap_200f_46
timestamp 1671378131
transform -1 0 351 0 1 12619
box -269 -53 6920 767
use tcap_200f  tcap_200f_47
timestamp 1671378131
transform -1 0 351 0 1 11905
box -269 -53 6920 767
use tcap_200f  tcap_200f_48
timestamp 1671378131
transform -1 0 351 0 1 11191
box -269 -53 6920 767
use tcap_200f  tcap_200f_49
timestamp 1671378131
transform -1 0 351 0 1 10477
box -269 -53 6920 767
use tcap_200f  tcap_200f_50
timestamp 1671378131
transform -1 0 351 0 1 9763
box -269 -53 6920 767
use tcap_200f  tcap_200f_51
timestamp 1671378131
transform -1 0 351 0 1 9049
box -269 -53 6920 767
use tcap_200f  tcap_200f_52
timestamp 1671378131
transform -1 0 351 0 1 8335
box -269 -53 6920 767
use tcap_200f  tcap_200f_53
timestamp 1671378131
transform -1 0 351 0 1 7621
box -269 -53 6920 767
use tcap_200f  tcap_200f_54
timestamp 1671378131
transform -1 0 351 0 1 6907
box -269 -53 6920 767
use tcap_200f  tcap_200f_55
timestamp 1671378131
transform -1 0 351 0 1 6193
box -269 -53 6920 767
use tcap_200f  tcap_200f_56
timestamp 1671378131
transform -1 0 351 0 1 5479
box -269 -53 6920 767
use tcap_200f  tcap_200f_57
timestamp 1671378131
transform -1 0 351 0 1 4765
box -269 -53 6920 767
use tcap_200f  tcap_200f_58
timestamp 1671378131
transform -1 0 351 0 1 4051
box -269 -53 6920 767
use tcap_200f  tcap_200f_59
timestamp 1671378131
transform -1 0 351 0 1 3337
box -269 -53 6920 767
use tcap_200f  tcap_200f_60
timestamp 1671378131
transform -1 0 351 0 1 2623
box -269 -53 6920 767
use tcap_200f  tcap_200f_61
timestamp 1671378131
transform -1 0 351 0 1 1909
box -269 -53 6920 767
use tcap_200f  tcap_200f_62
timestamp 1671378131
transform -1 0 351 0 1 1195
box -269 -53 6920 767
use tcap_200f  tcap_200f_63
timestamp 1671378131
transform -1 0 351 0 1 481
box -269 -53 6920 767
use tcap_200f  tcap_200f_64
timestamp 1671378131
transform -1 0 351 0 1 -233
box -269 -53 6920 767
use tcap_200f  tcap_200f_65
timestamp 1671378131
transform -1 0 351 0 1 -947
box -269 -53 6920 767
<< labels >>
rlabel metal2 400 -1060 440 -1020 1 B7
rlabel metal2 470 -1060 510 -1020 1 B6
rlabel metal2 540 -1060 580 -1020 1 B5
rlabel metal2 610 -1060 650 -1020 1 B4
rlabel metal2 680 -1060 720 -1020 1 B3
rlabel metal2 750 -1060 790 -1020 1 B2
rlabel metal2 820 -1060 860 -1020 1 B1
rlabel metal2 940 -1060 980 -1020 1 B0
rlabel metal3 460 23480 760 23570 1 VSUB
rlabel metal4 -1090 23250 -790 23340 1 C
<< end >>
