magic
tech sky130A
magscale 1 2
timestamp 1672473347
<< viali >>
rect 3249 27557 3283 27591
rect 4353 27557 4387 27591
rect 5825 27557 5859 27591
rect 7757 27557 7791 27591
rect 8493 27557 8527 27591
rect 9321 27557 9355 27591
rect 10793 27557 10827 27591
rect 11897 27557 11931 27591
rect 13369 27557 13403 27591
rect 1961 27421 1995 27455
rect 2421 27421 2455 27455
rect 3433 27421 3467 27455
rect 4537 27421 4571 27455
rect 5273 27421 5307 27455
rect 6009 27421 6043 27455
rect 6837 27421 6871 27455
rect 7573 27421 7607 27455
rect 8309 27421 8343 27455
rect 9137 27421 9171 27455
rect 9873 27421 9907 27455
rect 10609 27421 10643 27455
rect 11713 27421 11747 27455
rect 12449 27421 12483 27455
rect 13185 27421 13219 27455
rect 1777 27285 1811 27319
rect 2605 27285 2639 27319
rect 5089 27285 5123 27319
rect 7021 27285 7055 27319
rect 10057 27285 10091 27319
rect 12633 27285 12667 27319
rect 2145 27081 2179 27115
rect 3617 27081 3651 27115
rect 4353 27081 4387 27115
rect 5825 27081 5859 27115
rect 7205 27081 7239 27115
rect 7941 27081 7975 27115
rect 8677 27081 8711 27115
rect 10517 27081 10551 27115
rect 11897 27081 11931 27115
rect 14105 27081 14139 27115
rect 2329 26945 2363 26979
rect 3065 26945 3099 26979
rect 3801 26945 3835 26979
rect 4537 26945 4571 26979
rect 5273 26945 5307 26979
rect 6009 26945 6043 26979
rect 7021 26945 7055 26979
rect 7757 26945 7791 26979
rect 8493 26945 8527 26979
rect 9597 26945 9631 26979
rect 10333 26945 10367 26979
rect 11713 26945 11747 26979
rect 12449 26945 12483 26979
rect 13185 26945 13219 26979
rect 13921 26945 13955 26979
rect 2881 26809 2915 26843
rect 5089 26809 5123 26843
rect 12633 26809 12667 26843
rect 9781 26741 9815 26775
rect 13369 26741 13403 26775
rect 2513 26537 2547 26571
rect 4629 26537 4663 26571
rect 6193 26537 6227 26571
rect 7021 26537 7055 26571
rect 7757 26537 7791 26571
rect 8493 26537 8527 26571
rect 9413 26537 9447 26571
rect 10333 26537 10367 26571
rect 11069 26537 11103 26571
rect 11805 26537 11839 26571
rect 12541 26537 12575 26571
rect 1961 26469 1995 26503
rect 3157 26469 3191 26503
rect 5365 26469 5399 26503
rect 1961 26333 1995 26367
rect 2697 26333 2731 26367
rect 3249 26333 3283 26367
rect 4629 26333 4663 26367
rect 5365 26333 5399 26367
rect 6377 26333 6411 26367
rect 6837 26333 6871 26367
rect 7573 26333 7607 26367
rect 8493 26333 8527 26367
rect 9413 26333 9447 26367
rect 10241 26333 10275 26367
rect 10977 26333 11011 26367
rect 11805 26333 11839 26367
rect 12541 26333 12575 26367
rect 13093 26333 13127 26367
rect 13369 26265 13403 26299
rect 2421 25993 2455 26027
rect 6929 25993 6963 26027
rect 8493 25993 8527 26027
rect 13093 25993 13127 26027
rect 5181 25925 5215 25959
rect 1593 25857 1627 25891
rect 2605 25857 2639 25891
rect 3249 25857 3283 25891
rect 4261 25857 4295 25891
rect 5365 25857 5399 25891
rect 6837 25857 6871 25891
rect 8493 25857 8527 25891
rect 10425 25857 10459 25891
rect 10885 25857 10919 25891
rect 12173 25857 12207 25891
rect 12449 25857 12483 25891
rect 12909 25857 12943 25891
rect 13645 25857 13679 25891
rect 11069 25721 11103 25755
rect 1777 25653 1811 25687
rect 3249 25653 3283 25687
rect 4261 25653 4295 25687
rect 13645 25653 13679 25687
rect 2421 25449 2455 25483
rect 3065 25449 3099 25483
rect 4169 25449 4203 25483
rect 12817 25449 12851 25483
rect 13553 25381 13587 25415
rect 2237 25245 2271 25279
rect 3249 25245 3283 25279
rect 4353 25245 4387 25279
rect 11897 25245 11931 25279
rect 12633 25245 12667 25279
rect 13369 25245 13403 25279
rect 12081 25109 12115 25143
rect 1685 24769 1719 24803
rect 2421 24769 2455 24803
rect 12541 24769 12575 24803
rect 13093 24769 13127 24803
rect 13829 24769 13863 24803
rect 1869 24633 1903 24667
rect 2605 24633 2639 24667
rect 13277 24633 13311 24667
rect 14013 24565 14047 24599
rect 2053 24361 2087 24395
rect 13553 24361 13587 24395
rect 1869 24157 1903 24191
rect 13737 24157 13771 24191
rect 14197 23817 14231 23851
rect 14013 23681 14047 23715
rect 5365 21981 5399 22015
rect 5098 21913 5132 21947
rect 3985 21845 4019 21879
rect 5457 21641 5491 21675
rect 4077 21505 4111 21539
rect 4344 21505 4378 21539
rect 3433 21097 3467 21131
rect 4353 21097 4387 21131
rect 6745 21097 6779 21131
rect 8585 21097 8619 21131
rect 3249 20893 3283 20927
rect 4537 20893 4571 20927
rect 4721 20893 4755 20927
rect 4813 20893 4847 20927
rect 5365 20893 5399 20927
rect 7205 20893 7239 20927
rect 5632 20825 5666 20859
rect 7472 20825 7506 20859
rect 2789 20553 2823 20587
rect 6009 20553 6043 20587
rect 8769 20553 8803 20587
rect 3924 20485 3958 20519
rect 7656 20485 7690 20519
rect 4169 20417 4203 20451
rect 4629 20417 4663 20451
rect 4896 20417 4930 20451
rect 6561 20417 6595 20451
rect 6745 20417 6779 20451
rect 6929 20349 6963 20383
rect 7389 20349 7423 20383
rect 2053 20009 2087 20043
rect 4445 20009 4479 20043
rect 6745 20009 6779 20043
rect 8585 20009 8619 20043
rect 3433 19873 3467 19907
rect 4629 19805 4663 19839
rect 4905 19805 4939 19839
rect 5365 19805 5399 19839
rect 7205 19805 7239 19839
rect 3188 19737 3222 19771
rect 5632 19737 5666 19771
rect 7472 19737 7506 19771
rect 4813 19669 4847 19703
rect 4629 19465 4663 19499
rect 8769 19465 8803 19499
rect 5742 19397 5776 19431
rect 6009 19329 6043 19363
rect 7389 19329 7423 19363
rect 7656 19329 7690 19363
rect 6837 18921 6871 18955
rect 5457 18717 5491 18751
rect 5702 18649 5736 18683
rect 6653 18309 6687 18343
rect 6561 18241 6595 18275
rect 6837 18241 6871 18275
rect 7021 18037 7055 18071
rect 4353 17833 4387 17867
rect 5549 17833 5583 17867
rect 8585 17833 8619 17867
rect 5917 17697 5951 17731
rect 4537 17629 4571 17663
rect 4813 17629 4847 17663
rect 5733 17629 5767 17663
rect 5825 17629 5859 17663
rect 6009 17629 6043 17663
rect 7205 17629 7239 17663
rect 7472 17561 7506 17595
rect 4721 17493 4755 17527
rect 3709 17289 3743 17323
rect 7941 17289 7975 17323
rect 4822 17153 4856 17187
rect 5733 17153 5767 17187
rect 6561 17153 6595 17187
rect 6828 17153 6862 17187
rect 5089 17085 5123 17119
rect 5917 17085 5951 17119
rect 5549 16949 5583 16983
rect 4353 16745 4387 16779
rect 6929 16609 6963 16643
rect 7757 16609 7791 16643
rect 4169 16541 4203 16575
rect 7481 16541 7515 16575
rect 9321 16541 9355 16575
rect 5273 16473 5307 16507
rect 9137 16405 9171 16439
rect 4169 16201 4203 16235
rect 5365 16201 5399 16235
rect 8677 16201 8711 16235
rect 4353 16065 4387 16099
rect 4997 16065 5031 16099
rect 5089 16065 5123 16099
rect 7297 16065 7331 16099
rect 7564 16065 7598 16099
rect 4905 15997 4939 16031
rect 5181 15997 5215 16031
rect 6561 15657 6595 15691
rect 4721 15589 4755 15623
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 4537 15453 4571 15487
rect 4813 15453 4847 15487
rect 7665 15453 7699 15487
rect 7849 15453 7883 15487
rect 5273 15385 5307 15419
rect 4353 15317 4387 15351
rect 7481 15317 7515 15351
rect 3801 15113 3835 15147
rect 8401 15113 8435 15147
rect 9045 15113 9079 15147
rect 4914 15045 4948 15079
rect 5181 14977 5215 15011
rect 6561 14977 6595 15011
rect 6828 14977 6862 15011
rect 8585 14977 8619 15011
rect 9229 14977 9263 15011
rect 7941 14841 7975 14875
rect 6929 14569 6963 14603
rect 7389 14569 7423 14603
rect 8309 14569 8343 14603
rect 9321 14569 9355 14603
rect 4997 14433 5031 14467
rect 3985 14365 4019 14399
rect 4629 14365 4663 14399
rect 4813 14365 4847 14399
rect 5549 14365 5583 14399
rect 5816 14365 5850 14399
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 7849 14365 7883 14399
rect 8493 14365 8527 14399
rect 9137 14365 9171 14399
rect 4169 14229 4203 14263
rect 3893 14025 3927 14059
rect 5825 14025 5859 14059
rect 8401 14025 8435 14059
rect 8861 14025 8895 14059
rect 5006 13957 5040 13991
rect 5273 13889 5307 13923
rect 6009 13889 6043 13923
rect 7288 13889 7322 13923
rect 9045 13889 9079 13923
rect 7021 13821 7055 13855
rect 4813 13481 4847 13515
rect 7297 13481 7331 13515
rect 8493 13481 8527 13515
rect 9137 13481 9171 13515
rect 6193 13345 6227 13379
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 6469 13277 6503 13311
rect 6929 13277 6963 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 9321 13277 9355 13311
rect 7113 13209 7147 13243
rect 5089 12937 5123 12971
rect 6009 12937 6043 12971
rect 8493 12937 8527 12971
rect 9321 12937 9355 12971
rect 9781 12937 9815 12971
rect 4905 12801 4939 12835
rect 5549 12801 5583 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 8309 12801 8343 12835
rect 9137 12801 9171 12835
rect 9965 12801 9999 12835
rect 4721 12733 4755 12767
rect 6837 12733 6871 12767
rect 8125 12733 8159 12767
rect 8953 12733 8987 12767
rect 10149 12733 10183 12767
rect 4261 12665 4295 12699
rect 5641 12597 5675 12631
rect 4445 12393 4479 12427
rect 4629 12393 4663 12427
rect 6745 12393 6779 12427
rect 8401 12393 8435 12427
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 4261 12121 4295 12155
rect 5457 12121 5491 12155
rect 4471 12053 4505 12087
rect 4629 11849 4663 11883
rect 6745 11849 6779 11883
rect 9045 11849 9079 11883
rect 4445 11713 4479 11747
rect 5641 11713 5675 11747
rect 6561 11713 6595 11747
rect 7205 11713 7239 11747
rect 7472 11713 7506 11747
rect 9229 11713 9263 11747
rect 5917 11645 5951 11679
rect 8585 11577 8619 11611
rect 7573 11305 7607 11339
rect 6515 11237 6549 11271
rect 5549 11169 5583 11203
rect 8125 11169 8159 11203
rect 5825 11101 5859 11135
rect 6285 11101 6319 11135
rect 8033 11101 8067 11135
rect 7941 11033 7975 11067
rect 6561 10761 6595 10795
rect 8125 10761 8159 10795
rect 6929 10693 6963 10727
rect 4353 10625 4387 10659
rect 4609 10625 4643 10659
rect 7941 10625 7975 10659
rect 8769 10625 8803 10659
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 7757 10557 7791 10591
rect 8585 10489 8619 10523
rect 5733 10421 5767 10455
rect 9137 10217 9171 10251
rect 6469 10081 6503 10115
rect 6193 10013 6227 10047
rect 6929 10013 6963 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 7196 9945 7230 9979
rect 8309 9877 8343 9911
rect 7757 9673 7791 9707
rect 3985 9537 4019 9571
rect 4252 9537 4286 9571
rect 6929 9537 6963 9571
rect 7941 9537 7975 9571
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 5365 9401 5399 9435
rect 6561 9401 6595 9435
rect 4537 9129 4571 9163
rect 7297 9129 7331 9163
rect 7481 9129 7515 9163
rect 7941 9061 7975 9095
rect 6929 8993 6963 9027
rect 4721 8925 4755 8959
rect 5825 8925 5859 8959
rect 6009 8925 6043 8959
rect 8217 8925 8251 8959
rect 7941 8857 7975 8891
rect 5917 8789 5951 8823
rect 7297 8789 7331 8823
rect 8125 8789 8159 8823
rect 6009 8585 6043 8619
rect 8401 8585 8435 8619
rect 9137 8585 9171 8619
rect 7288 8517 7322 8551
rect 5733 8449 5767 8483
rect 7021 8449 7055 8483
rect 8861 8449 8895 8483
rect 6009 8381 6043 8415
rect 9137 8381 9171 8415
rect 5825 8313 5859 8347
rect 8953 8313 8987 8347
rect 4353 8041 4387 8075
rect 6745 8041 6779 8075
rect 7757 8041 7791 8075
rect 9321 8041 9355 8075
rect 9965 8041 9999 8075
rect 9137 7973 9171 8007
rect 4721 7905 4755 7939
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 5273 7837 5307 7871
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 10149 7837 10183 7871
rect 9305 7769 9339 7803
rect 9505 7769 9539 7803
rect 8125 7701 8159 7735
rect 3065 7497 3099 7531
rect 5457 7497 5491 7531
rect 8033 7497 8067 7531
rect 9321 7497 9355 7531
rect 4353 7429 4387 7463
rect 8861 7429 8895 7463
rect 5273 7361 5307 7395
rect 5549 7361 5583 7395
rect 6561 7361 6595 7395
rect 7849 7361 7883 7395
rect 8125 7361 8159 7395
rect 8953 7361 8987 7395
rect 6837 7293 6871 7327
rect 8769 7293 8803 7327
rect 7849 7225 7883 7259
rect 5089 7157 5123 7191
rect 4721 6817 4755 6851
rect 8585 6817 8619 6851
rect 9597 6817 9631 6851
rect 9689 6817 9723 6851
rect 4629 6749 4663 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 5549 6749 5583 6783
rect 8309 6749 8343 6783
rect 5816 6681 5850 6715
rect 9505 6681 9539 6715
rect 4445 6613 4479 6647
rect 4813 6613 4847 6647
rect 6929 6613 6963 6647
rect 9137 6613 9171 6647
rect 4629 6409 4663 6443
rect 5457 6409 5491 6443
rect 5733 6409 5767 6443
rect 8125 6409 8159 6443
rect 8677 6409 8711 6443
rect 3801 6341 3835 6375
rect 4261 6341 4295 6375
rect 4477 6341 4511 6375
rect 9137 6341 9171 6375
rect 3525 6273 3559 6307
rect 3617 6273 3651 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6745 6273 6779 6307
rect 7001 6273 7035 6307
rect 9045 6273 9079 6307
rect 9229 6205 9263 6239
rect 6009 6137 6043 6171
rect 3801 6069 3835 6103
rect 4445 6069 4479 6103
rect 4813 5865 4847 5899
rect 5549 5865 5583 5899
rect 6101 5865 6135 5899
rect 8585 5797 8619 5831
rect 7573 5729 7607 5763
rect 8033 5729 8067 5763
rect 4721 5661 4755 5695
rect 4997 5661 5031 5695
rect 5457 5661 5491 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 7297 5661 7331 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 4905 5593 4939 5627
rect 8309 5525 8343 5559
rect 6009 5321 6043 5355
rect 5641 5253 5675 5287
rect 5846 5253 5880 5287
rect 6929 5253 6963 5287
rect 6561 5185 6595 5219
rect 7573 5185 7607 5219
rect 7757 5185 7791 5219
rect 5825 4981 5859 5015
rect 6929 4981 6963 5015
rect 7113 4981 7147 5015
rect 7573 4981 7607 5015
rect 4813 4777 4847 4811
rect 5733 4777 5767 4811
rect 6745 4777 6779 4811
rect 9137 4777 9171 4811
rect 9689 4641 9723 4675
rect 4721 4573 4755 4607
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 6285 4573 6319 4607
rect 6561 4573 6595 4607
rect 7849 4573 7883 4607
rect 9597 4573 9631 4607
rect 8033 4505 8067 4539
rect 9505 4505 9539 4539
rect 5365 4437 5399 4471
rect 6377 4437 6411 4471
rect 5825 4233 5859 4267
rect 6561 4165 6595 4199
rect 8585 4165 8619 4199
rect 3985 4097 4019 4131
rect 4252 4097 4286 4131
rect 6009 4097 6043 4131
rect 6745 4097 6779 4131
rect 6837 4097 6871 4131
rect 7481 4097 7515 4131
rect 7757 4097 7791 4131
rect 8401 4029 8435 4063
rect 8493 4029 8527 4063
rect 6561 3961 6595 3995
rect 8953 3961 8987 3995
rect 5365 3893 5399 3927
rect 7297 3893 7331 3927
rect 7665 3893 7699 3927
rect 8493 3689 8527 3723
rect 4813 3621 4847 3655
rect 5273 3621 5307 3655
rect 4261 3553 4295 3587
rect 4353 3553 4387 3587
rect 6653 3553 6687 3587
rect 7113 3553 7147 3587
rect 7380 3485 7414 3519
rect 4445 3417 4479 3451
rect 6408 3417 6442 3451
rect 1869 3349 1903 3383
rect 13737 3349 13771 3383
rect 1777 3145 1811 3179
rect 6009 3145 6043 3179
rect 7205 3145 7239 3179
rect 7665 3145 7699 3179
rect 13461 3145 13495 3179
rect 14105 3145 14139 3179
rect 4896 3077 4930 3111
rect 1593 3009 1627 3043
rect 2237 3009 2271 3043
rect 4629 3009 4663 3043
rect 7297 3009 7331 3043
rect 13645 3009 13679 3043
rect 14289 3009 14323 3043
rect 7113 2941 7147 2975
rect 13001 2941 13035 2975
rect 3617 2873 3651 2907
rect 8125 2873 8159 2907
rect 3065 2805 3099 2839
rect 4169 2805 4203 2839
rect 8677 2805 8711 2839
rect 10701 2805 10735 2839
rect 11805 2805 11839 2839
rect 3433 2601 3467 2635
rect 6561 2601 6595 2635
rect 7481 2601 7515 2635
rect 8401 2601 8435 2635
rect 9689 2601 9723 2635
rect 10793 2601 10827 2635
rect 11897 2601 11931 2635
rect 13001 2601 13035 2635
rect 4629 2533 4663 2567
rect 6009 2533 6043 2567
rect 2237 2465 2271 2499
rect 5365 2465 5399 2499
rect 1961 2397 1995 2431
rect 3249 2397 3283 2431
rect 4445 2397 4479 2431
rect 5825 2397 5859 2431
rect 6745 2397 6779 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9873 2397 9907 2431
rect 10977 2397 11011 2431
rect 12081 2397 12115 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 5181 2329 5215 2363
rect 9229 2261 9263 2295
<< metal1 >>
rect 1104 27770 14812 27792
rect 1104 27718 2663 27770
rect 2715 27718 2727 27770
rect 2779 27718 2791 27770
rect 2843 27718 2855 27770
rect 2907 27718 2919 27770
rect 2971 27718 6090 27770
rect 6142 27718 6154 27770
rect 6206 27718 6218 27770
rect 6270 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 9517 27770
rect 9569 27718 9581 27770
rect 9633 27718 9645 27770
rect 9697 27718 9709 27770
rect 9761 27718 9773 27770
rect 9825 27718 12944 27770
rect 12996 27718 13008 27770
rect 13060 27718 13072 27770
rect 13124 27718 13136 27770
rect 13188 27718 13200 27770
rect 13252 27718 14812 27770
rect 1104 27696 14812 27718
rect 10318 27616 10324 27668
rect 10376 27656 10382 27668
rect 10376 27628 10916 27656
rect 10376 27616 10382 27628
rect 3237 27591 3295 27597
rect 3237 27557 3249 27591
rect 3283 27557 3295 27591
rect 3237 27551 3295 27557
rect 4341 27591 4399 27597
rect 4341 27557 4353 27591
rect 4387 27588 4399 27591
rect 5718 27588 5724 27600
rect 4387 27560 5724 27588
rect 4387 27557 4399 27560
rect 4341 27551 4399 27557
rect 3252 27520 3280 27551
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 5813 27591 5871 27597
rect 5813 27557 5825 27591
rect 5859 27588 5871 27591
rect 7006 27588 7012 27600
rect 5859 27560 7012 27588
rect 5859 27557 5871 27560
rect 5813 27551 5871 27557
rect 7006 27548 7012 27560
rect 7064 27548 7070 27600
rect 7745 27591 7803 27597
rect 7745 27557 7757 27591
rect 7791 27588 7803 27591
rect 8110 27588 8116 27600
rect 7791 27560 8116 27588
rect 7791 27557 7803 27560
rect 7745 27551 7803 27557
rect 8110 27548 8116 27560
rect 8168 27548 8174 27600
rect 8478 27588 8484 27600
rect 8439 27560 8484 27588
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 8938 27548 8944 27600
rect 8996 27588 9002 27600
rect 9309 27591 9367 27597
rect 9309 27588 9321 27591
rect 8996 27560 9321 27588
rect 8996 27548 9002 27560
rect 9309 27557 9321 27560
rect 9355 27557 9367 27591
rect 9309 27551 9367 27557
rect 9950 27548 9956 27600
rect 10008 27588 10014 27600
rect 10781 27591 10839 27597
rect 10781 27588 10793 27591
rect 10008 27560 10793 27588
rect 10008 27548 10014 27560
rect 10781 27557 10793 27560
rect 10827 27557 10839 27591
rect 10888 27588 10916 27628
rect 11606 27616 11612 27668
rect 11664 27656 11670 27668
rect 11664 27628 12296 27656
rect 11664 27616 11670 27628
rect 11885 27591 11943 27597
rect 11885 27588 11897 27591
rect 10888 27560 11897 27588
rect 10781 27551 10839 27557
rect 11885 27557 11897 27560
rect 11931 27557 11943 27591
rect 12268 27588 12296 27628
rect 13357 27591 13415 27597
rect 13357 27588 13369 27591
rect 12268 27560 13369 27588
rect 11885 27551 11943 27557
rect 13357 27557 13369 27560
rect 13403 27557 13415 27591
rect 13357 27551 13415 27557
rect 5350 27520 5356 27532
rect 3252 27492 5356 27520
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12032 27492 13216 27520
rect 12032 27480 12038 27492
rect 1946 27452 1952 27464
rect 1907 27424 1952 27452
rect 1946 27412 1952 27424
rect 2004 27412 2010 27464
rect 2406 27452 2412 27464
rect 2367 27424 2412 27452
rect 2406 27412 2412 27424
rect 2464 27412 2470 27464
rect 3421 27455 3479 27461
rect 3421 27421 3433 27455
rect 3467 27452 3479 27455
rect 4525 27455 4583 27461
rect 3467 27424 4476 27452
rect 3467 27421 3479 27424
rect 3421 27415 3479 27421
rect 4062 27384 4068 27396
rect 1780 27356 4068 27384
rect 1780 27325 1808 27356
rect 4062 27344 4068 27356
rect 4120 27344 4126 27396
rect 4448 27384 4476 27424
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 5166 27452 5172 27464
rect 4571 27424 5172 27452
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 5166 27412 5172 27424
rect 5224 27412 5230 27464
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27452 5319 27455
rect 5810 27452 5816 27464
rect 5307 27424 5816 27452
rect 5307 27421 5319 27424
rect 5261 27415 5319 27421
rect 5810 27412 5816 27424
rect 5868 27412 5874 27464
rect 5997 27455 6055 27461
rect 5997 27421 6009 27455
rect 6043 27421 6055 27455
rect 6822 27452 6828 27464
rect 6783 27424 6828 27452
rect 5997 27415 6055 27421
rect 5350 27384 5356 27396
rect 4448 27356 5356 27384
rect 5350 27344 5356 27356
rect 5408 27344 5414 27396
rect 6012 27384 6040 27415
rect 6822 27412 6828 27424
rect 6880 27412 6886 27464
rect 7558 27452 7564 27464
rect 7519 27424 7564 27452
rect 7558 27412 7564 27424
rect 7616 27412 7622 27464
rect 8297 27455 8355 27461
rect 8297 27421 8309 27455
rect 8343 27452 8355 27455
rect 8662 27452 8668 27464
rect 8343 27424 8668 27452
rect 8343 27421 8355 27424
rect 8297 27415 8355 27421
rect 8662 27412 8668 27424
rect 8720 27412 8726 27464
rect 9122 27452 9128 27464
rect 9083 27424 9128 27452
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 9861 27455 9919 27461
rect 9861 27421 9873 27455
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 6730 27384 6736 27396
rect 6012 27356 6736 27384
rect 6730 27344 6736 27356
rect 6788 27344 6794 27396
rect 8938 27344 8944 27396
rect 8996 27384 9002 27396
rect 9876 27384 9904 27415
rect 10502 27412 10508 27464
rect 10560 27452 10566 27464
rect 13188 27461 13216 27492
rect 10597 27455 10655 27461
rect 10597 27452 10609 27455
rect 10560 27424 10609 27452
rect 10560 27412 10566 27424
rect 10597 27421 10609 27424
rect 10643 27421 10655 27455
rect 11701 27455 11759 27461
rect 11701 27452 11713 27455
rect 10597 27415 10655 27421
rect 10704 27424 11713 27452
rect 8996 27356 9904 27384
rect 8996 27344 9002 27356
rect 10226 27344 10232 27396
rect 10284 27384 10290 27396
rect 10704 27384 10732 27424
rect 11701 27421 11713 27424
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27421 12495 27455
rect 12437 27415 12495 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 10284 27356 10732 27384
rect 10284 27344 10290 27356
rect 11606 27344 11612 27396
rect 11664 27384 11670 27396
rect 12452 27384 12480 27415
rect 11664 27356 12480 27384
rect 11664 27344 11670 27356
rect 1765 27319 1823 27325
rect 1765 27285 1777 27319
rect 1811 27285 1823 27319
rect 1765 27279 1823 27285
rect 2593 27319 2651 27325
rect 2593 27285 2605 27319
rect 2639 27316 2651 27319
rect 4614 27316 4620 27328
rect 2639 27288 4620 27316
rect 2639 27285 2651 27288
rect 2593 27279 2651 27285
rect 4614 27276 4620 27288
rect 4672 27276 4678 27328
rect 5077 27319 5135 27325
rect 5077 27285 5089 27319
rect 5123 27316 5135 27319
rect 6546 27316 6552 27328
rect 5123 27288 6552 27316
rect 5123 27285 5135 27288
rect 5077 27279 5135 27285
rect 6546 27276 6552 27288
rect 6604 27276 6610 27328
rect 7009 27319 7067 27325
rect 7009 27285 7021 27319
rect 7055 27316 7067 27319
rect 7466 27316 7472 27328
rect 7055 27288 7472 27316
rect 7055 27285 7067 27288
rect 7009 27279 7067 27285
rect 7466 27276 7472 27288
rect 7524 27276 7530 27328
rect 10045 27319 10103 27325
rect 10045 27285 10057 27319
rect 10091 27316 10103 27319
rect 10134 27316 10140 27328
rect 10091 27288 10140 27316
rect 10091 27285 10103 27288
rect 10045 27279 10103 27285
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 10594 27276 10600 27328
rect 10652 27316 10658 27328
rect 12621 27319 12679 27325
rect 12621 27316 12633 27319
rect 10652 27288 12633 27316
rect 10652 27276 10658 27288
rect 12621 27285 12633 27288
rect 12667 27285 12679 27319
rect 12621 27279 12679 27285
rect 1104 27226 14971 27248
rect 1104 27174 4376 27226
rect 4428 27174 4440 27226
rect 4492 27174 4504 27226
rect 4556 27174 4568 27226
rect 4620 27174 4632 27226
rect 4684 27174 7803 27226
rect 7855 27174 7867 27226
rect 7919 27174 7931 27226
rect 7983 27174 7995 27226
rect 8047 27174 8059 27226
rect 8111 27174 11230 27226
rect 11282 27174 11294 27226
rect 11346 27174 11358 27226
rect 11410 27174 11422 27226
rect 11474 27174 11486 27226
rect 11538 27174 14657 27226
rect 14709 27174 14721 27226
rect 14773 27174 14785 27226
rect 14837 27174 14849 27226
rect 14901 27174 14913 27226
rect 14965 27174 14971 27226
rect 1104 27152 14971 27174
rect 2133 27115 2191 27121
rect 2133 27081 2145 27115
rect 2179 27112 2191 27115
rect 3510 27112 3516 27124
rect 2179 27084 3516 27112
rect 2179 27081 2191 27084
rect 2133 27075 2191 27081
rect 3510 27072 3516 27084
rect 3568 27072 3574 27124
rect 3605 27115 3663 27121
rect 3605 27081 3617 27115
rect 3651 27081 3663 27115
rect 3605 27075 3663 27081
rect 4341 27115 4399 27121
rect 4341 27081 4353 27115
rect 4387 27112 4399 27115
rect 5626 27112 5632 27124
rect 4387 27084 5632 27112
rect 4387 27081 4399 27084
rect 4341 27075 4399 27081
rect 3620 27044 3648 27075
rect 5626 27072 5632 27084
rect 5684 27072 5690 27124
rect 5813 27115 5871 27121
rect 5813 27081 5825 27115
rect 5859 27112 5871 27115
rect 6454 27112 6460 27124
rect 5859 27084 6460 27112
rect 5859 27081 5871 27084
rect 5813 27075 5871 27081
rect 6454 27072 6460 27084
rect 6512 27072 6518 27124
rect 7190 27112 7196 27124
rect 7151 27084 7196 27112
rect 7190 27072 7196 27084
rect 7248 27072 7254 27124
rect 7650 27072 7656 27124
rect 7708 27112 7714 27124
rect 7929 27115 7987 27121
rect 7929 27112 7941 27115
rect 7708 27084 7941 27112
rect 7708 27072 7714 27084
rect 7929 27081 7941 27084
rect 7975 27081 7987 27115
rect 7929 27075 7987 27081
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 8665 27115 8723 27121
rect 8665 27112 8677 27115
rect 8444 27084 8677 27112
rect 8444 27072 8450 27084
rect 8665 27081 8677 27084
rect 8711 27081 8723 27115
rect 8665 27075 8723 27081
rect 10042 27072 10048 27124
rect 10100 27112 10106 27124
rect 10505 27115 10563 27121
rect 10505 27112 10517 27115
rect 10100 27084 10517 27112
rect 10100 27072 10106 27084
rect 10505 27081 10517 27084
rect 10551 27081 10563 27115
rect 10505 27075 10563 27081
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 11885 27115 11943 27121
rect 11885 27112 11897 27115
rect 11112 27084 11897 27112
rect 11112 27072 11118 27084
rect 11885 27081 11897 27084
rect 11931 27081 11943 27115
rect 11885 27075 11943 27081
rect 12158 27072 12164 27124
rect 12216 27112 12222 27124
rect 14093 27115 14151 27121
rect 14093 27112 14105 27115
rect 12216 27084 14105 27112
rect 12216 27072 12222 27084
rect 14093 27081 14105 27084
rect 14139 27081 14151 27115
rect 14093 27075 14151 27081
rect 5074 27044 5080 27056
rect 3620 27016 5080 27044
rect 5074 27004 5080 27016
rect 5132 27004 5138 27056
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26945 2375 26979
rect 2317 26939 2375 26945
rect 3053 26979 3111 26985
rect 3053 26945 3065 26979
rect 3099 26976 3111 26979
rect 3694 26976 3700 26988
rect 3099 26948 3700 26976
rect 3099 26945 3111 26948
rect 3053 26939 3111 26945
rect 2332 26908 2360 26939
rect 3694 26936 3700 26948
rect 3752 26936 3758 26988
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26976 3847 26979
rect 4154 26976 4160 26988
rect 3835 26948 4160 26976
rect 3835 26945 3847 26948
rect 3789 26939 3847 26945
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 4522 26976 4528 26988
rect 4483 26948 4528 26976
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 5258 26976 5264 26988
rect 5219 26948 5264 26976
rect 5258 26936 5264 26948
rect 5316 26936 5322 26988
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26976 6055 26979
rect 6914 26976 6920 26988
rect 6043 26948 6920 26976
rect 6043 26945 6055 26948
rect 5997 26939 6055 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 7006 26936 7012 26988
rect 7064 26976 7070 26988
rect 7742 26976 7748 26988
rect 7064 26948 7109 26976
rect 7703 26948 7748 26976
rect 7064 26936 7070 26948
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 8478 26976 8484 26988
rect 8439 26948 8484 26976
rect 8478 26936 8484 26948
rect 8536 26936 8542 26988
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 9585 26979 9643 26985
rect 9585 26976 9597 26979
rect 9456 26948 9597 26976
rect 9456 26936 9462 26948
rect 9585 26945 9597 26948
rect 9631 26945 9643 26979
rect 10318 26976 10324 26988
rect 10279 26948 10324 26976
rect 9585 26939 9643 26945
rect 10318 26936 10324 26948
rect 10376 26936 10382 26988
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11020 26948 11713 26976
rect 11020 26936 11026 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 11790 26936 11796 26988
rect 11848 26976 11854 26988
rect 12437 26979 12495 26985
rect 12437 26976 12449 26979
rect 11848 26948 12449 26976
rect 11848 26936 11854 26948
rect 12437 26945 12449 26948
rect 12483 26945 12495 26979
rect 12437 26939 12495 26945
rect 12526 26936 12532 26988
rect 12584 26976 12590 26988
rect 13173 26979 13231 26985
rect 13173 26976 13185 26979
rect 12584 26948 13185 26976
rect 12584 26936 12590 26948
rect 13173 26945 13185 26948
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13354 26936 13360 26988
rect 13412 26976 13418 26988
rect 13909 26979 13967 26985
rect 13909 26976 13921 26979
rect 13412 26948 13921 26976
rect 13412 26936 13418 26948
rect 13909 26945 13921 26948
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 3234 26908 3240 26920
rect 2332 26880 3240 26908
rect 3234 26868 3240 26880
rect 3292 26868 3298 26920
rect 2869 26843 2927 26849
rect 2869 26809 2881 26843
rect 2915 26840 2927 26843
rect 4246 26840 4252 26852
rect 2915 26812 4252 26840
rect 2915 26809 2927 26812
rect 2869 26803 2927 26809
rect 4246 26800 4252 26812
rect 4304 26800 4310 26852
rect 5077 26843 5135 26849
rect 5077 26809 5089 26843
rect 5123 26840 5135 26843
rect 5994 26840 6000 26852
rect 5123 26812 6000 26840
rect 5123 26809 5135 26812
rect 5077 26803 5135 26809
rect 5994 26800 6000 26812
rect 6052 26800 6058 26852
rect 11146 26800 11152 26852
rect 11204 26840 11210 26852
rect 12621 26843 12679 26849
rect 12621 26840 12633 26843
rect 11204 26812 12633 26840
rect 11204 26800 11210 26812
rect 12621 26809 12633 26812
rect 12667 26809 12679 26843
rect 12621 26803 12679 26809
rect 1946 26732 1952 26784
rect 2004 26772 2010 26784
rect 4706 26772 4712 26784
rect 2004 26744 4712 26772
rect 2004 26732 2010 26744
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 9769 26775 9827 26781
rect 9769 26741 9781 26775
rect 9815 26772 9827 26775
rect 9950 26772 9956 26784
rect 9815 26744 9956 26772
rect 9815 26741 9827 26744
rect 9769 26735 9827 26741
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 11698 26732 11704 26784
rect 11756 26772 11762 26784
rect 13357 26775 13415 26781
rect 13357 26772 13369 26775
rect 11756 26744 13369 26772
rect 11756 26732 11762 26744
rect 13357 26741 13369 26744
rect 13403 26741 13415 26775
rect 13357 26735 13415 26741
rect 1104 26682 14812 26704
rect 1104 26630 2663 26682
rect 2715 26630 2727 26682
rect 2779 26630 2791 26682
rect 2843 26630 2855 26682
rect 2907 26630 2919 26682
rect 2971 26630 6090 26682
rect 6142 26630 6154 26682
rect 6206 26630 6218 26682
rect 6270 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 9517 26682
rect 9569 26630 9581 26682
rect 9633 26630 9645 26682
rect 9697 26630 9709 26682
rect 9761 26630 9773 26682
rect 9825 26630 12944 26682
rect 12996 26630 13008 26682
rect 13060 26630 13072 26682
rect 13124 26630 13136 26682
rect 13188 26630 13200 26682
rect 13252 26630 14812 26682
rect 1104 26608 14812 26630
rect 2501 26571 2559 26577
rect 2501 26537 2513 26571
rect 2547 26568 2559 26571
rect 3418 26568 3424 26580
rect 2547 26540 3424 26568
rect 2547 26537 2559 26540
rect 2501 26531 2559 26537
rect 3418 26528 3424 26540
rect 3476 26528 3482 26580
rect 3694 26528 3700 26580
rect 3752 26568 3758 26580
rect 4617 26571 4675 26577
rect 4617 26568 4629 26571
rect 3752 26540 4629 26568
rect 3752 26528 3758 26540
rect 4617 26537 4629 26540
rect 4663 26537 4675 26571
rect 4617 26531 4675 26537
rect 5258 26528 5264 26580
rect 5316 26568 5322 26580
rect 6181 26571 6239 26577
rect 6181 26568 6193 26571
rect 5316 26540 6193 26568
rect 5316 26528 5322 26540
rect 6181 26537 6193 26540
rect 6227 26537 6239 26571
rect 7006 26568 7012 26580
rect 6967 26540 7012 26568
rect 6181 26531 6239 26537
rect 7006 26528 7012 26540
rect 7064 26528 7070 26580
rect 7742 26568 7748 26580
rect 7703 26540 7748 26568
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8481 26571 8539 26577
rect 8481 26537 8493 26571
rect 8527 26568 8539 26571
rect 9122 26568 9128 26580
rect 8527 26540 9128 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 9122 26528 9128 26540
rect 9180 26528 9186 26580
rect 9398 26568 9404 26580
rect 9359 26540 9404 26568
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 10318 26568 10324 26580
rect 10279 26540 10324 26568
rect 10318 26528 10324 26540
rect 10376 26528 10382 26580
rect 11057 26571 11115 26577
rect 11057 26537 11069 26571
rect 11103 26568 11115 26571
rect 11606 26568 11612 26580
rect 11103 26540 11612 26568
rect 11103 26537 11115 26540
rect 11057 26531 11115 26537
rect 11606 26528 11612 26540
rect 11664 26528 11670 26580
rect 11790 26568 11796 26580
rect 11751 26540 11796 26568
rect 11790 26528 11796 26540
rect 11848 26528 11854 26580
rect 12526 26568 12532 26580
rect 12487 26540 12532 26568
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 1946 26500 1952 26512
rect 1907 26472 1952 26500
rect 1946 26460 1952 26472
rect 2004 26460 2010 26512
rect 3145 26503 3203 26509
rect 3145 26469 3157 26503
rect 3191 26469 3203 26503
rect 3145 26463 3203 26469
rect 3160 26432 3188 26463
rect 4522 26460 4528 26512
rect 4580 26500 4586 26512
rect 5353 26503 5411 26509
rect 5353 26500 5365 26503
rect 4580 26472 5365 26500
rect 4580 26460 4586 26472
rect 5353 26469 5365 26472
rect 5399 26469 5411 26503
rect 5353 26463 5411 26469
rect 2700 26404 3188 26432
rect 1949 26367 2007 26373
rect 1949 26333 1961 26367
rect 1995 26364 2007 26367
rect 2222 26364 2228 26376
rect 1995 26336 2228 26364
rect 1995 26333 2007 26336
rect 1949 26327 2007 26333
rect 2222 26324 2228 26336
rect 2280 26324 2286 26376
rect 2700 26373 2728 26404
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 10502 26432 10508 26444
rect 6696 26404 10508 26432
rect 6696 26392 6702 26404
rect 2685 26367 2743 26373
rect 2685 26333 2697 26367
rect 2731 26333 2743 26367
rect 3234 26364 3240 26376
rect 3195 26336 3240 26364
rect 2685 26327 2743 26333
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 2038 26256 2044 26308
rect 2096 26296 2102 26308
rect 2406 26296 2412 26308
rect 2096 26268 2412 26296
rect 2096 26256 2102 26268
rect 2406 26256 2412 26268
rect 2464 26296 2470 26308
rect 4632 26296 4660 26327
rect 4798 26324 4804 26376
rect 4856 26364 4862 26376
rect 5166 26364 5172 26376
rect 4856 26336 5172 26364
rect 4856 26324 4862 26336
rect 5166 26324 5172 26336
rect 5224 26364 5230 26376
rect 5353 26367 5411 26373
rect 5353 26364 5365 26367
rect 5224 26336 5365 26364
rect 5224 26324 5230 26336
rect 5353 26333 5365 26336
rect 5399 26333 5411 26367
rect 5353 26327 5411 26333
rect 6365 26367 6423 26373
rect 6365 26333 6377 26367
rect 6411 26333 6423 26367
rect 6822 26364 6828 26376
rect 6783 26336 6828 26364
rect 6365 26327 6423 26333
rect 2464 26268 4660 26296
rect 6380 26296 6408 26327
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 6914 26324 6920 26376
rect 6972 26324 6978 26376
rect 7558 26364 7564 26376
rect 7519 26336 7564 26364
rect 7558 26324 7564 26336
rect 7616 26324 7622 26376
rect 8481 26367 8539 26373
rect 8481 26333 8493 26367
rect 8527 26364 8539 26367
rect 8938 26364 8944 26376
rect 8527 26336 8944 26364
rect 8527 26333 8539 26336
rect 8481 26327 8539 26333
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9416 26373 9444 26404
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 13354 26432 13360 26444
rect 12544 26404 13360 26432
rect 9401 26367 9459 26373
rect 9401 26333 9413 26367
rect 9447 26333 9459 26367
rect 10226 26364 10232 26376
rect 10187 26336 10232 26364
rect 9401 26327 9459 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 10318 26324 10324 26376
rect 10376 26364 10382 26376
rect 10962 26364 10968 26376
rect 10376 26336 10968 26364
rect 10376 26324 10382 26336
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 11606 26324 11612 26376
rect 11664 26364 11670 26376
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 11664 26336 11805 26364
rect 11664 26324 11670 26336
rect 11793 26333 11805 26336
rect 11839 26364 11851 26367
rect 11974 26364 11980 26376
rect 11839 26336 11980 26364
rect 11839 26333 11851 26336
rect 11793 26327 11851 26333
rect 11974 26324 11980 26336
rect 12032 26324 12038 26376
rect 12434 26324 12440 26376
rect 12492 26364 12498 26376
rect 12544 26373 12572 26404
rect 13354 26392 13360 26404
rect 13412 26392 13418 26444
rect 12529 26367 12587 26373
rect 12529 26364 12541 26367
rect 12492 26336 12541 26364
rect 12492 26324 12498 26336
rect 12529 26333 12541 26336
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 12618 26324 12624 26376
rect 12676 26364 12682 26376
rect 13081 26367 13139 26373
rect 13081 26364 13093 26367
rect 12676 26336 13093 26364
rect 12676 26324 12682 26336
rect 13081 26333 13093 26336
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 6932 26296 6960 26324
rect 7098 26296 7104 26308
rect 6380 26268 7104 26296
rect 2464 26256 2470 26268
rect 7098 26256 7104 26268
rect 7156 26256 7162 26308
rect 8570 26256 8576 26308
rect 8628 26296 8634 26308
rect 10244 26296 10272 26324
rect 13354 26296 13360 26308
rect 8628 26268 10272 26296
rect 13315 26268 13360 26296
rect 8628 26256 8634 26268
rect 13354 26256 13360 26268
rect 13412 26256 13418 26308
rect 6546 26188 6552 26240
rect 6604 26228 6610 26240
rect 6822 26228 6828 26240
rect 6604 26200 6828 26228
rect 6604 26188 6610 26200
rect 6822 26188 6828 26200
rect 6880 26188 6886 26240
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9950 26228 9956 26240
rect 9364 26200 9956 26228
rect 9364 26188 9370 26200
rect 9950 26188 9956 26200
rect 10008 26188 10014 26240
rect 1104 26138 14971 26160
rect 1104 26086 4376 26138
rect 4428 26086 4440 26138
rect 4492 26086 4504 26138
rect 4556 26086 4568 26138
rect 4620 26086 4632 26138
rect 4684 26086 7803 26138
rect 7855 26086 7867 26138
rect 7919 26086 7931 26138
rect 7983 26086 7995 26138
rect 8047 26086 8059 26138
rect 8111 26086 11230 26138
rect 11282 26086 11294 26138
rect 11346 26086 11358 26138
rect 11410 26086 11422 26138
rect 11474 26086 11486 26138
rect 11538 26086 14657 26138
rect 14709 26086 14721 26138
rect 14773 26086 14785 26138
rect 14837 26086 14849 26138
rect 14901 26086 14913 26138
rect 14965 26086 14971 26138
rect 1104 26064 14971 26086
rect 2409 26027 2467 26033
rect 2409 25993 2421 26027
rect 2455 26024 2467 26027
rect 3142 26024 3148 26036
rect 2455 25996 3148 26024
rect 2455 25993 2467 25996
rect 2409 25987 2467 25993
rect 3142 25984 3148 25996
rect 3200 25984 3206 26036
rect 5810 25984 5816 26036
rect 5868 26024 5874 26036
rect 6917 26027 6975 26033
rect 6917 26024 6929 26027
rect 5868 25996 6929 26024
rect 5868 25984 5874 25996
rect 6917 25993 6929 25996
rect 6963 25993 6975 26027
rect 8478 26024 8484 26036
rect 8439 25996 8484 26024
rect 6917 25987 6975 25993
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 10134 26024 10140 26036
rect 9272 25996 10140 26024
rect 9272 25984 9278 25996
rect 10134 25984 10140 25996
rect 10192 25984 10198 26036
rect 12250 25984 12256 26036
rect 12308 26024 12314 26036
rect 13081 26027 13139 26033
rect 13081 26024 13093 26027
rect 12308 25996 13093 26024
rect 12308 25984 12314 25996
rect 13081 25993 13093 25996
rect 13127 25993 13139 26027
rect 13081 25987 13139 25993
rect 4154 25916 4160 25968
rect 4212 25956 4218 25968
rect 5169 25959 5227 25965
rect 5169 25956 5181 25959
rect 4212 25928 5181 25956
rect 4212 25916 4218 25928
rect 5169 25925 5181 25928
rect 5215 25925 5227 25959
rect 5169 25919 5227 25925
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 3237 25891 3295 25897
rect 3237 25888 3249 25891
rect 2639 25860 3249 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 3237 25857 3249 25860
rect 3283 25888 3295 25891
rect 3326 25888 3332 25900
rect 3283 25860 3332 25888
rect 3283 25857 3295 25860
rect 3237 25851 3295 25857
rect 3326 25848 3332 25860
rect 3384 25848 3390 25900
rect 4246 25888 4252 25900
rect 4207 25860 4252 25888
rect 4246 25848 4252 25860
rect 4304 25888 4310 25900
rect 4706 25888 4712 25900
rect 4304 25860 4712 25888
rect 4304 25848 4310 25860
rect 4706 25848 4712 25860
rect 4764 25848 4770 25900
rect 5350 25888 5356 25900
rect 5311 25860 5356 25888
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 6822 25888 6828 25900
rect 6783 25860 6828 25888
rect 6822 25848 6828 25860
rect 6880 25848 6886 25900
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25888 8539 25891
rect 8662 25888 8668 25900
rect 8527 25860 8668 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 8662 25848 8668 25860
rect 8720 25848 8726 25900
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25888 10471 25891
rect 10870 25888 10876 25900
rect 10459 25860 10876 25888
rect 10459 25857 10471 25860
rect 10413 25851 10471 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 12158 25888 12164 25900
rect 12119 25860 12164 25888
rect 12158 25848 12164 25860
rect 12216 25848 12222 25900
rect 12437 25891 12495 25897
rect 12437 25857 12449 25891
rect 12483 25888 12495 25891
rect 12897 25891 12955 25897
rect 12897 25888 12909 25891
rect 12483 25860 12909 25888
rect 12483 25857 12495 25860
rect 12437 25851 12495 25857
rect 12897 25857 12909 25860
rect 12943 25857 12955 25891
rect 12897 25851 12955 25857
rect 13633 25891 13691 25897
rect 13633 25857 13645 25891
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 11882 25780 11888 25832
rect 11940 25820 11946 25832
rect 13648 25820 13676 25851
rect 11940 25792 13676 25820
rect 11940 25780 11946 25792
rect 11057 25755 11115 25761
rect 11057 25721 11069 25755
rect 11103 25752 11115 25755
rect 14182 25752 14188 25764
rect 11103 25724 14188 25752
rect 11103 25721 11115 25724
rect 11057 25715 11115 25721
rect 14182 25712 14188 25724
rect 14240 25712 14246 25764
rect 1762 25684 1768 25696
rect 1723 25656 1768 25684
rect 1762 25644 1768 25656
rect 1820 25644 1826 25696
rect 3234 25684 3240 25696
rect 3195 25656 3240 25684
rect 3234 25644 3240 25656
rect 3292 25644 3298 25696
rect 4249 25687 4307 25693
rect 4249 25653 4261 25687
rect 4295 25684 4307 25687
rect 4338 25684 4344 25696
rect 4295 25656 4344 25684
rect 4295 25653 4307 25656
rect 4249 25647 4307 25653
rect 4338 25644 4344 25656
rect 4396 25644 4402 25696
rect 13633 25687 13691 25693
rect 13633 25653 13645 25687
rect 13679 25684 13691 25687
rect 13722 25684 13728 25696
rect 13679 25656 13728 25684
rect 13679 25653 13691 25656
rect 13633 25647 13691 25653
rect 13722 25644 13728 25656
rect 13780 25644 13786 25696
rect 1104 25594 14812 25616
rect 1104 25542 2663 25594
rect 2715 25542 2727 25594
rect 2779 25542 2791 25594
rect 2843 25542 2855 25594
rect 2907 25542 2919 25594
rect 2971 25542 6090 25594
rect 6142 25542 6154 25594
rect 6206 25542 6218 25594
rect 6270 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 9517 25594
rect 9569 25542 9581 25594
rect 9633 25542 9645 25594
rect 9697 25542 9709 25594
rect 9761 25542 9773 25594
rect 9825 25542 12944 25594
rect 12996 25542 13008 25594
rect 13060 25542 13072 25594
rect 13124 25542 13136 25594
rect 13188 25542 13200 25594
rect 13252 25542 14812 25594
rect 1104 25520 14812 25542
rect 2409 25483 2467 25489
rect 2409 25449 2421 25483
rect 2455 25480 2467 25483
rect 2498 25480 2504 25492
rect 2455 25452 2504 25480
rect 2455 25449 2467 25452
rect 2409 25443 2467 25449
rect 2498 25440 2504 25452
rect 2556 25440 2562 25492
rect 3050 25480 3056 25492
rect 3011 25452 3056 25480
rect 3050 25440 3056 25452
rect 3108 25440 3114 25492
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 4157 25483 4215 25489
rect 4157 25480 4169 25483
rect 4028 25452 4169 25480
rect 4028 25440 4034 25452
rect 4157 25449 4169 25452
rect 4203 25449 4215 25483
rect 4157 25443 4215 25449
rect 12710 25440 12716 25492
rect 12768 25480 12774 25492
rect 12805 25483 12863 25489
rect 12805 25480 12817 25483
rect 12768 25452 12817 25480
rect 12768 25440 12774 25452
rect 12805 25449 12817 25452
rect 12851 25449 12863 25483
rect 12805 25443 12863 25449
rect 12894 25372 12900 25424
rect 12952 25412 12958 25424
rect 13541 25415 13599 25421
rect 13541 25412 13553 25415
rect 12952 25384 13553 25412
rect 12952 25372 12958 25384
rect 13541 25381 13553 25384
rect 13587 25381 13599 25415
rect 13541 25375 13599 25381
rect 2222 25276 2228 25288
rect 2135 25248 2228 25276
rect 2222 25236 2228 25248
rect 2280 25276 2286 25288
rect 3050 25276 3056 25288
rect 2280 25248 3056 25276
rect 2280 25236 2286 25248
rect 3050 25236 3056 25248
rect 3108 25236 3114 25288
rect 3234 25276 3240 25288
rect 3195 25248 3240 25276
rect 3234 25236 3240 25248
rect 3292 25236 3298 25288
rect 4338 25276 4344 25288
rect 4299 25248 4344 25276
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 11882 25276 11888 25288
rect 8812 25248 11888 25276
rect 8812 25236 8818 25248
rect 11882 25236 11888 25248
rect 11940 25236 11946 25288
rect 12158 25236 12164 25288
rect 12216 25276 12222 25288
rect 12621 25279 12679 25285
rect 12621 25276 12633 25279
rect 12216 25248 12633 25276
rect 12216 25236 12222 25248
rect 12621 25245 12633 25248
rect 12667 25245 12679 25279
rect 13354 25276 13360 25288
rect 13315 25248 13360 25276
rect 12621 25239 12679 25245
rect 13354 25236 13360 25248
rect 13412 25236 13418 25288
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 13630 25140 13636 25152
rect 12115 25112 13636 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 1104 25050 14971 25072
rect 1104 24998 4376 25050
rect 4428 24998 4440 25050
rect 4492 24998 4504 25050
rect 4556 24998 4568 25050
rect 4620 24998 4632 25050
rect 4684 24998 7803 25050
rect 7855 24998 7867 25050
rect 7919 24998 7931 25050
rect 7983 24998 7995 25050
rect 8047 24998 8059 25050
rect 8111 24998 11230 25050
rect 11282 24998 11294 25050
rect 11346 24998 11358 25050
rect 11410 24998 11422 25050
rect 11474 24998 11486 25050
rect 11538 24998 14657 25050
rect 14709 24998 14721 25050
rect 14773 24998 14785 25050
rect 14837 24998 14849 25050
rect 14901 24998 14913 25050
rect 14965 24998 14971 25050
rect 1104 24976 14971 24998
rect 1578 24760 1584 24812
rect 1636 24800 1642 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 1636 24772 1685 24800
rect 1636 24760 1642 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 1688 24732 1716 24763
rect 1946 24760 1952 24812
rect 2004 24800 2010 24812
rect 2409 24803 2467 24809
rect 2409 24800 2421 24803
rect 2004 24772 2421 24800
rect 2004 24760 2010 24772
rect 2409 24769 2421 24772
rect 2455 24769 2467 24803
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 2409 24763 2467 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 13081 24803 13139 24809
rect 13081 24800 13093 24803
rect 12860 24772 13093 24800
rect 12860 24760 12866 24772
rect 13081 24769 13093 24772
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 3878 24732 3884 24744
rect 1688 24704 3884 24732
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 12544 24732 12572 24760
rect 13832 24732 13860 24763
rect 12544 24704 13860 24732
rect 1854 24664 1860 24676
rect 1815 24636 1860 24664
rect 1854 24624 1860 24636
rect 1912 24624 1918 24676
rect 2314 24624 2320 24676
rect 2372 24664 2378 24676
rect 2593 24667 2651 24673
rect 2593 24664 2605 24667
rect 2372 24636 2605 24664
rect 2372 24624 2378 24636
rect 2593 24633 2605 24636
rect 2639 24633 2651 24667
rect 13262 24664 13268 24676
rect 13223 24636 13268 24664
rect 2593 24627 2651 24633
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 13998 24596 14004 24608
rect 13959 24568 14004 24596
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 1104 24506 14812 24528
rect 1104 24454 2663 24506
rect 2715 24454 2727 24506
rect 2779 24454 2791 24506
rect 2843 24454 2855 24506
rect 2907 24454 2919 24506
rect 2971 24454 6090 24506
rect 6142 24454 6154 24506
rect 6206 24454 6218 24506
rect 6270 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 9517 24506
rect 9569 24454 9581 24506
rect 9633 24454 9645 24506
rect 9697 24454 9709 24506
rect 9761 24454 9773 24506
rect 9825 24454 12944 24506
rect 12996 24454 13008 24506
rect 13060 24454 13072 24506
rect 13124 24454 13136 24506
rect 13188 24454 13200 24506
rect 13252 24454 14812 24506
rect 1104 24432 14812 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 2041 24395 2099 24401
rect 2041 24392 2053 24395
rect 1728 24364 2053 24392
rect 1728 24352 1734 24364
rect 2041 24361 2053 24364
rect 2087 24361 2099 24395
rect 2041 24355 2099 24361
rect 13446 24352 13452 24404
rect 13504 24392 13510 24404
rect 13541 24395 13599 24401
rect 13541 24392 13553 24395
rect 13504 24364 13553 24392
rect 13504 24352 13510 24364
rect 13541 24361 13553 24364
rect 13587 24361 13599 24395
rect 13541 24355 13599 24361
rect 1762 24148 1768 24200
rect 1820 24188 1826 24200
rect 1857 24191 1915 24197
rect 1857 24188 1869 24191
rect 1820 24160 1869 24188
rect 1820 24148 1826 24160
rect 1857 24157 1869 24160
rect 1903 24157 1915 24191
rect 13722 24188 13728 24200
rect 13683 24160 13728 24188
rect 1857 24151 1915 24157
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 1104 23962 14971 23984
rect 1104 23910 4376 23962
rect 4428 23910 4440 23962
rect 4492 23910 4504 23962
rect 4556 23910 4568 23962
rect 4620 23910 4632 23962
rect 4684 23910 7803 23962
rect 7855 23910 7867 23962
rect 7919 23910 7931 23962
rect 7983 23910 7995 23962
rect 8047 23910 8059 23962
rect 8111 23910 11230 23962
rect 11282 23910 11294 23962
rect 11346 23910 11358 23962
rect 11410 23910 11422 23962
rect 11474 23910 11486 23962
rect 11538 23910 14657 23962
rect 14709 23910 14721 23962
rect 14773 23910 14785 23962
rect 14837 23910 14849 23962
rect 14901 23910 14913 23962
rect 14965 23910 14971 23962
rect 1104 23888 14971 23910
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 14185 23851 14243 23857
rect 14185 23848 14197 23851
rect 13964 23820 14197 23848
rect 13964 23808 13970 23820
rect 14185 23817 14197 23820
rect 14231 23817 14243 23851
rect 14185 23811 14243 23817
rect 13998 23712 14004 23724
rect 13959 23684 14004 23712
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 1104 23418 14812 23440
rect 1104 23366 2663 23418
rect 2715 23366 2727 23418
rect 2779 23366 2791 23418
rect 2843 23366 2855 23418
rect 2907 23366 2919 23418
rect 2971 23366 6090 23418
rect 6142 23366 6154 23418
rect 6206 23366 6218 23418
rect 6270 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 9517 23418
rect 9569 23366 9581 23418
rect 9633 23366 9645 23418
rect 9697 23366 9709 23418
rect 9761 23366 9773 23418
rect 9825 23366 12944 23418
rect 12996 23366 13008 23418
rect 13060 23366 13072 23418
rect 13124 23366 13136 23418
rect 13188 23366 13200 23418
rect 13252 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14971 22896
rect 1104 22822 4376 22874
rect 4428 22822 4440 22874
rect 4492 22822 4504 22874
rect 4556 22822 4568 22874
rect 4620 22822 4632 22874
rect 4684 22822 7803 22874
rect 7855 22822 7867 22874
rect 7919 22822 7931 22874
rect 7983 22822 7995 22874
rect 8047 22822 8059 22874
rect 8111 22822 11230 22874
rect 11282 22822 11294 22874
rect 11346 22822 11358 22874
rect 11410 22822 11422 22874
rect 11474 22822 11486 22874
rect 11538 22822 14657 22874
rect 14709 22822 14721 22874
rect 14773 22822 14785 22874
rect 14837 22822 14849 22874
rect 14901 22822 14913 22874
rect 14965 22822 14971 22874
rect 1104 22800 14971 22822
rect 1104 22330 14812 22352
rect 1104 22278 2663 22330
rect 2715 22278 2727 22330
rect 2779 22278 2791 22330
rect 2843 22278 2855 22330
rect 2907 22278 2919 22330
rect 2971 22278 6090 22330
rect 6142 22278 6154 22330
rect 6206 22278 6218 22330
rect 6270 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 9517 22330
rect 9569 22278 9581 22330
rect 9633 22278 9645 22330
rect 9697 22278 9709 22330
rect 9761 22278 9773 22330
rect 9825 22278 12944 22330
rect 12996 22278 13008 22330
rect 13060 22278 13072 22330
rect 13124 22278 13136 22330
rect 13188 22278 13200 22330
rect 13252 22278 14812 22330
rect 1104 22256 14812 22278
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 5442 22012 5448 22024
rect 5399 21984 5448 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 3418 21904 3424 21956
rect 3476 21944 3482 21956
rect 5086 21947 5144 21953
rect 5086 21944 5098 21947
rect 3476 21916 5098 21944
rect 3476 21904 3482 21916
rect 5086 21913 5098 21916
rect 5132 21913 5144 21947
rect 5086 21907 5144 21913
rect 3326 21836 3332 21888
rect 3384 21876 3390 21888
rect 3973 21879 4031 21885
rect 3973 21876 3985 21879
rect 3384 21848 3985 21876
rect 3384 21836 3390 21848
rect 3973 21845 3985 21848
rect 4019 21845 4031 21879
rect 3973 21839 4031 21845
rect 1104 21786 14971 21808
rect 1104 21734 4376 21786
rect 4428 21734 4440 21786
rect 4492 21734 4504 21786
rect 4556 21734 4568 21786
rect 4620 21734 4632 21786
rect 4684 21734 7803 21786
rect 7855 21734 7867 21786
rect 7919 21734 7931 21786
rect 7983 21734 7995 21786
rect 8047 21734 8059 21786
rect 8111 21734 11230 21786
rect 11282 21734 11294 21786
rect 11346 21734 11358 21786
rect 11410 21734 11422 21786
rect 11474 21734 11486 21786
rect 11538 21734 14657 21786
rect 14709 21734 14721 21786
rect 14773 21734 14785 21786
rect 14837 21734 14849 21786
rect 14901 21734 14913 21786
rect 14965 21734 14971 21786
rect 1104 21712 14971 21734
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5445 21675 5503 21681
rect 5445 21672 5457 21675
rect 5408 21644 5457 21672
rect 5408 21632 5414 21644
rect 5445 21641 5457 21644
rect 5491 21641 5503 21675
rect 5445 21635 5503 21641
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21536 4123 21539
rect 4154 21536 4160 21548
rect 4111 21508 4160 21536
rect 4111 21505 4123 21508
rect 4065 21499 4123 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4338 21545 4344 21548
rect 4332 21499 4344 21545
rect 4396 21536 4402 21548
rect 4396 21508 4432 21536
rect 4338 21496 4344 21499
rect 4396 21496 4402 21508
rect 1104 21242 14812 21264
rect 1104 21190 2663 21242
rect 2715 21190 2727 21242
rect 2779 21190 2791 21242
rect 2843 21190 2855 21242
rect 2907 21190 2919 21242
rect 2971 21190 6090 21242
rect 6142 21190 6154 21242
rect 6206 21190 6218 21242
rect 6270 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 9517 21242
rect 9569 21190 9581 21242
rect 9633 21190 9645 21242
rect 9697 21190 9709 21242
rect 9761 21190 9773 21242
rect 9825 21190 12944 21242
rect 12996 21190 13008 21242
rect 13060 21190 13072 21242
rect 13124 21190 13136 21242
rect 13188 21190 13200 21242
rect 13252 21190 14812 21242
rect 1104 21168 14812 21190
rect 3418 21128 3424 21140
rect 3379 21100 3424 21128
rect 3418 21088 3424 21100
rect 3476 21088 3482 21140
rect 4338 21128 4344 21140
rect 4299 21100 4344 21128
rect 4338 21088 4344 21100
rect 4396 21088 4402 21140
rect 5718 21128 5724 21140
rect 4724 21100 5724 21128
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 4614 20924 4620 20936
rect 4571 20896 4620 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 3252 20856 3280 20887
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 4724 20933 4752 21100
rect 5718 21088 5724 21100
rect 5776 21088 5782 21140
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 6733 21131 6791 21137
rect 6733 21128 6745 21131
rect 6696 21100 6745 21128
rect 6696 21088 6702 21100
rect 6733 21097 6745 21100
rect 6779 21097 6791 21131
rect 8570 21128 8576 21140
rect 8531 21100 8576 21128
rect 6733 21091 6791 21097
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20893 4767 20927
rect 4709 20887 4767 20893
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20924 4859 20927
rect 4890 20924 4896 20936
rect 4847 20896 4896 20924
rect 4847 20893 4859 20896
rect 4801 20887 4859 20893
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 5442 20924 5448 20936
rect 5399 20896 5448 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 5442 20884 5448 20896
rect 5500 20884 5506 20936
rect 6178 20924 6184 20936
rect 5552 20896 6184 20924
rect 5552 20856 5580 20896
rect 6178 20884 6184 20896
rect 6236 20884 6242 20936
rect 7190 20924 7196 20936
rect 7151 20896 7196 20924
rect 7190 20884 7196 20896
rect 7248 20884 7254 20936
rect 3252 20828 5580 20856
rect 5620 20859 5678 20865
rect 5620 20825 5632 20859
rect 5666 20825 5678 20859
rect 5620 20819 5678 20825
rect 7460 20859 7518 20865
rect 7460 20825 7472 20859
rect 7506 20856 7518 20859
rect 9122 20856 9128 20868
rect 7506 20828 9128 20856
rect 7506 20825 7518 20828
rect 7460 20819 7518 20825
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 5644 20788 5672 20819
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 5592 20760 5672 20788
rect 5592 20748 5598 20760
rect 1104 20698 14971 20720
rect 1104 20646 4376 20698
rect 4428 20646 4440 20698
rect 4492 20646 4504 20698
rect 4556 20646 4568 20698
rect 4620 20646 4632 20698
rect 4684 20646 7803 20698
rect 7855 20646 7867 20698
rect 7919 20646 7931 20698
rect 7983 20646 7995 20698
rect 8047 20646 8059 20698
rect 8111 20646 11230 20698
rect 11282 20646 11294 20698
rect 11346 20646 11358 20698
rect 11410 20646 11422 20698
rect 11474 20646 11486 20698
rect 11538 20646 14657 20698
rect 14709 20646 14721 20698
rect 14773 20646 14785 20698
rect 14837 20646 14849 20698
rect 14901 20646 14913 20698
rect 14965 20646 14971 20698
rect 1104 20624 14971 20646
rect 2777 20587 2835 20593
rect 2777 20553 2789 20587
rect 2823 20584 2835 20587
rect 3142 20584 3148 20596
rect 2823 20556 3148 20584
rect 2823 20553 2835 20556
rect 2777 20547 2835 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 4706 20584 4712 20596
rect 4540 20556 4712 20584
rect 3912 20519 3970 20525
rect 3912 20485 3924 20519
rect 3958 20516 3970 20519
rect 4540 20516 4568 20556
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 5997 20587 6055 20593
rect 5997 20553 6009 20587
rect 6043 20584 6055 20587
rect 6546 20584 6552 20596
rect 6043 20556 6552 20584
rect 6043 20553 6055 20556
rect 5997 20547 6055 20553
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 8757 20587 8815 20593
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 12802 20584 12808 20596
rect 8803 20556 12808 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 5442 20516 5448 20528
rect 3958 20488 4568 20516
rect 4632 20488 5448 20516
rect 3958 20485 3970 20488
rect 3912 20479 3970 20485
rect 4154 20448 4160 20460
rect 4067 20420 4160 20448
rect 4154 20408 4160 20420
rect 4212 20448 4218 20460
rect 4632 20457 4660 20488
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 7644 20519 7702 20525
rect 7644 20485 7656 20519
rect 7690 20516 7702 20519
rect 8294 20516 8300 20528
rect 7690 20488 8300 20516
rect 7690 20485 7702 20488
rect 7644 20479 7702 20485
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 4212 20420 4629 20448
rect 4212 20408 4218 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 4884 20451 4942 20457
rect 4884 20417 4896 20451
rect 4930 20448 4942 20451
rect 5626 20448 5632 20460
rect 4930 20420 5632 20448
rect 4930 20417 4942 20420
rect 4884 20411 4942 20417
rect 5626 20408 5632 20420
rect 5684 20408 5690 20460
rect 6178 20408 6184 20460
rect 6236 20448 6242 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6236 20420 6561 20448
rect 6236 20408 6242 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 5810 20340 5816 20392
rect 5868 20380 5874 20392
rect 6748 20380 6776 20411
rect 5868 20352 6776 20380
rect 6917 20383 6975 20389
rect 5868 20340 5874 20352
rect 6917 20349 6929 20383
rect 6963 20349 6975 20383
rect 6917 20343 6975 20349
rect 4614 20204 4620 20256
rect 4672 20244 4678 20256
rect 6932 20244 6960 20343
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 7248 20352 7389 20380
rect 7248 20340 7254 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7377 20343 7435 20349
rect 4672 20216 6960 20244
rect 4672 20204 4678 20216
rect 1104 20154 14812 20176
rect 1104 20102 2663 20154
rect 2715 20102 2727 20154
rect 2779 20102 2791 20154
rect 2843 20102 2855 20154
rect 2907 20102 2919 20154
rect 2971 20102 6090 20154
rect 6142 20102 6154 20154
rect 6206 20102 6218 20154
rect 6270 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 9517 20154
rect 9569 20102 9581 20154
rect 9633 20102 9645 20154
rect 9697 20102 9709 20154
rect 9761 20102 9773 20154
rect 9825 20102 12944 20154
rect 12996 20102 13008 20154
rect 13060 20102 13072 20154
rect 13124 20102 13136 20154
rect 13188 20102 13200 20154
rect 13252 20102 14812 20154
rect 1104 20080 14812 20102
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20040 4491 20043
rect 5534 20040 5540 20052
rect 4479 20012 5540 20040
rect 4479 20009 4491 20012
rect 4433 20003 4491 20009
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 6733 20043 6791 20049
rect 6733 20009 6745 20043
rect 6779 20040 6791 20043
rect 7558 20040 7564 20052
rect 6779 20012 7564 20040
rect 6779 20009 6791 20012
rect 6733 20003 6791 20009
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 8573 20043 8631 20049
rect 8573 20009 8585 20043
rect 8619 20040 8631 20043
rect 12434 20040 12440 20052
rect 8619 20012 12440 20040
rect 8619 20009 8631 20012
rect 8573 20003 8631 20009
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 4154 19932 4160 19984
rect 4212 19932 4218 19984
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 4172 19904 4200 19932
rect 3467 19876 4200 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4890 19836 4896 19848
rect 4851 19808 4896 19836
rect 4617 19799 4675 19805
rect 3176 19771 3234 19777
rect 3176 19737 3188 19771
rect 3222 19768 3234 19771
rect 4632 19768 4660 19799
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19836 5411 19839
rect 5442 19836 5448 19848
rect 5399 19808 5448 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 7190 19836 7196 19848
rect 6972 19808 7196 19836
rect 6972 19796 6978 19808
rect 7190 19796 7196 19808
rect 7248 19796 7254 19848
rect 5620 19771 5678 19777
rect 5620 19768 5632 19771
rect 3222 19740 4292 19768
rect 4632 19740 5632 19768
rect 3222 19737 3234 19740
rect 3176 19731 3234 19737
rect 4264 19712 4292 19740
rect 5620 19737 5632 19740
rect 5666 19768 5678 19771
rect 6730 19768 6736 19780
rect 5666 19740 6736 19768
rect 5666 19737 5678 19740
rect 5620 19731 5678 19737
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 7460 19771 7518 19777
rect 7460 19737 7472 19771
rect 7506 19768 7518 19771
rect 8846 19768 8852 19780
rect 7506 19740 8852 19768
rect 7506 19737 7518 19740
rect 7460 19731 7518 19737
rect 8846 19728 8852 19740
rect 8904 19728 8910 19780
rect 4246 19660 4252 19712
rect 4304 19660 4310 19712
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 5902 19700 5908 19712
rect 4847 19672 5908 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 5902 19660 5908 19672
rect 5960 19660 5966 19712
rect 1104 19610 14971 19632
rect 1104 19558 4376 19610
rect 4428 19558 4440 19610
rect 4492 19558 4504 19610
rect 4556 19558 4568 19610
rect 4620 19558 4632 19610
rect 4684 19558 7803 19610
rect 7855 19558 7867 19610
rect 7919 19558 7931 19610
rect 7983 19558 7995 19610
rect 8047 19558 8059 19610
rect 8111 19558 11230 19610
rect 11282 19558 11294 19610
rect 11346 19558 11358 19610
rect 11410 19558 11422 19610
rect 11474 19558 11486 19610
rect 11538 19558 14657 19610
rect 14709 19558 14721 19610
rect 14773 19558 14785 19610
rect 14837 19558 14849 19610
rect 14901 19558 14913 19610
rect 14965 19558 14971 19610
rect 1104 19536 14971 19558
rect 4617 19499 4675 19505
rect 4617 19465 4629 19499
rect 4663 19496 4675 19499
rect 4798 19496 4804 19508
rect 4663 19468 4804 19496
rect 4663 19465 4675 19468
rect 4617 19459 4675 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 5810 19496 5816 19508
rect 4948 19468 5816 19496
rect 4948 19456 4954 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 5994 19456 6000 19508
rect 6052 19456 6058 19508
rect 8754 19496 8760 19508
rect 8715 19468 8760 19496
rect 8754 19456 8760 19468
rect 8812 19456 8818 19508
rect 5718 19388 5724 19440
rect 5776 19437 5782 19440
rect 5776 19428 5788 19437
rect 6012 19428 6040 19456
rect 5776 19400 6040 19428
rect 5776 19391 5788 19400
rect 5776 19388 5782 19391
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6914 19360 6920 19372
rect 6043 19332 6920 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6914 19320 6920 19332
rect 6972 19360 6978 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 6972 19332 7389 19360
rect 6972 19320 6978 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7644 19363 7702 19369
rect 7644 19329 7656 19363
rect 7690 19360 7702 19363
rect 9030 19360 9036 19372
rect 7690 19332 9036 19360
rect 7690 19329 7702 19332
rect 7644 19323 7702 19329
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 1104 19066 14812 19088
rect 1104 19014 2663 19066
rect 2715 19014 2727 19066
rect 2779 19014 2791 19066
rect 2843 19014 2855 19066
rect 2907 19014 2919 19066
rect 2971 19014 6090 19066
rect 6142 19014 6154 19066
rect 6206 19014 6218 19066
rect 6270 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 9517 19066
rect 9569 19014 9581 19066
rect 9633 19014 9645 19066
rect 9697 19014 9709 19066
rect 9761 19014 9773 19066
rect 9825 19014 12944 19066
rect 12996 19014 13008 19066
rect 13060 19014 13072 19066
rect 13124 19014 13136 19066
rect 13188 19014 13200 19066
rect 13252 19014 14812 19066
rect 1104 18992 14812 19014
rect 6822 18952 6828 18964
rect 6783 18924 6828 18952
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5534 18748 5540 18760
rect 5491 18720 5540 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5350 18640 5356 18692
rect 5408 18680 5414 18692
rect 5690 18683 5748 18689
rect 5690 18680 5702 18683
rect 5408 18652 5702 18680
rect 5408 18640 5414 18652
rect 5690 18649 5702 18652
rect 5736 18649 5748 18683
rect 5690 18643 5748 18649
rect 1104 18522 14971 18544
rect 1104 18470 4376 18522
rect 4428 18470 4440 18522
rect 4492 18470 4504 18522
rect 4556 18470 4568 18522
rect 4620 18470 4632 18522
rect 4684 18470 7803 18522
rect 7855 18470 7867 18522
rect 7919 18470 7931 18522
rect 7983 18470 7995 18522
rect 8047 18470 8059 18522
rect 8111 18470 11230 18522
rect 11282 18470 11294 18522
rect 11346 18470 11358 18522
rect 11410 18470 11422 18522
rect 11474 18470 11486 18522
rect 11538 18470 14657 18522
rect 14709 18470 14721 18522
rect 14773 18470 14785 18522
rect 14837 18470 14849 18522
rect 14901 18470 14913 18522
rect 14965 18470 14971 18522
rect 1104 18448 14971 18470
rect 5902 18300 5908 18352
rect 5960 18340 5966 18352
rect 6641 18343 6699 18349
rect 6641 18340 6653 18343
rect 5960 18312 6653 18340
rect 5960 18300 5966 18312
rect 6641 18309 6653 18312
rect 6687 18309 6699 18343
rect 6641 18303 6699 18309
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 5776 18244 6561 18272
rect 5776 18232 5782 18244
rect 6549 18241 6561 18244
rect 6595 18241 6607 18275
rect 6822 18272 6828 18284
rect 6783 18244 6828 18272
rect 6549 18235 6607 18241
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 7006 18068 7012 18080
rect 6967 18040 7012 18068
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 1104 17978 14812 18000
rect 1104 17926 2663 17978
rect 2715 17926 2727 17978
rect 2779 17926 2791 17978
rect 2843 17926 2855 17978
rect 2907 17926 2919 17978
rect 2971 17926 6090 17978
rect 6142 17926 6154 17978
rect 6206 17926 6218 17978
rect 6270 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 9517 17978
rect 9569 17926 9581 17978
rect 9633 17926 9645 17978
rect 9697 17926 9709 17978
rect 9761 17926 9773 17978
rect 9825 17926 12944 17978
rect 12996 17926 13008 17978
rect 13060 17926 13072 17978
rect 13124 17926 13136 17978
rect 13188 17926 13200 17978
rect 13252 17926 14812 17978
rect 1104 17904 14812 17926
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4341 17867 4399 17873
rect 4341 17864 4353 17867
rect 4304 17836 4353 17864
rect 4304 17824 4310 17836
rect 4341 17833 4353 17836
rect 4387 17833 4399 17867
rect 4341 17827 4399 17833
rect 5537 17867 5595 17873
rect 5537 17833 5549 17867
rect 5583 17864 5595 17867
rect 5626 17864 5632 17876
rect 5583 17836 5632 17864
rect 5583 17833 5595 17836
rect 5537 17827 5595 17833
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 11606 17864 11612 17876
rect 8619 17836 11612 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 5810 17796 5816 17808
rect 5723 17768 5816 17796
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4212 17632 4537 17660
rect 4212 17620 4218 17632
rect 4525 17629 4537 17632
rect 4571 17660 4583 17663
rect 4706 17660 4712 17672
rect 4571 17632 4712 17660
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 5166 17660 5172 17672
rect 4847 17632 5172 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 5166 17620 5172 17632
rect 5224 17660 5230 17672
rect 5626 17660 5632 17672
rect 5224 17632 5632 17660
rect 5224 17620 5230 17632
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5736 17669 5764 17768
rect 5810 17756 5816 17768
rect 5868 17796 5874 17808
rect 6086 17796 6092 17808
rect 5868 17768 6092 17796
rect 5868 17756 5874 17768
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 5902 17728 5908 17740
rect 5863 17700 5908 17728
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 5868 17632 5913 17660
rect 5868 17620 5874 17632
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6052 17632 6097 17660
rect 6052 17620 6058 17632
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6972 17632 7205 17660
rect 6972 17620 6978 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 4709 17527 4767 17533
rect 4709 17493 4721 17527
rect 4755 17524 4767 17527
rect 4890 17524 4896 17536
rect 4755 17496 4896 17524
rect 4755 17493 4767 17496
rect 4709 17487 4767 17493
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 6012 17524 6040 17620
rect 7460 17595 7518 17601
rect 7460 17561 7472 17595
rect 7506 17592 7518 17595
rect 9214 17592 9220 17604
rect 7506 17564 9220 17592
rect 7506 17561 7518 17564
rect 7460 17555 7518 17561
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 4948 17496 6040 17524
rect 4948 17484 4954 17496
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3108 17292 3709 17320
rect 3108 17280 3114 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 7929 17323 7987 17329
rect 7929 17289 7941 17323
rect 7975 17320 7987 17323
rect 8938 17320 8944 17332
rect 7975 17292 8944 17320
rect 7975 17289 7987 17292
rect 7929 17283 7987 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 6914 17252 6920 17264
rect 6564 17224 6920 17252
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 4810 17187 4868 17193
rect 4810 17184 4822 17187
rect 4396 17156 4822 17184
rect 4396 17144 4402 17156
rect 4810 17153 4822 17156
rect 4856 17153 4868 17187
rect 5718 17184 5724 17196
rect 5679 17156 5724 17184
rect 4810 17147 4868 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 6564 17193 6592 17224
rect 6914 17212 6920 17224
rect 6972 17212 6978 17264
rect 7006 17212 7012 17264
rect 7064 17212 7070 17264
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 5828 17156 6561 17184
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5828 17116 5856 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6816 17187 6874 17193
rect 6816 17153 6828 17187
rect 6862 17184 6874 17187
rect 7024 17184 7052 17212
rect 6862 17156 7052 17184
rect 6862 17153 6874 17156
rect 6816 17147 6874 17153
rect 5123 17088 5856 17116
rect 5905 17119 5963 17125
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 5920 17048 5948 17079
rect 5460 17020 5948 17048
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 5460 16980 5488 17020
rect 4212 16952 5488 16980
rect 5537 16983 5595 16989
rect 4212 16940 4218 16952
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 5626 16980 5632 16992
rect 5583 16952 5632 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 6086 16980 6092 16992
rect 5776 16952 6092 16980
rect 5776 16940 5782 16952
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 4338 16776 4344 16788
rect 4299 16748 4344 16776
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 6052 16680 7788 16708
rect 6052 16668 6058 16680
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 7760 16649 7788 16680
rect 7745 16643 7803 16649
rect 6972 16612 7017 16640
rect 6972 16600 6978 16612
rect 7745 16609 7757 16643
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 5644 16572 5672 16600
rect 7466 16572 7472 16584
rect 4203 16544 5672 16572
rect 7427 16544 7472 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 9306 16572 9312 16584
rect 9267 16544 9312 16572
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 5261 16507 5319 16513
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 5626 16504 5632 16516
rect 5307 16476 5632 16504
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 5626 16464 5632 16476
rect 5684 16464 5690 16516
rect 9122 16436 9128 16448
rect 9083 16408 9128 16436
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 8665 16235 8723 16241
rect 8665 16201 8677 16235
rect 8711 16232 8723 16235
rect 12158 16232 12164 16244
rect 8711 16204 12164 16232
rect 8711 16201 8723 16204
rect 8665 16195 8723 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 5902 16164 5908 16176
rect 5000 16136 5908 16164
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16096 4399 16099
rect 4706 16096 4712 16108
rect 4387 16068 4712 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 5000 16105 5028 16136
rect 5902 16124 5908 16136
rect 5960 16164 5966 16176
rect 6730 16164 6736 16176
rect 5960 16136 6736 16164
rect 5960 16124 5966 16136
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16065 5043 16099
rect 4985 16059 5043 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5810 16096 5816 16108
rect 5123 16068 5816 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6972 16068 7297 16096
rect 6972 16056 6978 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7552 16099 7610 16105
rect 7552 16065 7564 16099
rect 7598 16096 7610 16099
rect 8386 16096 8392 16108
rect 7598 16068 8392 16096
rect 7598 16065 7610 16068
rect 7552 16059 7610 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 4893 16031 4951 16037
rect 4893 15997 4905 16031
rect 4939 15997 4951 16031
rect 4893 15991 4951 15997
rect 4908 15960 4936 15991
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 5224 16000 5269 16028
rect 5224 15988 5230 16000
rect 4908 15932 5120 15960
rect 5092 15904 5120 15932
rect 5074 15852 5080 15904
rect 5132 15852 5138 15904
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 5592 15660 6561 15688
rect 5592 15648 5598 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6549 15651 6607 15657
rect 4709 15623 4767 15629
rect 4709 15589 4721 15623
rect 4755 15620 4767 15623
rect 4798 15620 4804 15632
rect 4755 15592 4804 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 4798 15580 4804 15592
rect 4856 15580 4862 15632
rect 7466 15620 7472 15632
rect 6886 15592 7472 15620
rect 4890 15552 4896 15564
rect 4540 15524 4896 15552
rect 4540 15493 4568 15524
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5074 15512 5080 15564
rect 5132 15552 5138 15564
rect 6886 15552 6914 15592
rect 7466 15580 7472 15592
rect 7524 15620 7530 15632
rect 7524 15592 7972 15620
rect 7524 15580 7530 15592
rect 7944 15561 7972 15592
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 5132 15524 6914 15552
rect 7300 15524 7757 15552
rect 5132 15512 5138 15524
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 5810 15484 5816 15496
rect 4847 15456 5816 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5810 15444 5816 15456
rect 5868 15484 5874 15496
rect 7300 15484 7328 15524
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 7650 15484 7656 15496
rect 5868 15456 7328 15484
rect 7611 15456 7656 15484
rect 5868 15444 5874 15456
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15484 7895 15487
rect 9398 15484 9404 15496
rect 7883 15456 9404 15484
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 5261 15419 5319 15425
rect 5261 15385 5273 15419
rect 5307 15416 5319 15419
rect 5626 15416 5632 15428
rect 5307 15388 5632 15416
rect 5307 15385 5319 15388
rect 5261 15379 5319 15385
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4890 15348 4896 15360
rect 4387 15320 4896 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4246 15144 4252 15156
rect 3835 15116 4252 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 8386 15144 8392 15156
rect 8347 15116 8392 15144
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 9030 15144 9036 15156
rect 8991 15116 9036 15144
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 4890 15036 4896 15088
rect 4948 15085 4954 15088
rect 4948 15076 4960 15085
rect 6914 15076 6920 15088
rect 4948 15048 4993 15076
rect 6564 15048 6920 15076
rect 4948 15039 4960 15048
rect 4948 15036 4954 15039
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 5534 15008 5540 15020
rect 5215 14980 5540 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 6564 15017 6592 15048
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6816 15011 6874 15017
rect 6816 14977 6828 15011
rect 6862 15008 6874 15011
rect 7374 15008 7380 15020
rect 6862 14980 7380 15008
rect 6862 14977 6874 14980
rect 6816 14971 6874 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 8570 15008 8576 15020
rect 8531 14980 8576 15008
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 9214 15008 9220 15020
rect 9175 14980 9220 15008
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 7929 14875 7987 14881
rect 7929 14841 7941 14875
rect 7975 14872 7987 14875
rect 8662 14872 8668 14884
rect 7975 14844 8668 14872
rect 7975 14841 7987 14844
rect 7929 14835 7987 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7098 14600 7104 14612
rect 6963 14572 7104 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7374 14600 7380 14612
rect 7335 14572 7380 14600
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 8294 14600 8300 14612
rect 8255 14572 8300 14600
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9306 14600 9312 14612
rect 9267 14572 9312 14600
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4764 14436 4997 14464
rect 4764 14424 4770 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 6788 14436 7788 14464
rect 6788 14424 6794 14436
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4019 14368 4629 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4798 14396 4804 14408
rect 4759 14368 4804 14396
rect 4617 14359 4675 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5316 14368 5549 14396
rect 5316 14356 5322 14368
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 5804 14399 5862 14405
rect 5804 14365 5816 14399
rect 5850 14396 5862 14399
rect 7466 14396 7472 14408
rect 5850 14368 7472 14396
rect 5850 14365 5862 14368
rect 5804 14359 5862 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 7760 14405 7788 14436
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 7837 14359 7895 14365
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 7576 14328 7604 14359
rect 6880 14300 7604 14328
rect 6880 14288 6886 14300
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 7650 14260 7656 14272
rect 4856 14232 7656 14260
rect 4856 14220 4862 14232
rect 7650 14220 7656 14232
rect 7708 14260 7714 14272
rect 7852 14260 7880 14359
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9398 14396 9404 14408
rect 9171 14368 9404 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 7708 14232 7880 14260
rect 7708 14220 7714 14232
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 3878 14056 3884 14068
rect 3839 14028 3884 14056
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 6822 14056 6828 14068
rect 5859 14028 6828 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14025 8447 14059
rect 8846 14056 8852 14068
rect 8807 14028 8852 14056
rect 8389 14019 8447 14025
rect 4154 13948 4160 14000
rect 4212 13988 4218 14000
rect 4994 13991 5052 13997
rect 4994 13988 5006 13991
rect 4212 13960 5006 13988
rect 4212 13948 4218 13960
rect 4994 13957 5006 13960
rect 5040 13957 5052 13991
rect 8404 13988 8432 14019
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 10318 13988 10324 14000
rect 8404 13960 10324 13988
rect 4994 13951 5052 13957
rect 10318 13948 10324 13960
rect 10376 13948 10382 14000
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 5994 13920 6000 13932
rect 5955 13892 6000 13920
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 7276 13923 7334 13929
rect 7276 13889 7288 13923
rect 7322 13920 7334 13923
rect 8754 13920 8760 13932
rect 7322 13892 8760 13920
rect 7322 13889 7334 13892
rect 7276 13883 7334 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 4798 13512 4804 13524
rect 4759 13484 4804 13512
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 5776 13484 7297 13512
rect 5776 13472 5782 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8570 13512 8576 13524
rect 8527 13484 8576 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 5166 13404 5172 13456
rect 5224 13404 5230 13456
rect 5184 13376 5212 13404
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 5000 13348 6193 13376
rect 5000 13317 5028 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13308 6515 13311
rect 6546 13308 6552 13320
rect 6503 13280 6552 13308
rect 6503 13277 6515 13280
rect 6457 13271 6515 13277
rect 5184 13240 5212 13271
rect 6546 13268 6552 13280
rect 6604 13308 6610 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6604 13280 6929 13308
rect 6604 13268 6610 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 6917 13271 6975 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 8662 13308 8668 13320
rect 8343 13280 8668 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9766 13308 9772 13320
rect 9355 13280 9772 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 6638 13240 6644 13252
rect 5184 13212 6644 13240
rect 6638 13200 6644 13212
rect 6696 13240 6702 13252
rect 7101 13243 7159 13249
rect 6696 13212 6914 13240
rect 6696 13200 6702 13212
rect 6886 13172 6914 13212
rect 7101 13209 7113 13243
rect 7147 13209 7159 13243
rect 7101 13203 7159 13209
rect 7116 13172 7144 13203
rect 6886 13144 7144 13172
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 5074 12968 5080 12980
rect 5035 12940 5080 12968
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5994 12968 6000 12980
rect 5955 12940 6000 12968
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9272 12940 9321 12968
rect 9272 12928 9278 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9766 12968 9772 12980
rect 9727 12940 9772 12968
rect 9309 12931 9367 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 4724 12872 5856 12900
rect 4724 12773 4752 12872
rect 4890 12832 4896 12844
rect 4851 12804 4896 12832
rect 4890 12792 4896 12804
rect 4948 12832 4954 12844
rect 5828 12841 5856 12872
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 4948 12804 5549 12832
rect 4948 12792 4954 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5859 12804 6561 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 8846 12832 8852 12844
rect 8343 12804 8852 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 9306 12832 9312 12844
rect 9171 12804 9312 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 4798 12764 4804 12776
rect 4755 12736 4804 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 4249 12699 4307 12705
rect 4249 12665 4261 12699
rect 4295 12696 4307 12699
rect 5442 12696 5448 12708
rect 4295 12668 5448 12696
rect 4295 12665 4307 12668
rect 4249 12659 4307 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 6840 12696 6868 12727
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7708 12736 8125 12764
rect 7708 12724 7714 12736
rect 8113 12733 8125 12736
rect 8159 12764 8171 12767
rect 8202 12764 8208 12776
rect 8159 12736 8208 12764
rect 8159 12733 8171 12736
rect 8113 12727 8171 12733
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8260 12736 8953 12764
rect 8260 12724 8266 12736
rect 8941 12733 8953 12736
rect 8987 12764 8999 12767
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 8987 12736 10149 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 9398 12696 9404 12708
rect 6840 12668 9404 12696
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 5626 12628 5632 12640
rect 5587 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 4706 12424 4712 12436
rect 4663 12396 4712 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 4448 12356 4476 12387
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 5592 12396 6745 12424
rect 5592 12384 5598 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 8389 12427 8447 12433
rect 8389 12393 8401 12427
rect 8435 12424 8447 12427
rect 9030 12424 9036 12436
rect 8435 12396 9036 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 4890 12356 4896 12368
rect 4448 12328 4896 12356
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7616 12192 8033 12220
rect 7616 12180 7622 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 8021 12183 8079 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 4246 12152 4252 12164
rect 4207 12124 4252 12152
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 5442 12152 5448 12164
rect 5403 12124 5448 12152
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 4459 12087 4517 12093
rect 4459 12053 4471 12087
rect 4505 12084 4517 12087
rect 5902 12084 5908 12096
rect 4505 12056 5908 12084
rect 4505 12053 4517 12056
rect 4459 12047 4517 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4798 11880 4804 11892
rect 4663 11852 4804 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 7558 11880 7564 11892
rect 6779 11852 7564 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8812 11852 9045 11880
rect 8812 11840 8818 11852
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 9033 11843 9091 11849
rect 4816 11812 4844 11840
rect 4816 11784 6592 11812
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4304 11716 4445 11744
rect 4304 11704 4310 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 4982 11744 4988 11756
rect 4479 11716 4988 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5626 11744 5632 11756
rect 5587 11716 5632 11744
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6564 11753 6592 11784
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6512 11716 6561 11744
rect 6512 11704 6518 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 7064 11716 7205 11744
rect 7064 11704 7070 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7460 11747 7518 11753
rect 7460 11713 7472 11747
rect 7506 11744 7518 11747
rect 8570 11744 8576 11756
rect 7506 11716 8576 11744
rect 7506 11713 7518 11716
rect 7460 11707 7518 11713
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 9214 11744 9220 11756
rect 9175 11716 9220 11744
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 5902 11676 5908 11688
rect 5863 11648 5908 11676
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 6730 11608 6736 11620
rect 5776 11580 6736 11608
rect 5776 11568 5782 11580
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 8573 11611 8631 11617
rect 8573 11577 8585 11611
rect 8619 11608 8631 11611
rect 10870 11608 10876 11620
rect 8619 11580 10876 11608
rect 8619 11577 8631 11580
rect 8573 11571 8631 11577
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 7561 11339 7619 11345
rect 7561 11336 7573 11339
rect 5960 11308 7573 11336
rect 5960 11296 5966 11308
rect 7561 11305 7573 11308
rect 7607 11305 7619 11339
rect 7561 11299 7619 11305
rect 6503 11271 6561 11277
rect 6503 11268 6515 11271
rect 5828 11240 6515 11268
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 5718 11200 5724 11212
rect 5583 11172 5724 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5828 11141 5856 11240
rect 6503 11237 6515 11240
rect 6549 11268 6561 11271
rect 6914 11268 6920 11280
rect 6549 11240 6920 11268
rect 6549 11237 6561 11240
rect 6503 11231 6561 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7248 11172 8125 11200
rect 7248 11160 7254 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6454 11132 6460 11144
rect 6319 11104 6460 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 6656 11104 8033 11132
rect 5166 11024 5172 11076
rect 5224 11064 5230 11076
rect 6656 11064 6684 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 7926 11064 7932 11076
rect 5224 11036 6684 11064
rect 7887 11036 7932 11064
rect 5224 11024 5230 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 6546 10792 6552 10804
rect 6507 10764 6552 10792
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8113 10795 8171 10801
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 9214 10792 9220 10804
rect 8159 10764 9220 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 5258 10724 5264 10736
rect 4356 10696 5264 10724
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4356 10665 4384 10696
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 7098 10724 7104 10736
rect 6963 10696 7104 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4212 10628 4353 10656
rect 4212 10616 4218 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4597 10659 4655 10665
rect 4597 10656 4609 10659
rect 4341 10619 4399 10625
rect 4448 10628 4609 10656
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4448 10588 4476 10628
rect 4597 10625 4609 10628
rect 4643 10625 4655 10659
rect 4597 10619 4655 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7616 10628 7941 10656
rect 7616 10616 7622 10628
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10656 8815 10659
rect 9122 10656 9128 10668
rect 8803 10628 9128 10656
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 4304 10560 4476 10588
rect 6472 10560 7021 10588
rect 4304 10548 4310 10560
rect 6472 10464 6500 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7009 10551 7067 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7760 10520 7788 10551
rect 8570 10520 8576 10532
rect 6972 10492 7788 10520
rect 8531 10492 8576 10520
rect 6972 10480 6978 10492
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 5721 10455 5779 10461
rect 5721 10421 5733 10455
rect 5767 10452 5779 10455
rect 6454 10452 6460 10464
rect 5767 10424 6460 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 6454 10112 6460 10124
rect 6415 10084 6460 10112
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5408 10016 6193 10044
rect 5408 10004 5414 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7006 10044 7012 10056
rect 6963 10016 7012 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 7184 9979 7242 9985
rect 7184 9945 7196 9979
rect 7230 9976 7242 9979
rect 7650 9976 7656 9988
rect 7230 9948 7656 9976
rect 7230 9945 7242 9948
rect 7184 9939 7242 9945
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 9324 9976 9352 10007
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9456 10016 9501 10044
rect 9456 10004 9462 10016
rect 13446 9976 13452 9988
rect 9324 9948 13452 9976
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8386 9908 8392 9920
rect 8343 9880 8392 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7708 9676 7757 9704
rect 7708 9664 7714 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4062 9568 4068 9580
rect 4019 9540 4068 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4240 9571 4298 9577
rect 4240 9537 4252 9571
rect 4286 9568 4298 9571
rect 4522 9568 4528 9580
rect 4286 9540 4528 9568
rect 4286 9537 4298 9540
rect 4240 9531 4298 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7190 9568 7196 9580
rect 6963 9540 7196 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7524 9540 7941 9568
rect 7524 9528 7530 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 7282 9500 7288 9512
rect 7147 9472 7288 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 5166 9392 5172 9444
rect 5224 9432 5230 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 5224 9404 5365 9432
rect 5224 9392 5230 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 6549 9435 6607 9441
rect 6549 9401 6561 9435
rect 6595 9432 6607 9435
rect 6638 9432 6644 9444
rect 6595 9404 6644 9432
rect 6595 9401 6607 9404
rect 6549 9395 6607 9401
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7024 9432 7052 9463
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 6972 9404 7052 9432
rect 6972 9392 6978 9404
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 6880 9132 7297 9160
rect 6880 9120 6886 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7285 9123 7343 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7432 9064 7941 9092
rect 7432 9052 7438 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 7929 9055 7987 9061
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 9030 9024 9036 9036
rect 6963 8996 9036 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7466 8956 7472 8968
rect 7340 8928 7472 8956
rect 7340 8916 7346 8928
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 7929 8891 7987 8897
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 9122 8888 9128 8900
rect 7975 8860 9128 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 5902 8820 5908 8832
rect 5863 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 7282 8820 7288 8832
rect 7243 8792 7288 8820
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8113 8823 8171 8829
rect 8113 8789 8125 8823
rect 8159 8820 8171 8823
rect 8754 8820 8760 8832
rect 8159 8792 8760 8820
rect 8159 8789 8171 8792
rect 8113 8783 8171 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5868 8588 6009 8616
rect 5868 8576 5874 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8585 8447 8619
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 8389 8579 8447 8585
rect 6914 8548 6920 8560
rect 5736 8520 6920 8548
rect 5736 8489 5764 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7276 8551 7334 8557
rect 7276 8517 7288 8551
rect 7322 8548 7334 8551
rect 7374 8548 7380 8560
rect 7322 8520 7380 8548
rect 7322 8517 7334 8520
rect 7276 8511 7334 8517
rect 7374 8508 7380 8520
rect 7432 8508 7438 8560
rect 8404 8548 8432 8579
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9858 8548 9864 8560
rect 8404 8520 9864 8548
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7006 8480 7012 8492
rect 6788 8452 7012 8480
rect 6788 8440 6794 8452
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7116 8452 8524 8480
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8412 6055 8415
rect 7116 8412 7144 8452
rect 6043 8384 7144 8412
rect 8496 8412 8524 8452
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8812 8452 8861 8480
rect 8812 8440 8818 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8496 8384 9137 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 9125 8381 9137 8384
rect 9171 8412 9183 8415
rect 9398 8412 9404 8424
rect 9171 8384 9404 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5776 8316 5825 8344
rect 5776 8304 5782 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7006 8344 7012 8356
rect 6880 8316 7012 8344
rect 6880 8304 6886 8316
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8938 8344 8944 8356
rect 8352 8316 8944 8344
rect 8352 8304 8358 8316
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4304 8044 4353 8072
rect 4304 8032 4310 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 6730 8072 6736 8084
rect 6691 8044 6736 8072
rect 4341 8035 4399 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7340 8044 7757 8072
rect 7340 8032 7346 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8996 8044 9321 8072
rect 8996 8032 9002 8044
rect 9309 8041 9321 8044
rect 9355 8072 9367 8075
rect 9398 8072 9404 8084
rect 9355 8044 9404 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9398 8032 9404 8044
rect 9456 8072 9462 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 9456 8044 9965 8072
rect 9456 8032 9462 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 9953 8035 10011 8041
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 9088 7976 9137 8004
rect 9088 7964 9094 7976
rect 9125 7973 9137 7976
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 5166 7936 5172 7948
rect 4755 7908 5172 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 8386 7936 8392 7948
rect 7944 7908 8392 7936
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4798 7868 4804 7880
rect 4759 7840 4804 7868
rect 4525 7831 4583 7837
rect 4540 7800 4568 7831
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5534 7868 5540 7880
rect 5307 7840 5540 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 7944 7877 7972 7908
rect 8386 7896 8392 7908
rect 8444 7936 8450 7948
rect 8444 7908 9352 7936
rect 8444 7896 8450 7908
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8294 7868 8300 7880
rect 8251 7840 8300 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 7650 7800 7656 7812
rect 4540 7772 7656 7800
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 9324 7809 9352 7908
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9916 7840 10149 7868
rect 9916 7828 9922 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 9293 7803 9352 7809
rect 9293 7769 9305 7803
rect 9339 7772 9352 7803
rect 9493 7803 9551 7809
rect 9339 7769 9351 7772
rect 9293 7763 9351 7769
rect 9493 7769 9505 7803
rect 9539 7769 9551 7803
rect 9493 7763 9551 7769
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8294 7732 8300 7744
rect 8159 7704 8300 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 9508 7732 9536 7763
rect 8628 7704 9536 7732
rect 8628 7692 8634 7704
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 4062 7528 4068 7540
rect 3099 7500 4068 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5350 7528 5356 7540
rect 4856 7500 5356 7528
rect 4856 7488 4862 7500
rect 5350 7488 5356 7500
rect 5408 7528 5414 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 5408 7500 5457 7528
rect 5408 7488 5414 7500
rect 5445 7497 5457 7500
rect 5491 7528 5503 7531
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 5491 7500 8033 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 9306 7528 9312 7540
rect 9267 7500 9312 7528
rect 8021 7491 8079 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 5626 7460 5632 7472
rect 4387 7432 5632 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 8754 7460 8760 7472
rect 8352 7432 8760 7460
rect 8352 7420 8358 7432
rect 8754 7420 8760 7432
rect 8812 7460 8818 7472
rect 8849 7463 8907 7469
rect 8849 7460 8861 7463
rect 8812 7432 8861 7460
rect 8812 7420 8818 7432
rect 8849 7429 8861 7432
rect 8895 7429 8907 7463
rect 8849 7423 8907 7429
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 5258 7392 5264 7404
rect 4672 7364 5264 7392
rect 4672 7352 4678 7364
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5592 7364 6561 7392
rect 5592 7352 5598 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 6696 7364 7849 7392
rect 6696 7352 6702 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 14090 7392 14096 7404
rect 8987 7364 14096 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5994 7324 6000 7336
rect 5224 7296 6000 7324
rect 5224 7284 5230 7296
rect 5994 7284 6000 7296
rect 6052 7324 6058 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6052 7296 6837 7324
rect 6052 7284 6058 7296
rect 6825 7293 6837 7296
rect 6871 7324 6883 7327
rect 8128 7324 8156 7355
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 6871 7296 8156 7324
rect 8757 7327 8815 7333
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7708 7228 7849 7256
rect 7708 7216 7714 7228
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 8772 7256 8800 7287
rect 9214 7256 9220 7268
rect 8772 7228 9220 7256
rect 7837 7219 7895 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 5258 6848 5264 6860
rect 4755 6820 5264 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9456 6820 9597 6848
rect 9456 6808 9462 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4632 6712 4660 6743
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4856 6752 4997 6780
rect 4856 6740 4862 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5166 6780 5172 6792
rect 5123 6752 5172 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 6730 6780 6736 6792
rect 5583 6752 6736 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 8294 6780 8300 6792
rect 8255 6752 8300 6780
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9692 6780 9720 6811
rect 9272 6752 9720 6780
rect 9272 6740 9278 6752
rect 5804 6715 5862 6721
rect 4212 6684 4568 6712
rect 4632 6684 4936 6712
rect 4212 6672 4218 6684
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4433 6647 4491 6653
rect 4433 6644 4445 6647
rect 3844 6616 4445 6644
rect 3844 6604 3850 6616
rect 4433 6613 4445 6616
rect 4479 6613 4491 6647
rect 4540 6644 4568 6684
rect 4614 6644 4620 6656
rect 4540 6616 4620 6644
rect 4433 6607 4491 6613
rect 4614 6604 4620 6616
rect 4672 6644 4678 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4672 6616 4813 6644
rect 4672 6604 4678 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4908 6644 4936 6684
rect 5804 6681 5816 6715
rect 5850 6712 5862 6715
rect 5902 6712 5908 6724
rect 5850 6684 5908 6712
rect 5850 6681 5862 6684
rect 5804 6675 5862 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 9493 6715 9551 6721
rect 9493 6681 9505 6715
rect 9539 6712 9551 6715
rect 9539 6684 12434 6712
rect 9539 6681 9551 6684
rect 9493 6675 9551 6681
rect 12406 6656 12434 6684
rect 6638 6644 6644 6656
rect 4908 6616 6644 6644
rect 4801 6607 4859 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8904 6616 9137 6644
rect 8904 6604 8910 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 12406 6616 12440 6656
rect 9125 6607 9183 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 4617 6443 4675 6449
rect 3528 6412 4384 6440
rect 3528 6313 3556 6412
rect 3786 6372 3792 6384
rect 3747 6344 3792 6372
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6341 4307 6375
rect 4356 6372 4384 6412
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4706 6440 4712 6452
rect 4663 6412 4712 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6440 5503 6443
rect 5534 6440 5540 6452
rect 5491 6412 5540 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 6914 6440 6920 6452
rect 5767 6412 6920 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8478 6440 8484 6452
rect 8159 6412 8484 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8662 6440 8668 6452
rect 8623 6412 8668 6440
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 4465 6375 4523 6381
rect 4465 6372 4477 6375
rect 4356 6344 4477 6372
rect 4249 6335 4307 6341
rect 4465 6341 4477 6344
rect 4511 6372 4523 6375
rect 4798 6372 4804 6384
rect 4511 6344 4804 6372
rect 4511 6341 4523 6344
rect 4465 6335 4523 6341
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 3620 6168 3648 6267
rect 4264 6236 4292 6335
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 8386 6332 8392 6384
rect 8444 6372 8450 6384
rect 9125 6375 9183 6381
rect 9125 6372 9137 6375
rect 8444 6344 9137 6372
rect 8444 6332 8450 6344
rect 9125 6341 9137 6344
rect 9171 6341 9183 6375
rect 9125 6335 9183 6341
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5684 6276 5729 6304
rect 5684 6264 5690 6276
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 6730 6304 6736 6316
rect 5868 6276 5913 6304
rect 6691 6276 6736 6304
rect 5868 6264 5874 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 6989 6307 7047 6313
rect 6989 6304 7001 6307
rect 6880 6276 7001 6304
rect 6880 6264 6886 6276
rect 6989 6273 7001 6276
rect 7035 6273 7047 6307
rect 6989 6267 7047 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 10962 6304 10968 6316
rect 9079 6276 10968 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 4264 6208 6776 6236
rect 5534 6168 5540 6180
rect 3620 6140 5540 6168
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 5994 6168 6000 6180
rect 5955 6140 6000 6168
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4246 6100 4252 6112
rect 3835 6072 4252 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 5074 6100 5080 6112
rect 4479 6072 5080 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 6748 6100 6776 6208
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9272 6208 9317 6236
rect 9272 6196 9278 6208
rect 7006 6100 7012 6112
rect 6748 6072 7012 6100
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 4798 5896 4804 5908
rect 4759 5868 4804 5896
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6822 5896 6828 5908
rect 6135 5868 6828 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8294 5828 8300 5840
rect 8128 5800 8300 5828
rect 5166 5760 5172 5772
rect 4724 5732 5172 5760
rect 4724 5701 4752 5732
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 5684 5732 7573 5760
rect 5684 5720 5690 5732
rect 7561 5729 7573 5732
rect 7607 5760 7619 5763
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7607 5732 8033 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4709 5655 4767 5661
rect 4816 5664 4997 5692
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4816 5624 4844 5664
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5316 5664 5457 5692
rect 5316 5652 5322 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 6273 5655 6331 5661
rect 4212 5596 4844 5624
rect 4893 5627 4951 5633
rect 4212 5584 4218 5596
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 5350 5624 5356 5636
rect 4939 5596 5356 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 6104 5556 6132 5655
rect 6288 5624 6316 5655
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 8128 5624 8156 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8570 5828 8576 5840
rect 8531 5800 8576 5828
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8294 5692 8300 5704
rect 8251 5664 8300 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9858 5692 9864 5704
rect 8435 5664 9864 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 6288 5596 8156 5624
rect 6638 5556 6644 5568
rect 5592 5528 6644 5556
rect 5592 5516 5598 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8386 5556 8392 5568
rect 8343 5528 8392 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5776 5324 6009 5352
rect 5776 5312 5782 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 5997 5315 6055 5321
rect 5626 5284 5632 5296
rect 5587 5256 5632 5284
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 5834 5287 5892 5293
rect 5834 5253 5846 5287
rect 5880 5284 5892 5287
rect 5880 5256 5948 5284
rect 5880 5253 5892 5256
rect 5834 5247 5892 5253
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 5920 5148 5948 5256
rect 6012 5216 6040 5315
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6696 5324 7696 5352
rect 6696 5312 6702 5324
rect 6914 5284 6920 5296
rect 6875 5256 6920 5284
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6012 5188 6561 5216
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7340 5188 7573 5216
rect 7340 5176 7346 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7668 5216 7696 5324
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7668 5188 7757 5216
rect 7561 5179 7619 5185
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 6822 5148 6828 5160
rect 5776 5120 6828 5148
rect 5776 5108 5782 5120
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7300 5148 7328 5176
rect 6880 5120 7328 5148
rect 6880 5108 6886 5120
rect 7006 5080 7012 5092
rect 6932 5052 7012 5080
rect 5810 5012 5816 5024
rect 5723 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 5012 5874 5024
rect 6454 5012 6460 5024
rect 5868 4984 6460 5012
rect 5868 4972 5874 4984
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 6932 5021 6960 5052
rect 7006 5040 7012 5052
rect 7064 5040 7070 5092
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 4981 6975 5015
rect 7098 5012 7104 5024
rect 7059 4984 7104 5012
rect 6917 4975 6975 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 7524 4984 7573 5012
rect 7524 4972 7530 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 5534 4808 5540 4820
rect 4847 4780 5540 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5718 4808 5724 4820
rect 5679 4780 5724 4808
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 6914 4808 6920 4820
rect 6779 4780 6920 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 8260 4780 9137 4808
rect 8260 4768 8266 4780
rect 9125 4777 9137 4780
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 5736 4672 5764 4768
rect 5736 4644 6316 4672
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4604 4770 4616
rect 4982 4604 4988 4616
rect 4764 4576 4988 4604
rect 4764 4564 4770 4576
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 6288 4613 6316 4644
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 9214 4672 9220 4684
rect 8444 4644 9220 4672
rect 8444 4632 8450 4644
rect 9214 4632 9220 4644
rect 9272 4672 9278 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9272 4644 9689 4672
rect 9272 4632 9278 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5684 4576 5825 4604
rect 5684 4564 5690 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 5828 4536 5856 4567
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6512 4576 6561 4604
rect 6512 4564 6518 4576
rect 6549 4573 6561 4576
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7432 4576 7849 4604
rect 7432 4564 7438 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 8352 4576 9597 4604
rect 8352 4564 8358 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 8021 4539 8079 4545
rect 5828 4508 6408 4536
rect 5350 4468 5356 4480
rect 5311 4440 5356 4468
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 6380 4477 6408 4508
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 8386 4536 8392 4548
rect 8067 4508 8392 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 10778 4536 10784 4548
rect 9539 4508 10784 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 6365 4471 6423 4477
rect 6365 4437 6377 4471
rect 6411 4468 6423 4471
rect 6638 4468 6644 4480
rect 6411 4440 6644 4468
rect 6411 4437 6423 4440
rect 6365 4431 6423 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 5813 4267 5871 4273
rect 5813 4233 5825 4267
rect 5859 4264 5871 4267
rect 6638 4264 6644 4276
rect 5859 4236 6644 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 6546 4196 6552 4208
rect 6507 4168 6552 4196
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 8294 4156 8300 4208
rect 8352 4156 8358 4208
rect 8573 4199 8631 4205
rect 8573 4165 8585 4199
rect 8619 4196 8631 4199
rect 9858 4196 9864 4208
rect 8619 4168 9864 4196
rect 8619 4165 8631 4168
rect 8573 4159 8631 4165
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4062 4128 4068 4140
rect 4019 4100 4068 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4246 4137 4252 4140
rect 4240 4128 4252 4137
rect 4207 4100 4252 4128
rect 4240 4091 4252 4100
rect 4246 4088 4252 4091
rect 4304 4088 4310 4140
rect 5994 4128 6000 4140
rect 5955 4100 6000 4128
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6696 4100 6745 4128
rect 6696 4088 6702 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6748 4060 6776 4091
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7466 4128 7472 4140
rect 6880 4100 6925 4128
rect 7427 4100 7472 4128
rect 6880 4088 6886 4100
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 8312 4128 8340 4156
rect 7791 4100 8340 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 8386 4060 8392 4072
rect 6748 4032 6868 4060
rect 8347 4032 8392 4060
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 6549 3995 6607 4001
rect 6549 3992 6561 3995
rect 5592 3964 6561 3992
rect 5592 3952 5598 3964
rect 6549 3961 6561 3964
rect 6595 3961 6607 3995
rect 6840 3992 6868 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 8496 3992 8524 4023
rect 6840 3964 8524 3992
rect 8941 3995 8999 4001
rect 6549 3955 6607 3961
rect 8941 3961 8953 3995
rect 8987 3992 8999 3995
rect 10042 3992 10048 4004
rect 8987 3964 10048 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5258 3924 5264 3936
rect 4396 3896 5264 3924
rect 4396 3884 4402 3896
rect 5258 3884 5264 3896
rect 5316 3924 5322 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5316 3896 5365 3924
rect 5316 3884 5322 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5353 3887 5411 3893
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 7374 3924 7380 3936
rect 7331 3896 7380 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 9030 3924 9036 3936
rect 7699 3896 9036 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 5442 3720 5448 3732
rect 3108 3692 5448 3720
rect 3108 3680 3114 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 6454 3720 6460 3732
rect 5736 3692 6460 3720
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 4890 3652 4896 3664
rect 4847 3624 4896 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5261 3655 5319 3661
rect 5261 3621 5273 3655
rect 5307 3652 5319 3655
rect 5736 3652 5764 3692
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8352 3692 8493 3720
rect 8352 3680 8358 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 5307 3624 5764 3652
rect 5307 3621 5319 3624
rect 5261 3615 5319 3621
rect 4246 3584 4252 3596
rect 4207 3556 4252 3584
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 6641 3587 6699 3593
rect 4396 3556 4441 3584
rect 4396 3544 4402 3556
rect 6641 3553 6653 3587
rect 6687 3584 6699 3587
rect 6730 3584 6736 3596
rect 6687 3556 6736 3584
rect 6687 3553 6699 3556
rect 6641 3547 6699 3553
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6788 3556 7113 3584
rect 6788 3544 6794 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7374 3525 7380 3528
rect 7368 3516 7380 3525
rect 7335 3488 7380 3516
rect 7368 3479 7380 3488
rect 7374 3476 7380 3479
rect 7432 3476 7438 3528
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4433 3451 4491 3457
rect 4433 3448 4445 3451
rect 4212 3420 4445 3448
rect 4212 3408 4218 3420
rect 4433 3417 4445 3420
rect 4479 3417 4491 3451
rect 4433 3411 4491 3417
rect 6396 3451 6454 3457
rect 6396 3417 6408 3451
rect 6442 3448 6454 3451
rect 6546 3448 6552 3460
rect 6442 3420 6552 3448
rect 6442 3417 6454 3420
rect 6396 3411 6454 3417
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 13998 3380 14004 3392
rect 13771 3352 14004 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 4246 3176 4252 3188
rect 1811 3148 4252 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5994 3176 6000 3188
rect 5955 3148 6000 3176
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 6512 3148 7205 3176
rect 6512 3136 6518 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7616 3148 7665 3176
rect 7616 3136 7622 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 7653 3139 7711 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 4884 3111 4942 3117
rect 4884 3077 4896 3111
rect 4930 3108 4942 3111
rect 5350 3108 5356 3120
rect 4930 3080 5356 3108
rect 4930 3077 4942 3080
rect 4884 3071 4942 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 750 3000 756 3052
rect 808 3040 814 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 808 3012 1593 3040
rect 808 3000 814 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1627 3012 2237 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4120 3012 4629 3040
rect 4120 3000 4126 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 8386 3040 8392 3052
rect 7331 3012 8392 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 7064 2944 7113 2972
rect 7064 2932 7070 2944
rect 7101 2941 7113 2944
rect 7147 2972 7159 2975
rect 7466 2972 7472 2984
rect 7147 2944 7472 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13648 2972 13676 3003
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14277 3043 14335 3049
rect 14277 3040 14289 3043
rect 14056 3012 14289 3040
rect 14056 3000 14062 3012
rect 14277 3009 14289 3012
rect 14323 3009 14335 3043
rect 14277 3003 14335 3009
rect 15102 2972 15108 2984
rect 13035 2944 15108 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4430 2904 4436 2916
rect 3651 2876 4436 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 7374 2864 7380 2916
rect 7432 2904 7438 2916
rect 8113 2907 8171 2913
rect 8113 2904 8125 2907
rect 7432 2876 8125 2904
rect 7432 2864 7438 2876
rect 8113 2873 8125 2876
rect 8159 2873 8171 2907
rect 8113 2867 8171 2873
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3234 2836 3240 2848
rect 3099 2808 3240 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 5810 2836 5816 2848
rect 4203 2808 5816 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8536 2808 8677 2836
rect 8536 2796 8542 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 10686 2836 10692 2848
rect 10647 2808 10692 2836
rect 8665 2799 8723 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11790 2836 11796 2848
rect 11751 2808 11796 2836
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 4154 2632 4160 2644
rect 3467 2604 4160 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 6546 2632 6552 2644
rect 6507 2604 6552 2632
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7248 2604 7481 2632
rect 7248 2592 7254 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 7469 2595 7527 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9677 2635 9735 2641
rect 9677 2601 9689 2635
rect 9723 2632 9735 2635
rect 9858 2632 9864 2644
rect 9723 2604 9864 2632
rect 9723 2601 9735 2604
rect 9677 2595 9735 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11020 2604 11897 2632
rect 11020 2592 11026 2604
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12492 2604 13001 2632
rect 12492 2592 12498 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 12989 2595 13047 2601
rect 4614 2564 4620 2576
rect 4575 2536 4620 2564
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 7282 2564 7288 2576
rect 6043 2536 7288 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 7282 2524 7288 2536
rect 7340 2524 7346 2576
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 4706 2496 4712 2508
rect 2271 2468 4712 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 7006 2496 7012 2508
rect 5399 2468 7012 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1912 2400 1961 2428
rect 1912 2388 1918 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 3234 2428 3240 2440
rect 3147 2400 3240 2428
rect 1949 2391 2007 2397
rect 3234 2388 3240 2400
rect 3292 2428 3298 2440
rect 4062 2428 4068 2440
rect 3292 2400 4068 2428
rect 3292 2388 3298 2400
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4430 2428 4436 2440
rect 4343 2400 4436 2428
rect 4430 2388 4436 2400
rect 4488 2428 4494 2440
rect 5074 2428 5080 2440
rect 4488 2400 5080 2428
rect 4488 2388 4494 2400
rect 5074 2388 5080 2400
rect 5132 2388 5138 2440
rect 5810 2428 5816 2440
rect 5723 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2428 5874 2440
rect 6270 2428 6276 2440
rect 5868 2400 6276 2428
rect 5868 2388 5874 2400
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7098 2428 7104 2440
rect 6779 2400 7104 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7432 2400 7665 2428
rect 7432 2388 7438 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8536 2400 8585 2428
rect 8536 2388 8542 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 8573 2391 8631 2397
rect 9600 2400 9873 2428
rect 4246 2320 4252 2372
rect 4304 2360 4310 2372
rect 5169 2363 5227 2369
rect 5169 2360 5181 2363
rect 4304 2332 5181 2360
rect 4304 2320 4310 2332
rect 5169 2329 5181 2332
rect 5215 2329 5227 2363
rect 5169 2323 5227 2329
rect 9600 2304 9628 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10744 2400 10977 2428
rect 10744 2388 10750 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11848 2400 12081 2428
rect 11848 2388 11854 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12952 2400 13185 2428
rect 12952 2388 12958 2400
rect 13173 2397 13185 2400
rect 13219 2428 13231 2431
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13219 2400 13645 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2292 9275 2295
rect 9582 2292 9588 2304
rect 9263 2264 9588 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
<< via1 >>
rect 2663 27718 2715 27770
rect 2727 27718 2779 27770
rect 2791 27718 2843 27770
rect 2855 27718 2907 27770
rect 2919 27718 2971 27770
rect 6090 27718 6142 27770
rect 6154 27718 6206 27770
rect 6218 27718 6270 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 9517 27718 9569 27770
rect 9581 27718 9633 27770
rect 9645 27718 9697 27770
rect 9709 27718 9761 27770
rect 9773 27718 9825 27770
rect 12944 27718 12996 27770
rect 13008 27718 13060 27770
rect 13072 27718 13124 27770
rect 13136 27718 13188 27770
rect 13200 27718 13252 27770
rect 10324 27616 10376 27668
rect 5724 27548 5776 27600
rect 7012 27548 7064 27600
rect 8116 27548 8168 27600
rect 8484 27591 8536 27600
rect 8484 27557 8493 27591
rect 8493 27557 8527 27591
rect 8527 27557 8536 27591
rect 8484 27548 8536 27557
rect 8944 27548 8996 27600
rect 9956 27548 10008 27600
rect 11612 27616 11664 27668
rect 5356 27480 5408 27532
rect 11980 27480 12032 27532
rect 1952 27455 2004 27464
rect 1952 27421 1961 27455
rect 1961 27421 1995 27455
rect 1995 27421 2004 27455
rect 1952 27412 2004 27421
rect 2412 27455 2464 27464
rect 2412 27421 2421 27455
rect 2421 27421 2455 27455
rect 2455 27421 2464 27455
rect 2412 27412 2464 27421
rect 4068 27344 4120 27396
rect 5172 27412 5224 27464
rect 5816 27412 5868 27464
rect 6828 27455 6880 27464
rect 5356 27344 5408 27396
rect 6828 27421 6837 27455
rect 6837 27421 6871 27455
rect 6871 27421 6880 27455
rect 6828 27412 6880 27421
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 7564 27412 7616 27421
rect 8668 27412 8720 27464
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 6736 27344 6788 27396
rect 8944 27344 8996 27396
rect 10508 27412 10560 27464
rect 10232 27344 10284 27396
rect 11612 27344 11664 27396
rect 4620 27276 4672 27328
rect 6552 27276 6604 27328
rect 7472 27276 7524 27328
rect 10140 27276 10192 27328
rect 10600 27276 10652 27328
rect 4376 27174 4428 27226
rect 4440 27174 4492 27226
rect 4504 27174 4556 27226
rect 4568 27174 4620 27226
rect 4632 27174 4684 27226
rect 7803 27174 7855 27226
rect 7867 27174 7919 27226
rect 7931 27174 7983 27226
rect 7995 27174 8047 27226
rect 8059 27174 8111 27226
rect 11230 27174 11282 27226
rect 11294 27174 11346 27226
rect 11358 27174 11410 27226
rect 11422 27174 11474 27226
rect 11486 27174 11538 27226
rect 14657 27174 14709 27226
rect 14721 27174 14773 27226
rect 14785 27174 14837 27226
rect 14849 27174 14901 27226
rect 14913 27174 14965 27226
rect 3516 27072 3568 27124
rect 5632 27072 5684 27124
rect 6460 27072 6512 27124
rect 7196 27115 7248 27124
rect 7196 27081 7205 27115
rect 7205 27081 7239 27115
rect 7239 27081 7248 27115
rect 7196 27072 7248 27081
rect 7656 27072 7708 27124
rect 8392 27072 8444 27124
rect 10048 27072 10100 27124
rect 11060 27072 11112 27124
rect 12164 27072 12216 27124
rect 5080 27004 5132 27056
rect 3700 26936 3752 26988
rect 4160 26936 4212 26988
rect 4528 26979 4580 26988
rect 4528 26945 4537 26979
rect 4537 26945 4571 26979
rect 4571 26945 4580 26979
rect 4528 26936 4580 26945
rect 5264 26979 5316 26988
rect 5264 26945 5273 26979
rect 5273 26945 5307 26979
rect 5307 26945 5316 26979
rect 5264 26936 5316 26945
rect 6920 26936 6972 26988
rect 7012 26979 7064 26988
rect 7012 26945 7021 26979
rect 7021 26945 7055 26979
rect 7055 26945 7064 26979
rect 7748 26979 7800 26988
rect 7012 26936 7064 26945
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 8484 26979 8536 26988
rect 8484 26945 8493 26979
rect 8493 26945 8527 26979
rect 8527 26945 8536 26979
rect 8484 26936 8536 26945
rect 9404 26936 9456 26988
rect 10324 26979 10376 26988
rect 10324 26945 10333 26979
rect 10333 26945 10367 26979
rect 10367 26945 10376 26979
rect 10324 26936 10376 26945
rect 10968 26936 11020 26988
rect 11796 26936 11848 26988
rect 12532 26936 12584 26988
rect 13360 26936 13412 26988
rect 3240 26868 3292 26920
rect 4252 26800 4304 26852
rect 6000 26800 6052 26852
rect 11152 26800 11204 26852
rect 1952 26732 2004 26784
rect 4712 26732 4764 26784
rect 9956 26732 10008 26784
rect 11704 26732 11756 26784
rect 2663 26630 2715 26682
rect 2727 26630 2779 26682
rect 2791 26630 2843 26682
rect 2855 26630 2907 26682
rect 2919 26630 2971 26682
rect 6090 26630 6142 26682
rect 6154 26630 6206 26682
rect 6218 26630 6270 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 9517 26630 9569 26682
rect 9581 26630 9633 26682
rect 9645 26630 9697 26682
rect 9709 26630 9761 26682
rect 9773 26630 9825 26682
rect 12944 26630 12996 26682
rect 13008 26630 13060 26682
rect 13072 26630 13124 26682
rect 13136 26630 13188 26682
rect 13200 26630 13252 26682
rect 3424 26528 3476 26580
rect 3700 26528 3752 26580
rect 5264 26528 5316 26580
rect 7012 26571 7064 26580
rect 7012 26537 7021 26571
rect 7021 26537 7055 26571
rect 7055 26537 7064 26571
rect 7012 26528 7064 26537
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 9128 26528 9180 26580
rect 9404 26571 9456 26580
rect 9404 26537 9413 26571
rect 9413 26537 9447 26571
rect 9447 26537 9456 26571
rect 9404 26528 9456 26537
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 11612 26528 11664 26580
rect 11796 26571 11848 26580
rect 11796 26537 11805 26571
rect 11805 26537 11839 26571
rect 11839 26537 11848 26571
rect 11796 26528 11848 26537
rect 12532 26571 12584 26580
rect 12532 26537 12541 26571
rect 12541 26537 12575 26571
rect 12575 26537 12584 26571
rect 12532 26528 12584 26537
rect 1952 26503 2004 26512
rect 1952 26469 1961 26503
rect 1961 26469 1995 26503
rect 1995 26469 2004 26503
rect 1952 26460 2004 26469
rect 4528 26460 4580 26512
rect 2228 26324 2280 26376
rect 6644 26392 6696 26444
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 2044 26256 2096 26308
rect 2412 26256 2464 26308
rect 4804 26324 4856 26376
rect 5172 26324 5224 26376
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 6920 26324 6972 26376
rect 7564 26367 7616 26376
rect 7564 26333 7573 26367
rect 7573 26333 7607 26367
rect 7607 26333 7616 26367
rect 7564 26324 7616 26333
rect 8944 26324 8996 26376
rect 10508 26392 10560 26444
rect 10232 26367 10284 26376
rect 10232 26333 10241 26367
rect 10241 26333 10275 26367
rect 10275 26333 10284 26367
rect 10232 26324 10284 26333
rect 10324 26324 10376 26376
rect 10968 26367 11020 26376
rect 10968 26333 10977 26367
rect 10977 26333 11011 26367
rect 11011 26333 11020 26367
rect 10968 26324 11020 26333
rect 11612 26324 11664 26376
rect 11980 26324 12032 26376
rect 12440 26324 12492 26376
rect 13360 26392 13412 26444
rect 12624 26324 12676 26376
rect 7104 26256 7156 26308
rect 8576 26256 8628 26308
rect 13360 26299 13412 26308
rect 13360 26265 13369 26299
rect 13369 26265 13403 26299
rect 13403 26265 13412 26299
rect 13360 26256 13412 26265
rect 6552 26188 6604 26240
rect 6828 26188 6880 26240
rect 9312 26188 9364 26240
rect 9956 26188 10008 26240
rect 4376 26086 4428 26138
rect 4440 26086 4492 26138
rect 4504 26086 4556 26138
rect 4568 26086 4620 26138
rect 4632 26086 4684 26138
rect 7803 26086 7855 26138
rect 7867 26086 7919 26138
rect 7931 26086 7983 26138
rect 7995 26086 8047 26138
rect 8059 26086 8111 26138
rect 11230 26086 11282 26138
rect 11294 26086 11346 26138
rect 11358 26086 11410 26138
rect 11422 26086 11474 26138
rect 11486 26086 11538 26138
rect 14657 26086 14709 26138
rect 14721 26086 14773 26138
rect 14785 26086 14837 26138
rect 14849 26086 14901 26138
rect 14913 26086 14965 26138
rect 3148 25984 3200 26036
rect 5816 25984 5868 26036
rect 8484 26027 8536 26036
rect 8484 25993 8493 26027
rect 8493 25993 8527 26027
rect 8527 25993 8536 26027
rect 8484 25984 8536 25993
rect 9220 25984 9272 26036
rect 10140 25984 10192 26036
rect 12256 25984 12308 26036
rect 4160 25916 4212 25968
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 3332 25848 3384 25900
rect 4252 25891 4304 25900
rect 4252 25857 4261 25891
rect 4261 25857 4295 25891
rect 4295 25857 4304 25891
rect 4252 25848 4304 25857
rect 4712 25848 4764 25900
rect 5356 25891 5408 25900
rect 5356 25857 5365 25891
rect 5365 25857 5399 25891
rect 5399 25857 5408 25891
rect 5356 25848 5408 25857
rect 6828 25891 6880 25900
rect 6828 25857 6837 25891
rect 6837 25857 6871 25891
rect 6871 25857 6880 25891
rect 6828 25848 6880 25857
rect 8668 25848 8720 25900
rect 10876 25891 10928 25900
rect 10876 25857 10885 25891
rect 10885 25857 10919 25891
rect 10919 25857 10928 25891
rect 10876 25848 10928 25857
rect 12164 25891 12216 25900
rect 12164 25857 12173 25891
rect 12173 25857 12207 25891
rect 12207 25857 12216 25891
rect 12164 25848 12216 25857
rect 11888 25780 11940 25832
rect 14188 25712 14240 25764
rect 1768 25687 1820 25696
rect 1768 25653 1777 25687
rect 1777 25653 1811 25687
rect 1811 25653 1820 25687
rect 1768 25644 1820 25653
rect 3240 25687 3292 25696
rect 3240 25653 3249 25687
rect 3249 25653 3283 25687
rect 3283 25653 3292 25687
rect 3240 25644 3292 25653
rect 4344 25644 4396 25696
rect 13728 25644 13780 25696
rect 2663 25542 2715 25594
rect 2727 25542 2779 25594
rect 2791 25542 2843 25594
rect 2855 25542 2907 25594
rect 2919 25542 2971 25594
rect 6090 25542 6142 25594
rect 6154 25542 6206 25594
rect 6218 25542 6270 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 9517 25542 9569 25594
rect 9581 25542 9633 25594
rect 9645 25542 9697 25594
rect 9709 25542 9761 25594
rect 9773 25542 9825 25594
rect 12944 25542 12996 25594
rect 13008 25542 13060 25594
rect 13072 25542 13124 25594
rect 13136 25542 13188 25594
rect 13200 25542 13252 25594
rect 2504 25440 2556 25492
rect 3056 25483 3108 25492
rect 3056 25449 3065 25483
rect 3065 25449 3099 25483
rect 3099 25449 3108 25483
rect 3056 25440 3108 25449
rect 3976 25440 4028 25492
rect 12716 25440 12768 25492
rect 12900 25372 12952 25424
rect 2228 25279 2280 25288
rect 2228 25245 2237 25279
rect 2237 25245 2271 25279
rect 2271 25245 2280 25279
rect 2228 25236 2280 25245
rect 3056 25236 3108 25288
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 4344 25279 4396 25288
rect 4344 25245 4353 25279
rect 4353 25245 4387 25279
rect 4387 25245 4396 25279
rect 4344 25236 4396 25245
rect 8760 25236 8812 25288
rect 11888 25279 11940 25288
rect 11888 25245 11897 25279
rect 11897 25245 11931 25279
rect 11931 25245 11940 25279
rect 11888 25236 11940 25245
rect 12164 25236 12216 25288
rect 13360 25279 13412 25288
rect 13360 25245 13369 25279
rect 13369 25245 13403 25279
rect 13403 25245 13412 25279
rect 13360 25236 13412 25245
rect 13636 25100 13688 25152
rect 4376 24998 4428 25050
rect 4440 24998 4492 25050
rect 4504 24998 4556 25050
rect 4568 24998 4620 25050
rect 4632 24998 4684 25050
rect 7803 24998 7855 25050
rect 7867 24998 7919 25050
rect 7931 24998 7983 25050
rect 7995 24998 8047 25050
rect 8059 24998 8111 25050
rect 11230 24998 11282 25050
rect 11294 24998 11346 25050
rect 11358 24998 11410 25050
rect 11422 24998 11474 25050
rect 11486 24998 11538 25050
rect 14657 24998 14709 25050
rect 14721 24998 14773 25050
rect 14785 24998 14837 25050
rect 14849 24998 14901 25050
rect 14913 24998 14965 25050
rect 1584 24760 1636 24812
rect 1952 24760 2004 24812
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 12808 24760 12860 24812
rect 3884 24692 3936 24744
rect 1860 24667 1912 24676
rect 1860 24633 1869 24667
rect 1869 24633 1903 24667
rect 1903 24633 1912 24667
rect 1860 24624 1912 24633
rect 2320 24624 2372 24676
rect 13268 24667 13320 24676
rect 13268 24633 13277 24667
rect 13277 24633 13311 24667
rect 13311 24633 13320 24667
rect 13268 24624 13320 24633
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 2663 24454 2715 24506
rect 2727 24454 2779 24506
rect 2791 24454 2843 24506
rect 2855 24454 2907 24506
rect 2919 24454 2971 24506
rect 6090 24454 6142 24506
rect 6154 24454 6206 24506
rect 6218 24454 6270 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 9517 24454 9569 24506
rect 9581 24454 9633 24506
rect 9645 24454 9697 24506
rect 9709 24454 9761 24506
rect 9773 24454 9825 24506
rect 12944 24454 12996 24506
rect 13008 24454 13060 24506
rect 13072 24454 13124 24506
rect 13136 24454 13188 24506
rect 13200 24454 13252 24506
rect 1676 24352 1728 24404
rect 13452 24352 13504 24404
rect 1768 24148 1820 24200
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 4376 23910 4428 23962
rect 4440 23910 4492 23962
rect 4504 23910 4556 23962
rect 4568 23910 4620 23962
rect 4632 23910 4684 23962
rect 7803 23910 7855 23962
rect 7867 23910 7919 23962
rect 7931 23910 7983 23962
rect 7995 23910 8047 23962
rect 8059 23910 8111 23962
rect 11230 23910 11282 23962
rect 11294 23910 11346 23962
rect 11358 23910 11410 23962
rect 11422 23910 11474 23962
rect 11486 23910 11538 23962
rect 14657 23910 14709 23962
rect 14721 23910 14773 23962
rect 14785 23910 14837 23962
rect 14849 23910 14901 23962
rect 14913 23910 14965 23962
rect 13912 23808 13964 23860
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 2663 23366 2715 23418
rect 2727 23366 2779 23418
rect 2791 23366 2843 23418
rect 2855 23366 2907 23418
rect 2919 23366 2971 23418
rect 6090 23366 6142 23418
rect 6154 23366 6206 23418
rect 6218 23366 6270 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 9517 23366 9569 23418
rect 9581 23366 9633 23418
rect 9645 23366 9697 23418
rect 9709 23366 9761 23418
rect 9773 23366 9825 23418
rect 12944 23366 12996 23418
rect 13008 23366 13060 23418
rect 13072 23366 13124 23418
rect 13136 23366 13188 23418
rect 13200 23366 13252 23418
rect 4376 22822 4428 22874
rect 4440 22822 4492 22874
rect 4504 22822 4556 22874
rect 4568 22822 4620 22874
rect 4632 22822 4684 22874
rect 7803 22822 7855 22874
rect 7867 22822 7919 22874
rect 7931 22822 7983 22874
rect 7995 22822 8047 22874
rect 8059 22822 8111 22874
rect 11230 22822 11282 22874
rect 11294 22822 11346 22874
rect 11358 22822 11410 22874
rect 11422 22822 11474 22874
rect 11486 22822 11538 22874
rect 14657 22822 14709 22874
rect 14721 22822 14773 22874
rect 14785 22822 14837 22874
rect 14849 22822 14901 22874
rect 14913 22822 14965 22874
rect 2663 22278 2715 22330
rect 2727 22278 2779 22330
rect 2791 22278 2843 22330
rect 2855 22278 2907 22330
rect 2919 22278 2971 22330
rect 6090 22278 6142 22330
rect 6154 22278 6206 22330
rect 6218 22278 6270 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 9517 22278 9569 22330
rect 9581 22278 9633 22330
rect 9645 22278 9697 22330
rect 9709 22278 9761 22330
rect 9773 22278 9825 22330
rect 12944 22278 12996 22330
rect 13008 22278 13060 22330
rect 13072 22278 13124 22330
rect 13136 22278 13188 22330
rect 13200 22278 13252 22330
rect 5448 21972 5500 22024
rect 3424 21904 3476 21956
rect 3332 21836 3384 21888
rect 4376 21734 4428 21786
rect 4440 21734 4492 21786
rect 4504 21734 4556 21786
rect 4568 21734 4620 21786
rect 4632 21734 4684 21786
rect 7803 21734 7855 21786
rect 7867 21734 7919 21786
rect 7931 21734 7983 21786
rect 7995 21734 8047 21786
rect 8059 21734 8111 21786
rect 11230 21734 11282 21786
rect 11294 21734 11346 21786
rect 11358 21734 11410 21786
rect 11422 21734 11474 21786
rect 11486 21734 11538 21786
rect 14657 21734 14709 21786
rect 14721 21734 14773 21786
rect 14785 21734 14837 21786
rect 14849 21734 14901 21786
rect 14913 21734 14965 21786
rect 5356 21632 5408 21684
rect 4160 21496 4212 21548
rect 4344 21539 4396 21548
rect 4344 21505 4378 21539
rect 4378 21505 4396 21539
rect 4344 21496 4396 21505
rect 2663 21190 2715 21242
rect 2727 21190 2779 21242
rect 2791 21190 2843 21242
rect 2855 21190 2907 21242
rect 2919 21190 2971 21242
rect 6090 21190 6142 21242
rect 6154 21190 6206 21242
rect 6218 21190 6270 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 9517 21190 9569 21242
rect 9581 21190 9633 21242
rect 9645 21190 9697 21242
rect 9709 21190 9761 21242
rect 9773 21190 9825 21242
rect 12944 21190 12996 21242
rect 13008 21190 13060 21242
rect 13072 21190 13124 21242
rect 13136 21190 13188 21242
rect 13200 21190 13252 21242
rect 3424 21131 3476 21140
rect 3424 21097 3433 21131
rect 3433 21097 3467 21131
rect 3467 21097 3476 21131
rect 3424 21088 3476 21097
rect 4344 21131 4396 21140
rect 4344 21097 4353 21131
rect 4353 21097 4387 21131
rect 4387 21097 4396 21131
rect 4344 21088 4396 21097
rect 4620 20884 4672 20936
rect 5724 21088 5776 21140
rect 6644 21088 6696 21140
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 4896 20884 4948 20936
rect 5448 20884 5500 20936
rect 6184 20884 6236 20936
rect 7196 20927 7248 20936
rect 7196 20893 7205 20927
rect 7205 20893 7239 20927
rect 7239 20893 7248 20927
rect 7196 20884 7248 20893
rect 5540 20748 5592 20800
rect 9128 20816 9180 20868
rect 4376 20646 4428 20698
rect 4440 20646 4492 20698
rect 4504 20646 4556 20698
rect 4568 20646 4620 20698
rect 4632 20646 4684 20698
rect 7803 20646 7855 20698
rect 7867 20646 7919 20698
rect 7931 20646 7983 20698
rect 7995 20646 8047 20698
rect 8059 20646 8111 20698
rect 11230 20646 11282 20698
rect 11294 20646 11346 20698
rect 11358 20646 11410 20698
rect 11422 20646 11474 20698
rect 11486 20646 11538 20698
rect 14657 20646 14709 20698
rect 14721 20646 14773 20698
rect 14785 20646 14837 20698
rect 14849 20646 14901 20698
rect 14913 20646 14965 20698
rect 3148 20544 3200 20596
rect 4712 20544 4764 20596
rect 6552 20544 6604 20596
rect 12808 20544 12860 20596
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 5448 20476 5500 20528
rect 8300 20476 8352 20528
rect 4160 20408 4212 20417
rect 5632 20408 5684 20460
rect 6184 20408 6236 20460
rect 5816 20340 5868 20392
rect 4620 20204 4672 20256
rect 7196 20340 7248 20392
rect 2663 20102 2715 20154
rect 2727 20102 2779 20154
rect 2791 20102 2843 20154
rect 2855 20102 2907 20154
rect 2919 20102 2971 20154
rect 6090 20102 6142 20154
rect 6154 20102 6206 20154
rect 6218 20102 6270 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 9517 20102 9569 20154
rect 9581 20102 9633 20154
rect 9645 20102 9697 20154
rect 9709 20102 9761 20154
rect 9773 20102 9825 20154
rect 12944 20102 12996 20154
rect 13008 20102 13060 20154
rect 13072 20102 13124 20154
rect 13136 20102 13188 20154
rect 13200 20102 13252 20154
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 5540 20000 5592 20052
rect 7564 20000 7616 20052
rect 12440 20000 12492 20052
rect 4160 19932 4212 19984
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 5448 19796 5500 19848
rect 6920 19796 6972 19848
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 6736 19728 6788 19780
rect 8852 19728 8904 19780
rect 4252 19660 4304 19712
rect 5908 19660 5960 19712
rect 4376 19558 4428 19610
rect 4440 19558 4492 19610
rect 4504 19558 4556 19610
rect 4568 19558 4620 19610
rect 4632 19558 4684 19610
rect 7803 19558 7855 19610
rect 7867 19558 7919 19610
rect 7931 19558 7983 19610
rect 7995 19558 8047 19610
rect 8059 19558 8111 19610
rect 11230 19558 11282 19610
rect 11294 19558 11346 19610
rect 11358 19558 11410 19610
rect 11422 19558 11474 19610
rect 11486 19558 11538 19610
rect 14657 19558 14709 19610
rect 14721 19558 14773 19610
rect 14785 19558 14837 19610
rect 14849 19558 14901 19610
rect 14913 19558 14965 19610
rect 4804 19456 4856 19508
rect 4896 19456 4948 19508
rect 5816 19456 5868 19508
rect 6000 19456 6052 19508
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 5724 19431 5776 19440
rect 5724 19397 5742 19431
rect 5742 19397 5776 19431
rect 5724 19388 5776 19397
rect 6920 19320 6972 19372
rect 9036 19320 9088 19372
rect 2663 19014 2715 19066
rect 2727 19014 2779 19066
rect 2791 19014 2843 19066
rect 2855 19014 2907 19066
rect 2919 19014 2971 19066
rect 6090 19014 6142 19066
rect 6154 19014 6206 19066
rect 6218 19014 6270 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 9517 19014 9569 19066
rect 9581 19014 9633 19066
rect 9645 19014 9697 19066
rect 9709 19014 9761 19066
rect 9773 19014 9825 19066
rect 12944 19014 12996 19066
rect 13008 19014 13060 19066
rect 13072 19014 13124 19066
rect 13136 19014 13188 19066
rect 13200 19014 13252 19066
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 5540 18708 5592 18760
rect 5356 18640 5408 18692
rect 4376 18470 4428 18522
rect 4440 18470 4492 18522
rect 4504 18470 4556 18522
rect 4568 18470 4620 18522
rect 4632 18470 4684 18522
rect 7803 18470 7855 18522
rect 7867 18470 7919 18522
rect 7931 18470 7983 18522
rect 7995 18470 8047 18522
rect 8059 18470 8111 18522
rect 11230 18470 11282 18522
rect 11294 18470 11346 18522
rect 11358 18470 11410 18522
rect 11422 18470 11474 18522
rect 11486 18470 11538 18522
rect 14657 18470 14709 18522
rect 14721 18470 14773 18522
rect 14785 18470 14837 18522
rect 14849 18470 14901 18522
rect 14913 18470 14965 18522
rect 5908 18300 5960 18352
rect 5724 18232 5776 18284
rect 6828 18275 6880 18284
rect 6828 18241 6837 18275
rect 6837 18241 6871 18275
rect 6871 18241 6880 18275
rect 6828 18232 6880 18241
rect 7012 18071 7064 18080
rect 7012 18037 7021 18071
rect 7021 18037 7055 18071
rect 7055 18037 7064 18071
rect 7012 18028 7064 18037
rect 2663 17926 2715 17978
rect 2727 17926 2779 17978
rect 2791 17926 2843 17978
rect 2855 17926 2907 17978
rect 2919 17926 2971 17978
rect 6090 17926 6142 17978
rect 6154 17926 6206 17978
rect 6218 17926 6270 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 9517 17926 9569 17978
rect 9581 17926 9633 17978
rect 9645 17926 9697 17978
rect 9709 17926 9761 17978
rect 9773 17926 9825 17978
rect 12944 17926 12996 17978
rect 13008 17926 13060 17978
rect 13072 17926 13124 17978
rect 13136 17926 13188 17978
rect 13200 17926 13252 17978
rect 4252 17824 4304 17876
rect 5632 17824 5684 17876
rect 11612 17824 11664 17876
rect 4160 17620 4212 17672
rect 4712 17620 4764 17672
rect 5172 17620 5224 17672
rect 5632 17620 5684 17672
rect 5816 17756 5868 17808
rect 6092 17756 6144 17808
rect 5908 17731 5960 17740
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 6920 17620 6972 17672
rect 4896 17484 4948 17536
rect 9220 17552 9272 17604
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 3056 17280 3108 17332
rect 8944 17280 8996 17332
rect 4344 17144 4396 17196
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 6920 17212 6972 17264
rect 7012 17212 7064 17264
rect 4160 16940 4212 16992
rect 5632 16940 5684 16992
rect 5724 16940 5776 16992
rect 6092 16940 6144 16992
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 4344 16779 4396 16788
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 6000 16668 6052 16720
rect 5632 16600 5684 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 9312 16575 9364 16584
rect 9312 16541 9321 16575
rect 9321 16541 9355 16575
rect 9355 16541 9364 16575
rect 9312 16532 9364 16541
rect 5632 16464 5684 16516
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 12164 16192 12216 16244
rect 4712 16056 4764 16108
rect 5908 16124 5960 16176
rect 6736 16124 6788 16176
rect 5816 16056 5868 16108
rect 6920 16056 6972 16108
rect 8392 16056 8444 16108
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5080 15852 5132 15904
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 5540 15648 5592 15700
rect 4804 15580 4856 15632
rect 4896 15512 4948 15564
rect 5080 15512 5132 15564
rect 7472 15580 7524 15632
rect 5816 15444 5868 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 9404 15444 9456 15496
rect 5632 15376 5684 15428
rect 4896 15308 4948 15360
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 4252 15104 4304 15156
rect 8392 15147 8444 15156
rect 8392 15113 8401 15147
rect 8401 15113 8435 15147
rect 8435 15113 8444 15147
rect 8392 15104 8444 15113
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9036 15104 9088 15113
rect 4896 15079 4948 15088
rect 4896 15045 4914 15079
rect 4914 15045 4948 15079
rect 4896 15036 4948 15045
rect 5540 14968 5592 15020
rect 6920 15036 6972 15088
rect 7380 14968 7432 15020
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 8668 14832 8720 14884
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 7104 14560 7156 14612
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 8300 14603 8352 14612
rect 8300 14569 8309 14603
rect 8309 14569 8343 14603
rect 8343 14569 8352 14603
rect 8300 14560 8352 14569
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 4712 14424 4764 14476
rect 6736 14424 6788 14476
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 5264 14356 5316 14408
rect 7472 14356 7524 14408
rect 8484 14399 8536 14408
rect 6828 14288 6880 14340
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4804 14220 4856 14272
rect 7656 14220 7708 14272
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 9404 14356 9456 14408
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 3884 14059 3936 14068
rect 3884 14025 3893 14059
rect 3893 14025 3927 14059
rect 3927 14025 3936 14059
rect 3884 14016 3936 14025
rect 6828 14016 6880 14068
rect 8852 14059 8904 14068
rect 4160 13948 4212 14000
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 10324 13948 10376 14000
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 6000 13923 6052 13932
rect 6000 13889 6009 13923
rect 6009 13889 6043 13923
rect 6043 13889 6052 13923
rect 6000 13880 6052 13889
rect 8760 13880 8812 13932
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 4804 13515 4856 13524
rect 4804 13481 4813 13515
rect 4813 13481 4847 13515
rect 4847 13481 4856 13515
rect 4804 13472 4856 13481
rect 5724 13472 5776 13524
rect 8576 13472 8628 13524
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 5172 13404 5224 13456
rect 6552 13268 6604 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 8668 13268 8720 13320
rect 9772 13268 9824 13320
rect 6644 13200 6696 13252
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 5080 12971 5132 12980
rect 5080 12937 5089 12971
rect 5089 12937 5123 12971
rect 5123 12937 5132 12971
rect 5080 12928 5132 12937
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 9220 12928 9272 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 8852 12792 8904 12844
rect 9312 12792 9364 12844
rect 10048 12792 10100 12844
rect 4804 12724 4856 12776
rect 5448 12656 5500 12708
rect 7656 12724 7708 12776
rect 8208 12724 8260 12776
rect 9404 12656 9456 12708
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 4712 12384 4764 12436
rect 5540 12384 5592 12436
rect 9036 12384 9088 12436
rect 4896 12316 4948 12368
rect 7564 12180 7616 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 5908 12044 5960 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 4804 11840 4856 11892
rect 7564 11840 7616 11892
rect 8760 11840 8812 11892
rect 4252 11704 4304 11756
rect 4988 11704 5040 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 6460 11704 6512 11756
rect 7012 11704 7064 11756
rect 8576 11704 8628 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 5724 11568 5776 11620
rect 6736 11568 6788 11620
rect 10876 11568 10928 11620
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 5908 11296 5960 11348
rect 5724 11160 5776 11212
rect 6920 11228 6972 11280
rect 7196 11160 7248 11212
rect 6460 11092 6512 11144
rect 5172 11024 5224 11076
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 9220 10752 9272 10804
rect 4160 10616 4212 10668
rect 5264 10684 5316 10736
rect 7104 10684 7156 10736
rect 4252 10548 4304 10600
rect 7564 10616 7616 10668
rect 9128 10616 9180 10668
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 6920 10480 6972 10532
rect 8576 10523 8628 10532
rect 8576 10489 8585 10523
rect 8585 10489 8619 10523
rect 8619 10489 8628 10523
rect 8576 10480 8628 10489
rect 6460 10412 6512 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 6460 10115 6512 10124
rect 6460 10081 6469 10115
rect 6469 10081 6503 10115
rect 6503 10081 6512 10115
rect 6460 10072 6512 10081
rect 5356 10004 5408 10056
rect 7012 10004 7064 10056
rect 7656 9936 7708 9988
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 13452 9936 13504 9988
rect 8392 9868 8444 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 7656 9664 7708 9716
rect 4068 9528 4120 9580
rect 4528 9528 4580 9580
rect 7196 9528 7248 9580
rect 7472 9528 7524 9580
rect 5172 9392 5224 9444
rect 6644 9392 6696 9444
rect 6920 9392 6972 9444
rect 7288 9460 7340 9512
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 6828 9120 6880 9172
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 7380 9052 7432 9104
rect 9036 8984 9088 9036
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 7288 8916 7340 8968
rect 7472 8916 7524 8968
rect 8300 8916 8352 8968
rect 9128 8848 9180 8900
rect 5908 8823 5960 8832
rect 5908 8789 5917 8823
rect 5917 8789 5951 8823
rect 5951 8789 5960 8823
rect 5908 8780 5960 8789
rect 7288 8823 7340 8832
rect 7288 8789 7297 8823
rect 7297 8789 7331 8823
rect 7331 8789 7340 8823
rect 7288 8780 7340 8789
rect 8760 8780 8812 8832
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 5816 8576 5868 8628
rect 9128 8619 9180 8628
rect 6920 8508 6972 8560
rect 7380 8508 7432 8560
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 9864 8508 9916 8560
rect 6736 8440 6788 8492
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 8760 8440 8812 8492
rect 9404 8372 9456 8424
rect 5724 8304 5776 8356
rect 6828 8304 6880 8356
rect 7012 8304 7064 8356
rect 8300 8304 8352 8356
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 8944 8304 8996 8313
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 4252 8032 4304 8084
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7288 8032 7340 8084
rect 8944 8032 8996 8084
rect 9404 8032 9456 8084
rect 9036 7964 9088 8016
rect 5172 7896 5224 7948
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5540 7828 5592 7880
rect 8392 7896 8444 7948
rect 8300 7828 8352 7880
rect 7656 7760 7708 7812
rect 9864 7828 9916 7880
rect 8300 7692 8352 7744
rect 8576 7692 8628 7744
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 4068 7488 4120 7540
rect 4804 7488 4856 7540
rect 5356 7488 5408 7540
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 5632 7420 5684 7472
rect 8300 7420 8352 7472
rect 8760 7420 8812 7472
rect 4620 7352 4672 7404
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 6644 7352 6696 7404
rect 5172 7284 5224 7336
rect 6000 7284 6052 7336
rect 14096 7352 14148 7404
rect 7656 7216 7708 7268
rect 9220 7216 9272 7268
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 5264 6808 5316 6860
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 9404 6808 9456 6860
rect 4160 6672 4212 6724
rect 4804 6740 4856 6792
rect 5172 6740 5224 6792
rect 6736 6740 6788 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 9220 6740 9272 6792
rect 3792 6604 3844 6656
rect 4620 6604 4672 6656
rect 5908 6672 5960 6724
rect 6644 6604 6696 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 8852 6604 8904 6656
rect 12440 6604 12492 6656
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 3792 6375 3844 6384
rect 3792 6341 3801 6375
rect 3801 6341 3835 6375
rect 3835 6341 3844 6375
rect 3792 6332 3844 6341
rect 4712 6400 4764 6452
rect 5540 6400 5592 6452
rect 6920 6400 6972 6452
rect 8484 6400 8536 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 4804 6332 4856 6384
rect 8392 6332 8444 6384
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 6736 6307 6788 6316
rect 5816 6264 5868 6273
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 6828 6264 6880 6316
rect 10968 6264 11020 6316
rect 5540 6128 5592 6180
rect 6000 6171 6052 6180
rect 6000 6137 6009 6171
rect 6009 6137 6043 6171
rect 6043 6137 6052 6171
rect 6000 6128 6052 6137
rect 4252 6060 4304 6112
rect 5080 6060 5132 6112
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 7012 6060 7064 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 4804 5899 4856 5908
rect 4804 5865 4813 5899
rect 4813 5865 4847 5899
rect 4847 5865 4856 5899
rect 4804 5856 4856 5865
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6828 5856 6880 5908
rect 5172 5720 5224 5772
rect 5632 5720 5684 5772
rect 4160 5584 4212 5636
rect 5264 5652 5316 5704
rect 7288 5695 7340 5704
rect 5356 5584 5408 5636
rect 5540 5516 5592 5568
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 8300 5788 8352 5840
rect 8576 5831 8628 5840
rect 8576 5797 8585 5831
rect 8585 5797 8619 5831
rect 8619 5797 8628 5831
rect 8576 5788 8628 5797
rect 8300 5652 8352 5704
rect 9864 5652 9916 5704
rect 6644 5516 6696 5568
rect 8392 5516 8444 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 5724 5312 5776 5364
rect 5632 5287 5684 5296
rect 5632 5253 5641 5287
rect 5641 5253 5675 5287
rect 5675 5253 5684 5287
rect 5632 5244 5684 5253
rect 5724 5108 5776 5160
rect 6644 5312 6696 5364
rect 6920 5287 6972 5296
rect 6920 5253 6929 5287
rect 6929 5253 6963 5287
rect 6963 5253 6972 5287
rect 6920 5244 6972 5253
rect 7288 5176 7340 5228
rect 6828 5108 6880 5160
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 6460 4972 6512 5024
rect 7012 5040 7064 5092
rect 7104 5015 7156 5024
rect 7104 4981 7113 5015
rect 7113 4981 7147 5015
rect 7147 4981 7156 5015
rect 7104 4972 7156 4981
rect 7472 4972 7524 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 5540 4768 5592 4820
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 6920 4768 6972 4820
rect 8208 4768 8260 4820
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4988 4564 5040 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5632 4564 5684 4616
rect 8392 4632 8444 4684
rect 9220 4632 9272 4684
rect 6460 4564 6512 4616
rect 7380 4564 7432 4616
rect 8300 4564 8352 4616
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 5356 4428 5408 4437
rect 8392 4496 8444 4548
rect 10784 4496 10836 4548
rect 6644 4428 6696 4480
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 6644 4224 6696 4276
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 8300 4156 8352 4208
rect 9864 4156 9916 4208
rect 4068 4088 4120 4140
rect 4252 4131 4304 4140
rect 4252 4097 4286 4131
rect 4286 4097 4304 4131
rect 4252 4088 4304 4097
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6644 4088 6696 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 7472 4131 7524 4140
rect 6828 4088 6880 4097
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 8392 4063 8444 4072
rect 5540 3952 5592 4004
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 10048 3952 10100 4004
rect 4344 3884 4396 3936
rect 5264 3884 5316 3936
rect 7380 3884 7432 3936
rect 9036 3884 9088 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 3056 3680 3108 3732
rect 5448 3680 5500 3732
rect 4896 3612 4948 3664
rect 6460 3680 6512 3732
rect 8300 3680 8352 3732
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 6736 3544 6788 3596
rect 7380 3519 7432 3528
rect 7380 3485 7414 3519
rect 7414 3485 7432 3519
rect 7380 3476 7432 3485
rect 4160 3408 4212 3460
rect 6552 3408 6604 3460
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 14004 3340 14056 3392
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 4252 3136 4304 3188
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6460 3136 6512 3188
rect 7564 3136 7616 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 5356 3068 5408 3120
rect 756 3000 808 3052
rect 4068 3000 4120 3052
rect 8392 3000 8444 3052
rect 7012 2932 7064 2984
rect 7472 2932 7524 2984
rect 14004 3000 14056 3052
rect 15108 2932 15160 2984
rect 4436 2864 4488 2916
rect 7380 2864 7432 2916
rect 3240 2796 3292 2848
rect 5816 2796 5868 2848
rect 8484 2796 8536 2848
rect 10692 2839 10744 2848
rect 10692 2805 10701 2839
rect 10701 2805 10735 2839
rect 10735 2805 10744 2839
rect 10692 2796 10744 2805
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 4160 2592 4212 2644
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 7196 2592 7248 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 9864 2592 9916 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 10968 2592 11020 2644
rect 12440 2592 12492 2644
rect 4620 2567 4672 2576
rect 4620 2533 4629 2567
rect 4629 2533 4663 2567
rect 4663 2533 4672 2567
rect 4620 2524 4672 2533
rect 7288 2524 7340 2576
rect 4712 2456 4764 2508
rect 7012 2456 7064 2508
rect 1860 2388 1912 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4068 2388 4120 2440
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 5080 2388 5132 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6276 2388 6328 2440
rect 7104 2388 7156 2440
rect 7380 2388 7432 2440
rect 8484 2388 8536 2440
rect 4252 2320 4304 2372
rect 10692 2388 10744 2440
rect 11796 2388 11848 2440
rect 12900 2388 12952 2440
rect 9588 2252 9640 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
<< metal2 >>
rect 1766 29322 1822 30000
rect 2042 29322 2098 30000
rect 1688 29294 1822 29322
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 24818 1624 25842
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1688 24410 1716 29294
rect 1766 29200 1822 29294
rect 1872 29294 2098 29322
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1780 24206 1808 25638
rect 1872 24682 1900 29294
rect 2042 29200 2098 29294
rect 2318 29200 2374 30000
rect 2594 29322 2650 30000
rect 2516 29294 2650 29322
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1964 26790 1992 27406
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 1952 26512 2004 26518
rect 1952 26454 2004 26460
rect 1964 24818 1992 26454
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2044 26308 2096 26314
rect 2044 26250 2096 26256
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 2056 20058 2084 26250
rect 2240 25294 2268 26318
rect 2228 25288 2280 25294
rect 2228 25230 2280 25236
rect 2332 24682 2360 29200
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 2424 26314 2452 27406
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 2516 25498 2544 29294
rect 2594 29200 2650 29294
rect 2870 29322 2926 30000
rect 2870 29294 3096 29322
rect 2870 29200 2926 29294
rect 2663 27772 2971 27781
rect 2663 27770 2669 27772
rect 2725 27770 2749 27772
rect 2805 27770 2829 27772
rect 2885 27770 2909 27772
rect 2965 27770 2971 27772
rect 2725 27718 2727 27770
rect 2907 27718 2909 27770
rect 2663 27716 2669 27718
rect 2725 27716 2749 27718
rect 2805 27716 2829 27718
rect 2885 27716 2909 27718
rect 2965 27716 2971 27718
rect 2663 27707 2971 27716
rect 2663 26684 2971 26693
rect 2663 26682 2669 26684
rect 2725 26682 2749 26684
rect 2805 26682 2829 26684
rect 2885 26682 2909 26684
rect 2965 26682 2971 26684
rect 2725 26630 2727 26682
rect 2907 26630 2909 26682
rect 2663 26628 2669 26630
rect 2725 26628 2749 26630
rect 2805 26628 2829 26630
rect 2885 26628 2909 26630
rect 2965 26628 2971 26630
rect 2663 26619 2971 26628
rect 2663 25596 2971 25605
rect 2663 25594 2669 25596
rect 2725 25594 2749 25596
rect 2805 25594 2829 25596
rect 2885 25594 2909 25596
rect 2965 25594 2971 25596
rect 2725 25542 2727 25594
rect 2907 25542 2909 25594
rect 2663 25540 2669 25542
rect 2725 25540 2749 25542
rect 2805 25540 2829 25542
rect 2885 25540 2909 25542
rect 2965 25540 2971 25542
rect 2663 25531 2971 25540
rect 3068 25498 3096 29294
rect 3146 29200 3202 30000
rect 3422 29200 3478 30000
rect 3698 29322 3754 30000
rect 3528 29294 3754 29322
rect 3160 26042 3188 29200
rect 3240 26920 3292 26926
rect 3240 26862 3292 26868
rect 3252 26382 3280 26862
rect 3436 26586 3464 29200
rect 3528 27130 3556 29294
rect 3698 29200 3754 29294
rect 3974 29200 4030 30000
rect 4250 29322 4306 30000
rect 4172 29294 4306 29322
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3700 26988 3752 26994
rect 3700 26930 3752 26936
rect 3712 26586 3740 26930
rect 3424 26580 3476 26586
rect 3424 26522 3476 26528
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3148 26036 3200 26042
rect 3148 25978 3200 25984
rect 3252 25786 3280 26318
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 3160 25758 3280 25786
rect 2504 25492 2556 25498
rect 2504 25434 2556 25440
rect 3056 25492 3108 25498
rect 3056 25434 3108 25440
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 2320 24676 2372 24682
rect 2320 24618 2372 24624
rect 2663 24508 2971 24517
rect 2663 24506 2669 24508
rect 2725 24506 2749 24508
rect 2805 24506 2829 24508
rect 2885 24506 2909 24508
rect 2965 24506 2971 24508
rect 2725 24454 2727 24506
rect 2907 24454 2909 24506
rect 2663 24452 2669 24454
rect 2725 24452 2749 24454
rect 2805 24452 2829 24454
rect 2885 24452 2909 24454
rect 2965 24452 2971 24454
rect 2663 24443 2971 24452
rect 2663 23420 2971 23429
rect 2663 23418 2669 23420
rect 2725 23418 2749 23420
rect 2805 23418 2829 23420
rect 2885 23418 2909 23420
rect 2965 23418 2971 23420
rect 2725 23366 2727 23418
rect 2907 23366 2909 23418
rect 2663 23364 2669 23366
rect 2725 23364 2749 23366
rect 2805 23364 2829 23366
rect 2885 23364 2909 23366
rect 2965 23364 2971 23366
rect 2663 23355 2971 23364
rect 2663 22332 2971 22341
rect 2663 22330 2669 22332
rect 2725 22330 2749 22332
rect 2805 22330 2829 22332
rect 2885 22330 2909 22332
rect 2965 22330 2971 22332
rect 2725 22278 2727 22330
rect 2907 22278 2909 22330
rect 2663 22276 2669 22278
rect 2725 22276 2749 22278
rect 2805 22276 2829 22278
rect 2885 22276 2909 22278
rect 2965 22276 2971 22278
rect 2663 22267 2971 22276
rect 2663 21244 2971 21253
rect 2663 21242 2669 21244
rect 2725 21242 2749 21244
rect 2805 21242 2829 21244
rect 2885 21242 2909 21244
rect 2965 21242 2971 21244
rect 2725 21190 2727 21242
rect 2907 21190 2909 21242
rect 2663 21188 2669 21190
rect 2725 21188 2749 21190
rect 2805 21188 2829 21190
rect 2885 21188 2909 21190
rect 2965 21188 2971 21190
rect 2663 21179 2971 21188
rect 2663 20156 2971 20165
rect 2663 20154 2669 20156
rect 2725 20154 2749 20156
rect 2805 20154 2829 20156
rect 2885 20154 2909 20156
rect 2965 20154 2971 20156
rect 2725 20102 2727 20154
rect 2907 20102 2909 20154
rect 2663 20100 2669 20102
rect 2725 20100 2749 20102
rect 2805 20100 2829 20102
rect 2885 20100 2909 20102
rect 2965 20100 2971 20102
rect 2663 20091 2971 20100
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2663 19068 2971 19077
rect 2663 19066 2669 19068
rect 2725 19066 2749 19068
rect 2805 19066 2829 19068
rect 2885 19066 2909 19068
rect 2965 19066 2971 19068
rect 2725 19014 2727 19066
rect 2907 19014 2909 19066
rect 2663 19012 2669 19014
rect 2725 19012 2749 19014
rect 2805 19012 2829 19014
rect 2885 19012 2909 19014
rect 2965 19012 2971 19014
rect 2663 19003 2971 19012
rect 2663 17980 2971 17989
rect 2663 17978 2669 17980
rect 2725 17978 2749 17980
rect 2805 17978 2829 17980
rect 2885 17978 2909 17980
rect 2965 17978 2971 17980
rect 2725 17926 2727 17978
rect 2907 17926 2909 17978
rect 2663 17924 2669 17926
rect 2725 17924 2749 17926
rect 2805 17924 2829 17926
rect 2885 17924 2909 17926
rect 2965 17924 2971 17926
rect 2663 17915 2971 17924
rect 3068 17338 3096 25230
rect 3160 20602 3188 25758
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3252 25294 3280 25638
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3344 21894 3372 25842
rect 3988 25498 4016 29200
rect 4172 27554 4200 29294
rect 4250 29200 4306 29294
rect 4526 29200 4582 30000
rect 4802 29322 4858 30000
rect 4632 29294 4858 29322
rect 4080 27526 4200 27554
rect 4080 27402 4108 27526
rect 4540 27418 4568 29200
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 4264 27390 4568 27418
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 25974 4200 26930
rect 4264 26858 4292 27390
rect 4632 27334 4660 29294
rect 4802 29200 4858 29294
rect 5078 29200 5134 30000
rect 5354 29200 5410 30000
rect 5630 29200 5686 30000
rect 5906 29322 5962 30000
rect 6182 29322 6238 30000
rect 5736 29294 5962 29322
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4376 27228 4684 27237
rect 4376 27226 4382 27228
rect 4438 27226 4462 27228
rect 4518 27226 4542 27228
rect 4598 27226 4622 27228
rect 4678 27226 4684 27228
rect 4438 27174 4440 27226
rect 4620 27174 4622 27226
rect 4376 27172 4382 27174
rect 4438 27172 4462 27174
rect 4518 27172 4542 27174
rect 4598 27172 4622 27174
rect 4678 27172 4684 27174
rect 4376 27163 4684 27172
rect 5092 27062 5120 29200
rect 5368 27538 5396 29200
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5080 27056 5132 27062
rect 5080 26998 5132 27004
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4252 26852 4304 26858
rect 4252 26794 4304 26800
rect 4540 26518 4568 26930
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4376 26140 4684 26149
rect 4376 26138 4382 26140
rect 4438 26138 4462 26140
rect 4518 26138 4542 26140
rect 4598 26138 4622 26140
rect 4678 26138 4684 26140
rect 4438 26086 4440 26138
rect 4620 26086 4622 26138
rect 4376 26084 4382 26086
rect 4438 26084 4462 26086
rect 4518 26084 4542 26086
rect 4598 26084 4622 26086
rect 4678 26084 4684 26086
rect 4376 26075 4684 26084
rect 4160 25968 4212 25974
rect 4160 25910 4212 25916
rect 4724 25906 4752 26726
rect 5184 26382 5212 27406
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 5264 26988 5316 26994
rect 5264 26930 5316 26936
rect 5276 26586 5304 26930
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 4252 25900 4304 25906
rect 4252 25842 4304 25848
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3424 21956 3476 21962
rect 3424 21898 3476 21904
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3436 21146 3464 21898
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 3896 14074 3924 24686
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4172 20466 4200 21490
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4172 19990 4200 20402
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4264 19836 4292 25842
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 4356 25294 4384 25638
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4376 25052 4684 25061
rect 4376 25050 4382 25052
rect 4438 25050 4462 25052
rect 4518 25050 4542 25052
rect 4598 25050 4622 25052
rect 4678 25050 4684 25052
rect 4438 24998 4440 25050
rect 4620 24998 4622 25050
rect 4376 24996 4382 24998
rect 4438 24996 4462 24998
rect 4518 24996 4542 24998
rect 4598 24996 4622 24998
rect 4678 24996 4684 24998
rect 4376 24987 4684 24996
rect 4376 23964 4684 23973
rect 4376 23962 4382 23964
rect 4438 23962 4462 23964
rect 4518 23962 4542 23964
rect 4598 23962 4622 23964
rect 4678 23962 4684 23964
rect 4438 23910 4440 23962
rect 4620 23910 4622 23962
rect 4376 23908 4382 23910
rect 4438 23908 4462 23910
rect 4518 23908 4542 23910
rect 4598 23908 4622 23910
rect 4678 23908 4684 23910
rect 4376 23899 4684 23908
rect 4376 22876 4684 22885
rect 4376 22874 4382 22876
rect 4438 22874 4462 22876
rect 4518 22874 4542 22876
rect 4598 22874 4622 22876
rect 4678 22874 4684 22876
rect 4438 22822 4440 22874
rect 4620 22822 4622 22874
rect 4376 22820 4382 22822
rect 4438 22820 4462 22822
rect 4518 22820 4542 22822
rect 4598 22820 4622 22822
rect 4678 22820 4684 22822
rect 4376 22811 4684 22820
rect 4376 21788 4684 21797
rect 4376 21786 4382 21788
rect 4438 21786 4462 21788
rect 4518 21786 4542 21788
rect 4598 21786 4622 21788
rect 4678 21786 4684 21788
rect 4438 21734 4440 21786
rect 4620 21734 4622 21786
rect 4376 21732 4382 21734
rect 4438 21732 4462 21734
rect 4518 21732 4542 21734
rect 4598 21732 4622 21734
rect 4678 21732 4684 21734
rect 4376 21723 4684 21732
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4356 21146 4384 21490
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 4620 20936 4672 20942
rect 4672 20896 4752 20924
rect 4620 20878 4672 20884
rect 4376 20700 4684 20709
rect 4376 20698 4382 20700
rect 4438 20698 4462 20700
rect 4518 20698 4542 20700
rect 4598 20698 4622 20700
rect 4678 20698 4684 20700
rect 4438 20646 4440 20698
rect 4620 20646 4622 20698
rect 4376 20644 4382 20646
rect 4438 20644 4462 20646
rect 4518 20644 4542 20646
rect 4598 20644 4622 20646
rect 4678 20644 4684 20646
rect 4376 20635 4684 20644
rect 4724 20602 4752 20896
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4620 20256 4672 20262
rect 4724 20210 4752 20538
rect 4672 20204 4752 20210
rect 4620 20198 4752 20204
rect 4632 20182 4752 20198
rect 4172 19808 4292 19836
rect 4172 17762 4200 19808
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4264 17882 4292 19654
rect 4376 19612 4684 19621
rect 4376 19610 4382 19612
rect 4438 19610 4462 19612
rect 4518 19610 4542 19612
rect 4598 19610 4622 19612
rect 4678 19610 4684 19612
rect 4438 19558 4440 19610
rect 4620 19558 4622 19610
rect 4376 19556 4382 19558
rect 4438 19556 4462 19558
rect 4518 19556 4542 19558
rect 4598 19556 4622 19558
rect 4678 19556 4684 19558
rect 4376 19547 4684 19556
rect 4376 18524 4684 18533
rect 4376 18522 4382 18524
rect 4438 18522 4462 18524
rect 4518 18522 4542 18524
rect 4598 18522 4622 18524
rect 4678 18522 4684 18524
rect 4438 18470 4440 18522
rect 4620 18470 4622 18522
rect 4376 18468 4382 18470
rect 4438 18468 4462 18470
rect 4518 18468 4542 18470
rect 4598 18468 4622 18470
rect 4678 18468 4684 18470
rect 4376 18459 4684 18468
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4172 17734 4292 17762
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 16998 4200 17614
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16250 4200 16934
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4264 15162 4292 17734
rect 4724 17678 4752 20182
rect 4816 19514 4844 26318
rect 5368 25906 5396 27338
rect 5644 27130 5672 29200
rect 5736 27606 5764 29294
rect 5906 29200 5962 29294
rect 6012 29294 6238 29322
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 5828 26042 5856 27406
rect 6012 26858 6040 29294
rect 6182 29200 6238 29294
rect 6458 29200 6514 30000
rect 6734 29322 6790 30000
rect 6564 29294 6790 29322
rect 6090 27772 6398 27781
rect 6090 27770 6096 27772
rect 6152 27770 6176 27772
rect 6232 27770 6256 27772
rect 6312 27770 6336 27772
rect 6392 27770 6398 27772
rect 6152 27718 6154 27770
rect 6334 27718 6336 27770
rect 6090 27716 6096 27718
rect 6152 27716 6176 27718
rect 6232 27716 6256 27718
rect 6312 27716 6336 27718
rect 6392 27716 6398 27718
rect 6090 27707 6398 27716
rect 6472 27130 6500 29200
rect 6564 27334 6592 29294
rect 6734 29200 6790 29294
rect 7010 29200 7066 30000
rect 7286 29322 7342 30000
rect 7208 29294 7342 29322
rect 7024 27606 7052 29200
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6552 27328 6604 27334
rect 6552 27270 6604 27276
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6000 26852 6052 26858
rect 6000 26794 6052 26800
rect 6090 26684 6398 26693
rect 6090 26682 6096 26684
rect 6152 26682 6176 26684
rect 6232 26682 6256 26684
rect 6312 26682 6336 26684
rect 6392 26682 6398 26684
rect 6152 26630 6154 26682
rect 6334 26630 6336 26682
rect 6090 26628 6096 26630
rect 6152 26628 6176 26630
rect 6232 26628 6256 26630
rect 6312 26628 6336 26630
rect 6392 26628 6398 26630
rect 6090 26619 6398 26628
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5368 21690 5396 25842
rect 6090 25596 6398 25605
rect 6090 25594 6096 25596
rect 6152 25594 6176 25596
rect 6232 25594 6256 25596
rect 6312 25594 6336 25596
rect 6392 25594 6398 25596
rect 6152 25542 6154 25594
rect 6334 25542 6336 25594
rect 6090 25540 6096 25542
rect 6152 25540 6176 25542
rect 6232 25540 6256 25542
rect 6312 25540 6336 25542
rect 6392 25540 6398 25542
rect 6090 25531 6398 25540
rect 6090 24508 6398 24517
rect 6090 24506 6096 24508
rect 6152 24506 6176 24508
rect 6232 24506 6256 24508
rect 6312 24506 6336 24508
rect 6392 24506 6398 24508
rect 6152 24454 6154 24506
rect 6334 24454 6336 24506
rect 6090 24452 6096 24454
rect 6152 24452 6176 24454
rect 6232 24452 6256 24454
rect 6312 24452 6336 24454
rect 6392 24452 6398 24454
rect 6090 24443 6398 24452
rect 6090 23420 6398 23429
rect 6090 23418 6096 23420
rect 6152 23418 6176 23420
rect 6232 23418 6256 23420
rect 6312 23418 6336 23420
rect 6392 23418 6398 23420
rect 6152 23366 6154 23418
rect 6334 23366 6336 23418
rect 6090 23364 6096 23366
rect 6152 23364 6176 23366
rect 6232 23364 6256 23366
rect 6312 23364 6336 23366
rect 6392 23364 6398 23366
rect 6090 23355 6398 23364
rect 6090 22332 6398 22341
rect 6090 22330 6096 22332
rect 6152 22330 6176 22332
rect 6232 22330 6256 22332
rect 6312 22330 6336 22332
rect 6392 22330 6398 22332
rect 6152 22278 6154 22330
rect 6334 22278 6336 22330
rect 6090 22276 6096 22278
rect 6152 22276 6176 22278
rect 6232 22276 6256 22278
rect 6312 22276 6336 22278
rect 6392 22276 6398 22278
rect 6090 22267 6398 22276
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5460 20942 5488 21966
rect 6090 21244 6398 21253
rect 6090 21242 6096 21244
rect 6152 21242 6176 21244
rect 6232 21242 6256 21244
rect 6312 21242 6336 21244
rect 6392 21242 6398 21244
rect 6152 21190 6154 21242
rect 6334 21190 6336 21242
rect 6090 21188 6096 21190
rect 6152 21188 6176 21190
rect 6232 21188 6256 21190
rect 6312 21188 6336 21190
rect 6392 21188 6398 21190
rect 6090 21179 6398 21188
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 4908 19854 4936 20878
rect 5460 20534 5488 20878
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5460 19854 5488 20470
rect 5552 20058 5580 20742
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 4908 19514 4936 19790
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 5460 19258 5488 19790
rect 5460 19230 5580 19258
rect 5552 18766 5580 19230
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4356 16794 4384 17138
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4724 14482 4752 16050
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4172 14006 4200 14214
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 4724 12442 4752 14418
rect 4816 14414 4844 15574
rect 4908 15570 4936 17478
rect 5184 16046 5212 17614
rect 5368 16250 5396 18634
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15570 5120 15846
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4908 15094 4936 15302
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4816 14278 4844 14350
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 13530 4844 14214
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 5092 12986 5120 15506
rect 5184 13462 5212 15982
rect 5552 15706 5580 18702
rect 5644 17882 5672 20402
rect 5736 19446 5764 21082
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 20466 6224 20878
rect 6564 20602 6592 26182
rect 6656 21146 6684 26386
rect 6748 25922 6776 27338
rect 6840 26382 6868 27406
rect 7208 27130 7236 29294
rect 7286 29200 7342 29294
rect 7562 29200 7618 30000
rect 7838 29322 7894 30000
rect 7668 29294 7894 29322
rect 7576 27554 7604 29200
rect 7484 27526 7604 27554
rect 7484 27334 7512 27526
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7472 27328 7524 27334
rect 7472 27270 7524 27276
rect 7196 27124 7248 27130
rect 7196 27066 7248 27072
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 6932 26382 6960 26930
rect 7024 26586 7052 26930
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 7576 26382 7604 27406
rect 7668 27130 7696 29294
rect 7838 29200 7894 29294
rect 8114 29200 8170 30000
rect 8390 29200 8446 30000
rect 8666 29322 8722 30000
rect 8496 29294 8722 29322
rect 8128 27606 8156 29200
rect 8116 27600 8168 27606
rect 8116 27542 8168 27548
rect 7803 27228 8111 27237
rect 7803 27226 7809 27228
rect 7865 27226 7889 27228
rect 7945 27226 7969 27228
rect 8025 27226 8049 27228
rect 8105 27226 8111 27228
rect 7865 27174 7867 27226
rect 8047 27174 8049 27226
rect 7803 27172 7809 27174
rect 7865 27172 7889 27174
rect 7945 27172 7969 27174
rect 8025 27172 8049 27174
rect 8105 27172 8111 27174
rect 7803 27163 8111 27172
rect 8404 27130 8432 29200
rect 8496 27606 8524 29294
rect 8666 29200 8722 29294
rect 8942 29200 8998 30000
rect 9218 29200 9274 30000
rect 9494 29322 9550 30000
rect 9324 29294 9550 29322
rect 8956 27606 8984 29200
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 7760 26586 7788 26930
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 7564 26376 7616 26382
rect 7564 26318 7616 26324
rect 6840 26246 6868 26318
rect 7104 26308 7156 26314
rect 7104 26250 7156 26256
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6748 25906 6868 25922
rect 6748 25900 6880 25906
rect 6748 25894 6828 25900
rect 6828 25842 6880 25848
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6184 20460 6236 20466
rect 6184 20402 6236 20408
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5828 19514 5856 20334
rect 6090 20156 6398 20165
rect 6090 20154 6096 20156
rect 6152 20154 6176 20156
rect 6232 20154 6256 20156
rect 6312 20154 6336 20156
rect 6392 20154 6398 20156
rect 6152 20102 6154 20154
rect 6334 20102 6336 20154
rect 6090 20100 6096 20102
rect 6152 20100 6176 20102
rect 6232 20100 6256 20102
rect 6312 20100 6336 20102
rect 6392 20100 6398 20102
rect 6090 20091 6398 20100
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5724 19440 5776 19446
rect 5724 19382 5776 19388
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5632 17672 5684 17678
rect 5736 17626 5764 18226
rect 5828 17814 5856 19450
rect 5920 18358 5948 19654
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5920 17746 5948 18294
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5684 17620 5764 17626
rect 5632 17614 5764 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5644 17598 5764 17614
rect 5736 17202 5764 17598
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5644 16658 5672 16934
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5552 15026 5580 15642
rect 5644 15434 5672 16458
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5644 14906 5672 15370
rect 5552 14878 5672 14906
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5276 13938 5304 14350
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11762 4292 12106
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4816 11898 4844 12718
rect 4908 12374 4936 12786
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 4172 9602 4200 10610
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4080 9586 4200 9602
rect 4068 9580 4200 9586
rect 4120 9574 4200 9580
rect 4068 9522 4120 9528
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 4080 7546 4108 9522
rect 4264 8090 4292 10542
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9178 4568 9522
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6390 3832 6598
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 4080 4146 4108 7482
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 5642 4200 6666
rect 4632 6662 4660 7346
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4724 6458 4752 8910
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7546 4844 7822
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4816 6798 4844 7482
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4264 4146 4292 6054
rect 4816 5914 4844 6326
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 756 3052 808 3058
rect 756 2994 808 3000
rect 768 800 796 2994
rect 1872 2446 1900 3334
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 3068 2632 3096 3674
rect 4080 3058 4108 4082
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3602 4384 3878
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2976 2604 3096 2632
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1872 800 1900 2382
rect 2976 800 3004 2604
rect 3252 2446 3280 2790
rect 4172 2650 4200 3402
rect 4264 3194 4292 3538
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 800 4108 2382
rect 4264 2378 4292 3130
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4448 2446 4476 2858
rect 4620 2576 4672 2582
rect 4618 2544 4620 2553
rect 4672 2544 4674 2553
rect 4724 2514 4752 4558
rect 4908 3670 4936 12310
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 4622 5028 11698
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 9450 5212 11018
rect 5276 10742 5304 13874
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 12170 5488 12650
rect 5552 12442 5580 14878
rect 5736 13530 5764 16934
rect 5828 16114 5856 17614
rect 5920 16182 5948 17682
rect 6012 17678 6040 19450
rect 6090 19068 6398 19077
rect 6090 19066 6096 19068
rect 6152 19066 6176 19068
rect 6232 19066 6256 19068
rect 6312 19066 6336 19068
rect 6392 19066 6398 19068
rect 6152 19014 6154 19066
rect 6334 19014 6336 19066
rect 6090 19012 6096 19014
rect 6152 19012 6176 19014
rect 6232 19012 6256 19014
rect 6312 19012 6336 19014
rect 6392 19012 6398 19014
rect 6090 19003 6398 19012
rect 6748 18850 6776 19722
rect 6840 18970 6868 25842
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6932 19378 6960 19790
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6748 18822 6868 18850
rect 6840 18290 6868 18822
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6090 17980 6398 17989
rect 6090 17978 6096 17980
rect 6152 17978 6176 17980
rect 6232 17978 6256 17980
rect 6312 17978 6336 17980
rect 6392 17978 6398 17980
rect 6152 17926 6154 17978
rect 6334 17926 6336 17978
rect 6090 17924 6096 17926
rect 6152 17924 6176 17926
rect 6232 17924 6256 17926
rect 6312 17924 6336 17926
rect 6392 17924 6398 17926
rect 6090 17915 6398 17924
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 16726 6040 17614
rect 6104 16998 6132 17750
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5828 15502 5856 16050
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 13410 5856 15438
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6748 14482 6776 16118
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5644 13382 5856 13410
rect 5644 12646 5672 13382
rect 6012 12986 6040 13874
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5184 8106 5212 9386
rect 5184 8078 5304 8106
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7342 5212 7890
rect 5276 7410 5304 8078
rect 5368 7546 5396 9998
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6118 5120 7142
rect 5184 6798 5212 7278
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5184 5778 5212 6734
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5276 5710 5304 6802
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5276 3942 5304 5646
rect 5368 5642 5396 7482
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 5368 3126 5396 4422
rect 5460 3738 5488 12106
rect 5552 7886 5580 12378
rect 5644 11762 5672 12582
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5920 11694 5948 12038
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11218 5764 11562
rect 5920 11354 5948 11630
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 6472 11150 6500 11698
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6564 10810 6592 13262
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6472 10130 6500 10406
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6656 9450 6684 13194
rect 6748 11626 6776 14418
rect 6840 14346 6868 18226
rect 6932 17678 6960 19314
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17270 6960 17614
rect 7024 17270 7052 18022
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 6932 16658 6960 17206
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6932 16114 6960 16594
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 15094 6960 16050
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7116 14618 7144 26250
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7208 20398 7236 20878
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7208 19854 7236 20334
rect 7576 20058 7604 26318
rect 7803 26140 8111 26149
rect 7803 26138 7809 26140
rect 7865 26138 7889 26140
rect 7945 26138 7969 26140
rect 8025 26138 8049 26140
rect 8105 26138 8111 26140
rect 7865 26086 7867 26138
rect 8047 26086 8049 26138
rect 7803 26084 7809 26086
rect 7865 26084 7889 26086
rect 7945 26084 7969 26086
rect 8025 26084 8049 26086
rect 8105 26084 8111 26086
rect 7803 26075 8111 26084
rect 8496 26042 8524 26930
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 7803 25052 8111 25061
rect 7803 25050 7809 25052
rect 7865 25050 7889 25052
rect 7945 25050 7969 25052
rect 8025 25050 8049 25052
rect 8105 25050 8111 25052
rect 7865 24998 7867 25050
rect 8047 24998 8049 25050
rect 7803 24996 7809 24998
rect 7865 24996 7889 24998
rect 7945 24996 7969 24998
rect 8025 24996 8049 24998
rect 8105 24996 8111 24998
rect 7803 24987 8111 24996
rect 7803 23964 8111 23973
rect 7803 23962 7809 23964
rect 7865 23962 7889 23964
rect 7945 23962 7969 23964
rect 8025 23962 8049 23964
rect 8105 23962 8111 23964
rect 7865 23910 7867 23962
rect 8047 23910 8049 23962
rect 7803 23908 7809 23910
rect 7865 23908 7889 23910
rect 7945 23908 7969 23910
rect 8025 23908 8049 23910
rect 8105 23908 8111 23910
rect 7803 23899 8111 23908
rect 7803 22876 8111 22885
rect 7803 22874 7809 22876
rect 7865 22874 7889 22876
rect 7945 22874 7969 22876
rect 8025 22874 8049 22876
rect 8105 22874 8111 22876
rect 7865 22822 7867 22874
rect 8047 22822 8049 22874
rect 7803 22820 7809 22822
rect 7865 22820 7889 22822
rect 7945 22820 7969 22822
rect 8025 22820 8049 22822
rect 8105 22820 8111 22822
rect 7803 22811 8111 22820
rect 7803 21788 8111 21797
rect 7803 21786 7809 21788
rect 7865 21786 7889 21788
rect 7945 21786 7969 21788
rect 8025 21786 8049 21788
rect 8105 21786 8111 21788
rect 7865 21734 7867 21786
rect 8047 21734 8049 21786
rect 7803 21732 7809 21734
rect 7865 21732 7889 21734
rect 7945 21732 7969 21734
rect 8025 21732 8049 21734
rect 8105 21732 8111 21734
rect 7803 21723 8111 21732
rect 8588 21146 8616 26250
rect 8680 25906 8708 27406
rect 8944 27396 8996 27402
rect 8944 27338 8996 27344
rect 8956 26382 8984 27338
rect 9140 26586 9168 27406
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8668 25900 8720 25906
rect 8668 25842 8720 25848
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 7803 20700 8111 20709
rect 7803 20698 7809 20700
rect 7865 20698 7889 20700
rect 7945 20698 7969 20700
rect 8025 20698 8049 20700
rect 8105 20698 8111 20700
rect 7865 20646 7867 20698
rect 8047 20646 8049 20698
rect 7803 20644 7809 20646
rect 7865 20644 7889 20646
rect 7945 20644 7969 20646
rect 8025 20644 8049 20646
rect 8105 20644 8111 20646
rect 7803 20635 8111 20644
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7803 19612 8111 19621
rect 7803 19610 7809 19612
rect 7865 19610 7889 19612
rect 7945 19610 7969 19612
rect 8025 19610 8049 19612
rect 8105 19610 8111 19612
rect 7865 19558 7867 19610
rect 8047 19558 8049 19610
rect 7803 19556 7809 19558
rect 7865 19556 7889 19558
rect 7945 19556 7969 19558
rect 8025 19556 8049 19558
rect 8105 19556 8111 19558
rect 7803 19547 8111 19556
rect 7803 18524 8111 18533
rect 7803 18522 7809 18524
rect 7865 18522 7889 18524
rect 7945 18522 7969 18524
rect 8025 18522 8049 18524
rect 8105 18522 8111 18524
rect 7865 18470 7867 18522
rect 8047 18470 8049 18522
rect 7803 18468 7809 18470
rect 7865 18468 7889 18470
rect 7945 18468 7969 18470
rect 8025 18468 8049 18470
rect 8105 18468 8111 18470
rect 7803 18459 8111 18468
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 15638 7512 16526
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14618 7420 14962
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7484 14414 7512 15302
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6840 14074 6868 14282
rect 7668 14278 7696 15438
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 8312 14618 8340 20470
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8404 15162 8432 16050
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 11762 7052 13806
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 8220 12782 8248 13262
rect 8496 12986 8524 14350
rect 8588 13530 8616 14962
rect 8680 14890 8708 25842
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8772 19514 8800 25230
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8864 14074 8892 19722
rect 8956 17338 8984 26318
rect 9232 26042 9260 29200
rect 9324 26246 9352 29294
rect 9494 29200 9550 29294
rect 9770 29322 9826 30000
rect 9770 29294 9996 29322
rect 9770 29200 9826 29294
rect 9517 27772 9825 27781
rect 9517 27770 9523 27772
rect 9579 27770 9603 27772
rect 9659 27770 9683 27772
rect 9739 27770 9763 27772
rect 9819 27770 9825 27772
rect 9579 27718 9581 27770
rect 9761 27718 9763 27770
rect 9517 27716 9523 27718
rect 9579 27716 9603 27718
rect 9659 27716 9683 27718
rect 9739 27716 9763 27718
rect 9819 27716 9825 27718
rect 9517 27707 9825 27716
rect 9968 27606 9996 29294
rect 10046 29200 10102 30000
rect 10322 29200 10378 30000
rect 10598 29200 10654 30000
rect 10874 29322 10930 30000
rect 10874 29294 11008 29322
rect 10874 29200 10930 29294
rect 9956 27600 10008 27606
rect 9956 27542 10008 27548
rect 10060 27130 10088 29200
rect 10336 27674 10364 29200
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9416 26586 9444 26930
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9517 26684 9825 26693
rect 9517 26682 9523 26684
rect 9579 26682 9603 26684
rect 9659 26682 9683 26684
rect 9739 26682 9763 26684
rect 9819 26682 9825 26684
rect 9579 26630 9581 26682
rect 9761 26630 9763 26682
rect 9517 26628 9523 26630
rect 9579 26628 9603 26630
rect 9659 26628 9683 26630
rect 9739 26628 9763 26630
rect 9819 26628 9825 26630
rect 9517 26619 9825 26628
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9968 26246 9996 26726
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9956 26240 10008 26246
rect 9956 26182 10008 26188
rect 10152 26042 10180 27270
rect 10244 26382 10272 27338
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10336 26586 10364 26930
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10520 26450 10548 27406
rect 10612 27334 10640 29200
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10980 27112 11008 29294
rect 11150 29200 11206 30000
rect 11426 29322 11482 30000
rect 11426 29294 11652 29322
rect 11426 29200 11482 29294
rect 11060 27124 11112 27130
rect 10980 27084 11060 27112
rect 11060 27066 11112 27072
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10980 26382 11008 26930
rect 11164 26858 11192 29200
rect 11624 27674 11652 29294
rect 11702 29200 11758 30000
rect 11978 29322 12034 30000
rect 11978 29294 12204 29322
rect 11978 29200 12034 29294
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11612 27396 11664 27402
rect 11612 27338 11664 27344
rect 11230 27228 11538 27237
rect 11230 27226 11236 27228
rect 11292 27226 11316 27228
rect 11372 27226 11396 27228
rect 11452 27226 11476 27228
rect 11532 27226 11538 27228
rect 11292 27174 11294 27226
rect 11474 27174 11476 27226
rect 11230 27172 11236 27174
rect 11292 27172 11316 27174
rect 11372 27172 11396 27174
rect 11452 27172 11476 27174
rect 11532 27172 11538 27174
rect 11230 27163 11538 27172
rect 11152 26852 11204 26858
rect 11152 26794 11204 26800
rect 11624 26586 11652 27338
rect 11716 26790 11744 29200
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11796 26988 11848 26994
rect 11796 26930 11848 26936
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11808 26586 11836 26930
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 11992 26382 12020 27474
rect 12176 27130 12204 29294
rect 12254 29200 12310 30000
rect 12530 29322 12586 30000
rect 12530 29294 12756 29322
rect 12530 29200 12586 29294
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 9517 25596 9825 25605
rect 9517 25594 9523 25596
rect 9579 25594 9603 25596
rect 9659 25594 9683 25596
rect 9739 25594 9763 25596
rect 9819 25594 9825 25596
rect 9579 25542 9581 25594
rect 9761 25542 9763 25594
rect 9517 25540 9523 25542
rect 9579 25540 9603 25542
rect 9659 25540 9683 25542
rect 9739 25540 9763 25542
rect 9819 25540 9825 25542
rect 9517 25531 9825 25540
rect 9517 24508 9825 24517
rect 9517 24506 9523 24508
rect 9579 24506 9603 24508
rect 9659 24506 9683 24508
rect 9739 24506 9763 24508
rect 9819 24506 9825 24508
rect 9579 24454 9581 24506
rect 9761 24454 9763 24506
rect 9517 24452 9523 24454
rect 9579 24452 9603 24454
rect 9659 24452 9683 24454
rect 9739 24452 9763 24454
rect 9819 24452 9825 24454
rect 9517 24443 9825 24452
rect 9517 23420 9825 23429
rect 9517 23418 9523 23420
rect 9579 23418 9603 23420
rect 9659 23418 9683 23420
rect 9739 23418 9763 23420
rect 9819 23418 9825 23420
rect 9579 23366 9581 23418
rect 9761 23366 9763 23418
rect 9517 23364 9523 23366
rect 9579 23364 9603 23366
rect 9659 23364 9683 23366
rect 9739 23364 9763 23366
rect 9819 23364 9825 23366
rect 9517 23355 9825 23364
rect 9517 22332 9825 22341
rect 9517 22330 9523 22332
rect 9579 22330 9603 22332
rect 9659 22330 9683 22332
rect 9739 22330 9763 22332
rect 9819 22330 9825 22332
rect 9579 22278 9581 22330
rect 9761 22278 9763 22330
rect 9517 22276 9523 22278
rect 9579 22276 9603 22278
rect 9659 22276 9683 22278
rect 9739 22276 9763 22278
rect 9819 22276 9825 22278
rect 9517 22267 9825 22276
rect 9517 21244 9825 21253
rect 9517 21242 9523 21244
rect 9579 21242 9603 21244
rect 9659 21242 9683 21244
rect 9739 21242 9763 21244
rect 9819 21242 9825 21244
rect 9579 21190 9581 21242
rect 9761 21190 9763 21242
rect 9517 21188 9523 21190
rect 9579 21188 9603 21190
rect 9659 21188 9683 21190
rect 9739 21188 9763 21190
rect 9819 21188 9825 21190
rect 9517 21179 9825 21188
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9048 15162 9076 19314
rect 9140 16454 9168 20810
rect 9517 20156 9825 20165
rect 9517 20154 9523 20156
rect 9579 20154 9603 20156
rect 9659 20154 9683 20156
rect 9739 20154 9763 20156
rect 9819 20154 9825 20156
rect 9579 20102 9581 20154
rect 9761 20102 9763 20154
rect 9517 20100 9523 20102
rect 9579 20100 9603 20102
rect 9659 20100 9683 20102
rect 9739 20100 9763 20102
rect 9819 20100 9825 20102
rect 9517 20091 9825 20100
rect 9517 19068 9825 19077
rect 9517 19066 9523 19068
rect 9579 19066 9603 19068
rect 9659 19066 9683 19068
rect 9739 19066 9763 19068
rect 9819 19066 9825 19068
rect 9579 19014 9581 19066
rect 9761 19014 9763 19066
rect 9517 19012 9523 19014
rect 9579 19012 9603 19014
rect 9659 19012 9683 19014
rect 9739 19012 9763 19014
rect 9819 19012 9825 19014
rect 9517 19003 9825 19012
rect 9517 17980 9825 17989
rect 9517 17978 9523 17980
rect 9579 17978 9603 17980
rect 9659 17978 9683 17980
rect 9739 17978 9763 17980
rect 9819 17978 9825 17980
rect 9579 17926 9581 17978
rect 9761 17926 9763 17978
rect 9517 17924 9523 17926
rect 9579 17924 9603 17926
rect 9659 17924 9683 17926
rect 9739 17924 9763 17926
rect 9819 17924 9825 17926
rect 9517 17915 9825 17924
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9232 15178 9260 17546
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9140 15150 9260 15178
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 7668 12434 7696 12718
rect 7576 12406 7696 12434
rect 7576 12238 7604 12406
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7576 11898 7604 12174
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6932 10538 6960 11222
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 9602 6960 10474
rect 7024 10062 7052 11698
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6840 9574 6960 9602
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6840 9178 6868 9574
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5828 8634 5856 8910
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7562 5580 7822
rect 5552 7534 5672 7562
rect 5644 7478 5672 7534
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5552 6458 5580 7346
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5552 5914 5580 6122
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5778 5672 6258
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 4826 5580 5510
rect 5736 5370 5764 8298
rect 5920 6730 5948 8774
rect 6012 7342 6040 8910
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6748 8090 6776 8434
rect 6840 8362 6868 9114
rect 6932 8566 6960 9386
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 6656 6662 6684 7346
rect 6748 6798 6776 8026
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 4622 5672 5238
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5736 4826 5764 5102
rect 5828 5030 5856 6258
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5552 4010 5580 4558
rect 6012 4146 6040 6122
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6656 5574 6684 6598
rect 6748 6322 6776 6734
rect 6932 6662 6960 8502
rect 7024 8498 7052 9998
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6458 6960 6598
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5370 6684 5510
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6656 5250 6684 5306
rect 6564 5222 6684 5250
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6472 4622 6500 4966
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 6012 3194 6040 4082
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6472 3738 6500 4558
rect 6564 4214 6592 5222
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4282 6684 4422
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4146 6684 4218
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6472 3194 6500 3674
rect 6748 3602 6776 6258
rect 6840 5914 6868 6258
rect 7024 6118 7052 8298
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4146 6868 5102
rect 6932 4826 6960 5238
rect 7024 5098 7052 6054
rect 7116 5137 7144 10678
rect 7208 10606 7236 11154
rect 7930 11112 7986 11121
rect 7930 11047 7932 11056
rect 7984 11047 7986 11056
rect 7932 11018 7984 11024
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 9738 7236 10542
rect 7208 9710 7328 9738
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7102 5128 7158 5137
rect 7012 5092 7064 5098
rect 7102 5063 7158 5072
rect 7012 5034 7064 5040
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 4618 2479 4674 2488
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5828 2446 5856 2790
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6564 2650 6592 3402
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7024 2514 7052 2926
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7116 2446 7144 4966
rect 7208 2650 7236 9522
rect 7300 9518 7328 9710
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 8974 7328 9454
rect 7484 9178 7512 9522
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8090 7328 8774
rect 7392 8566 7420 9046
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5234 7328 5646
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7286 5128 7342 5137
rect 7484 5114 7512 8910
rect 7286 5063 7342 5072
rect 7392 5086 7512 5114
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 2582 7328 5063
rect 7392 4622 7420 5086
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4026 7420 4558
rect 7484 4146 7512 4966
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7392 3998 7512 4026
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3534 7420 3878
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 2990 7512 3998
rect 7576 3194 7604 10610
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9722 7696 9930
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7668 7274 7696 7754
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 8220 4826 8248 12174
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8588 10538 8616 11698
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8362 8340 8910
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 7886 8340 8298
rect 8404 7954 8432 9862
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7478 8340 7686
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 6798 8340 7414
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 5846 8340 6734
rect 8404 6390 8432 7890
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 6866 8616 7686
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6474 8616 6802
rect 8496 6458 8616 6474
rect 8680 6458 8708 13262
rect 8772 11898 8800 13874
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8498 8800 8774
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 7478 8800 8434
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8864 6662 8892 12786
rect 9048 12442 9076 13874
rect 9140 13530 9168 15150
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 12986 9260 14962
rect 9324 14618 9352 16526
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14414 9444 15438
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9232 10810 9260 11698
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9140 10266 9168 10610
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8956 8090 8984 8298
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9048 8022 9076 8978
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 8634 9168 8842
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8484 6452 8616 6458
rect 8536 6446 8616 6452
rect 8484 6394 8536 6400
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4622 8340 5646
rect 8404 5574 8432 6326
rect 8588 5846 8616 6446
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 8312 4214 8340 4558
rect 8404 4554 8432 4626
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8312 3738 8340 4150
rect 8404 4078 8432 4490
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 9048 3942 9076 7958
rect 9324 7546 9352 12786
rect 9416 12714 9444 14350
rect 10336 14006 10364 26318
rect 11230 26140 11538 26149
rect 11230 26138 11236 26140
rect 11292 26138 11316 26140
rect 11372 26138 11396 26140
rect 11452 26138 11476 26140
rect 11532 26138 11538 26140
rect 11292 26086 11294 26138
rect 11474 26086 11476 26138
rect 11230 26084 11236 26086
rect 11292 26084 11316 26086
rect 11372 26084 11396 26086
rect 11452 26084 11476 26086
rect 11532 26084 11538 26086
rect 11230 26075 11538 26084
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10888 25265 10916 25842
rect 10874 25256 10930 25265
rect 10874 25191 10930 25200
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12986 9812 13262
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 10062 9444 12650
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 8430 9444 9998
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9232 6798 9260 7210
rect 9416 6866 9444 8026
rect 9876 7886 9904 8502
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6254 9260 6734
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 4690 9260 6190
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9876 5710 9904 7822
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7392 2446 7420 2858
rect 8404 2650 8432 2994
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8496 2446 8524 2790
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 9876 2650 9904 4150
rect 10060 4010 10088 12786
rect 10888 11626 10916 25191
rect 11230 25052 11538 25061
rect 11230 25050 11236 25052
rect 11292 25050 11316 25052
rect 11372 25050 11396 25052
rect 11452 25050 11476 25052
rect 11532 25050 11538 25052
rect 11292 24998 11294 25050
rect 11474 24998 11476 25050
rect 11230 24996 11236 24998
rect 11292 24996 11316 24998
rect 11372 24996 11396 24998
rect 11452 24996 11476 24998
rect 11532 24996 11538 24998
rect 11230 24987 11538 24996
rect 11230 23964 11538 23973
rect 11230 23962 11236 23964
rect 11292 23962 11316 23964
rect 11372 23962 11396 23964
rect 11452 23962 11476 23964
rect 11532 23962 11538 23964
rect 11292 23910 11294 23962
rect 11474 23910 11476 23962
rect 11230 23908 11236 23910
rect 11292 23908 11316 23910
rect 11372 23908 11396 23910
rect 11452 23908 11476 23910
rect 11532 23908 11538 23910
rect 11230 23899 11538 23908
rect 11230 22876 11538 22885
rect 11230 22874 11236 22876
rect 11292 22874 11316 22876
rect 11372 22874 11396 22876
rect 11452 22874 11476 22876
rect 11532 22874 11538 22876
rect 11292 22822 11294 22874
rect 11474 22822 11476 22874
rect 11230 22820 11236 22822
rect 11292 22820 11316 22822
rect 11372 22820 11396 22822
rect 11452 22820 11476 22822
rect 11532 22820 11538 22822
rect 11230 22811 11538 22820
rect 11230 21788 11538 21797
rect 11230 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11396 21788
rect 11452 21786 11476 21788
rect 11532 21786 11538 21788
rect 11292 21734 11294 21786
rect 11474 21734 11476 21786
rect 11230 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11396 21734
rect 11452 21732 11476 21734
rect 11532 21732 11538 21734
rect 11230 21723 11538 21732
rect 11230 20700 11538 20709
rect 11230 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11396 20700
rect 11452 20698 11476 20700
rect 11532 20698 11538 20700
rect 11292 20646 11294 20698
rect 11474 20646 11476 20698
rect 11230 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11396 20646
rect 11452 20644 11476 20646
rect 11532 20644 11538 20646
rect 11230 20635 11538 20644
rect 11230 19612 11538 19621
rect 11230 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11396 19612
rect 11452 19610 11476 19612
rect 11532 19610 11538 19612
rect 11292 19558 11294 19610
rect 11474 19558 11476 19610
rect 11230 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11396 19558
rect 11452 19556 11476 19558
rect 11532 19556 11538 19558
rect 11230 19547 11538 19556
rect 11230 18524 11538 18533
rect 11230 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11396 18524
rect 11452 18522 11476 18524
rect 11532 18522 11538 18524
rect 11292 18470 11294 18522
rect 11474 18470 11476 18522
rect 11230 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11396 18470
rect 11452 18468 11476 18470
rect 11532 18468 11538 18470
rect 11230 18459 11538 18468
rect 11624 17882 11652 26318
rect 12268 26042 12296 29200
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12544 26586 12572 26930
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 11888 25832 11940 25838
rect 11888 25774 11940 25780
rect 11900 25294 11928 25774
rect 12176 25294 12204 25842
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 12176 16250 12204 25230
rect 12452 20058 12480 26318
rect 12530 25256 12586 25265
rect 12530 25191 12586 25200
rect 12544 24818 12572 25191
rect 12636 24834 12664 26318
rect 12728 25498 12756 29294
rect 12806 29200 12862 30000
rect 13082 29322 13138 30000
rect 13358 29322 13414 30000
rect 13082 29294 13308 29322
rect 13082 29200 13138 29294
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12820 25378 12848 29200
rect 12944 27772 13252 27781
rect 12944 27770 12950 27772
rect 13006 27770 13030 27772
rect 13086 27770 13110 27772
rect 13166 27770 13190 27772
rect 13246 27770 13252 27772
rect 13006 27718 13008 27770
rect 13188 27718 13190 27770
rect 12944 27716 12950 27718
rect 13006 27716 13030 27718
rect 13086 27716 13110 27718
rect 13166 27716 13190 27718
rect 13246 27716 13252 27718
rect 12944 27707 13252 27716
rect 12944 26684 13252 26693
rect 12944 26682 12950 26684
rect 13006 26682 13030 26684
rect 13086 26682 13110 26684
rect 13166 26682 13190 26684
rect 13246 26682 13252 26684
rect 13006 26630 13008 26682
rect 13188 26630 13190 26682
rect 12944 26628 12950 26630
rect 13006 26628 13030 26630
rect 13086 26628 13110 26630
rect 13166 26628 13190 26630
rect 13246 26628 13252 26630
rect 12944 26619 13252 26628
rect 12944 25596 13252 25605
rect 12944 25594 12950 25596
rect 13006 25594 13030 25596
rect 13086 25594 13110 25596
rect 13166 25594 13190 25596
rect 13246 25594 13252 25596
rect 13006 25542 13008 25594
rect 13188 25542 13190 25594
rect 12944 25540 12950 25542
rect 13006 25540 13030 25542
rect 13086 25540 13110 25542
rect 13166 25540 13190 25542
rect 13246 25540 13252 25542
rect 12944 25531 13252 25540
rect 12900 25424 12952 25430
rect 12820 25372 12900 25378
rect 12820 25366 12952 25372
rect 12820 25350 12940 25366
rect 12636 24818 12848 24834
rect 12532 24812 12584 24818
rect 12636 24812 12860 24818
rect 12636 24806 12808 24812
rect 12532 24754 12584 24760
rect 12808 24754 12860 24760
rect 12820 20602 12848 24754
rect 13280 24682 13308 29294
rect 13358 29294 13492 29322
rect 13358 29200 13414 29294
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13372 26450 13400 26930
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13372 25294 13400 26250
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 12944 24508 13252 24517
rect 12944 24506 12950 24508
rect 13006 24506 13030 24508
rect 13086 24506 13110 24508
rect 13166 24506 13190 24508
rect 13246 24506 13252 24508
rect 13006 24454 13008 24506
rect 13188 24454 13190 24506
rect 12944 24452 12950 24454
rect 13006 24452 13030 24454
rect 13086 24452 13110 24454
rect 13166 24452 13190 24454
rect 13246 24452 13252 24454
rect 12944 24443 13252 24452
rect 13464 24410 13492 29294
rect 13634 29200 13690 30000
rect 13910 29200 13966 30000
rect 14186 29200 14242 30000
rect 13648 25158 13676 29200
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13740 24206 13768 25638
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13924 23866 13952 29200
rect 14200 25770 14228 29200
rect 14657 27228 14965 27237
rect 14657 27226 14663 27228
rect 14719 27226 14743 27228
rect 14799 27226 14823 27228
rect 14879 27226 14903 27228
rect 14959 27226 14965 27228
rect 14719 27174 14721 27226
rect 14901 27174 14903 27226
rect 14657 27172 14663 27174
rect 14719 27172 14743 27174
rect 14799 27172 14823 27174
rect 14879 27172 14903 27174
rect 14959 27172 14965 27174
rect 14657 27163 14965 27172
rect 14657 26140 14965 26149
rect 14657 26138 14663 26140
rect 14719 26138 14743 26140
rect 14799 26138 14823 26140
rect 14879 26138 14903 26140
rect 14959 26138 14965 26140
rect 14719 26086 14721 26138
rect 14901 26086 14903 26138
rect 14657 26084 14663 26086
rect 14719 26084 14743 26086
rect 14799 26084 14823 26086
rect 14879 26084 14903 26086
rect 14959 26084 14965 26086
rect 14657 26075 14965 26084
rect 14188 25764 14240 25770
rect 14188 25706 14240 25712
rect 14657 25052 14965 25061
rect 14657 25050 14663 25052
rect 14719 25050 14743 25052
rect 14799 25050 14823 25052
rect 14879 25050 14903 25052
rect 14959 25050 14965 25052
rect 14719 24998 14721 25050
rect 14901 24998 14903 25050
rect 14657 24996 14663 24998
rect 14719 24996 14743 24998
rect 14799 24996 14823 24998
rect 14879 24996 14903 24998
rect 14959 24996 14965 24998
rect 14657 24987 14965 24996
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14016 23730 14044 24550
rect 14657 23964 14965 23973
rect 14657 23962 14663 23964
rect 14719 23962 14743 23964
rect 14799 23962 14823 23964
rect 14879 23962 14903 23964
rect 14959 23962 14965 23964
rect 14719 23910 14721 23962
rect 14901 23910 14903 23962
rect 14657 23908 14663 23910
rect 14719 23908 14743 23910
rect 14799 23908 14823 23910
rect 14879 23908 14903 23910
rect 14959 23908 14965 23910
rect 14657 23899 14965 23908
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 12944 23420 13252 23429
rect 12944 23418 12950 23420
rect 13006 23418 13030 23420
rect 13086 23418 13110 23420
rect 13166 23418 13190 23420
rect 13246 23418 13252 23420
rect 13006 23366 13008 23418
rect 13188 23366 13190 23418
rect 12944 23364 12950 23366
rect 13006 23364 13030 23366
rect 13086 23364 13110 23366
rect 13166 23364 13190 23366
rect 13246 23364 13252 23366
rect 12944 23355 13252 23364
rect 14657 22876 14965 22885
rect 14657 22874 14663 22876
rect 14719 22874 14743 22876
rect 14799 22874 14823 22876
rect 14879 22874 14903 22876
rect 14959 22874 14965 22876
rect 14719 22822 14721 22874
rect 14901 22822 14903 22874
rect 14657 22820 14663 22822
rect 14719 22820 14743 22822
rect 14799 22820 14823 22822
rect 14879 22820 14903 22822
rect 14959 22820 14965 22822
rect 14657 22811 14965 22820
rect 12944 22332 13252 22341
rect 12944 22330 12950 22332
rect 13006 22330 13030 22332
rect 13086 22330 13110 22332
rect 13166 22330 13190 22332
rect 13246 22330 13252 22332
rect 13006 22278 13008 22330
rect 13188 22278 13190 22330
rect 12944 22276 12950 22278
rect 13006 22276 13030 22278
rect 13086 22276 13110 22278
rect 13166 22276 13190 22278
rect 13246 22276 13252 22278
rect 12944 22267 13252 22276
rect 14657 21788 14965 21797
rect 14657 21786 14663 21788
rect 14719 21786 14743 21788
rect 14799 21786 14823 21788
rect 14879 21786 14903 21788
rect 14959 21786 14965 21788
rect 14719 21734 14721 21786
rect 14901 21734 14903 21786
rect 14657 21732 14663 21734
rect 14719 21732 14743 21734
rect 14799 21732 14823 21734
rect 14879 21732 14903 21734
rect 14959 21732 14965 21734
rect 14657 21723 14965 21732
rect 12944 21244 13252 21253
rect 12944 21242 12950 21244
rect 13006 21242 13030 21244
rect 13086 21242 13110 21244
rect 13166 21242 13190 21244
rect 13246 21242 13252 21244
rect 13006 21190 13008 21242
rect 13188 21190 13190 21242
rect 12944 21188 12950 21190
rect 13006 21188 13030 21190
rect 13086 21188 13110 21190
rect 13166 21188 13190 21190
rect 13246 21188 13252 21190
rect 12944 21179 13252 21188
rect 14657 20700 14965 20709
rect 14657 20698 14663 20700
rect 14719 20698 14743 20700
rect 14799 20698 14823 20700
rect 14879 20698 14903 20700
rect 14959 20698 14965 20700
rect 14719 20646 14721 20698
rect 14901 20646 14903 20698
rect 14657 20644 14663 20646
rect 14719 20644 14743 20646
rect 14799 20644 14823 20646
rect 14879 20644 14903 20646
rect 14959 20644 14965 20646
rect 14657 20635 14965 20644
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12944 20156 13252 20165
rect 12944 20154 12950 20156
rect 13006 20154 13030 20156
rect 13086 20154 13110 20156
rect 13166 20154 13190 20156
rect 13246 20154 13252 20156
rect 13006 20102 13008 20154
rect 13188 20102 13190 20154
rect 12944 20100 12950 20102
rect 13006 20100 13030 20102
rect 13086 20100 13110 20102
rect 13166 20100 13190 20102
rect 13246 20100 13252 20102
rect 12944 20091 13252 20100
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 14657 19612 14965 19621
rect 14657 19610 14663 19612
rect 14719 19610 14743 19612
rect 14799 19610 14823 19612
rect 14879 19610 14903 19612
rect 14959 19610 14965 19612
rect 14719 19558 14721 19610
rect 14901 19558 14903 19610
rect 14657 19556 14663 19558
rect 14719 19556 14743 19558
rect 14799 19556 14823 19558
rect 14879 19556 14903 19558
rect 14959 19556 14965 19558
rect 14657 19547 14965 19556
rect 12944 19068 13252 19077
rect 12944 19066 12950 19068
rect 13006 19066 13030 19068
rect 13086 19066 13110 19068
rect 13166 19066 13190 19068
rect 13246 19066 13252 19068
rect 13006 19014 13008 19066
rect 13188 19014 13190 19066
rect 12944 19012 12950 19014
rect 13006 19012 13030 19014
rect 13086 19012 13110 19014
rect 13166 19012 13190 19014
rect 13246 19012 13252 19014
rect 12944 19003 13252 19012
rect 14657 18524 14965 18533
rect 14657 18522 14663 18524
rect 14719 18522 14743 18524
rect 14799 18522 14823 18524
rect 14879 18522 14903 18524
rect 14959 18522 14965 18524
rect 14719 18470 14721 18522
rect 14901 18470 14903 18522
rect 14657 18468 14663 18470
rect 14719 18468 14743 18470
rect 14799 18468 14823 18470
rect 14879 18468 14903 18470
rect 14959 18468 14965 18470
rect 14657 18459 14965 18468
rect 12944 17980 13252 17989
rect 12944 17978 12950 17980
rect 13006 17978 13030 17980
rect 13086 17978 13110 17980
rect 13166 17978 13190 17980
rect 13246 17978 13252 17980
rect 13006 17926 13008 17978
rect 13188 17926 13190 17978
rect 12944 17924 12950 17926
rect 13006 17924 13030 17926
rect 13086 17924 13110 17926
rect 13166 17924 13190 17926
rect 13246 17924 13252 17926
rect 12944 17915 13252 17924
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10704 2446 10732 2790
rect 10796 2650 10824 4490
rect 10980 2650 11008 6258
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11808 2446 11836 2790
rect 12452 2650 12480 6598
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 13464 3194 13492 9930
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 14016 3058 14044 3334
rect 14108 3194 14136 7346
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 5080 2440 5132 2446
rect 5816 2440 5868 2446
rect 5132 2400 5212 2428
rect 5080 2382 5132 2388
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 5184 800 5212 2400
rect 5816 2382 5868 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 6288 800 6316 2382
rect 7392 800 7420 2382
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 8496 800 8524 2382
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9600 800 9628 2246
rect 10704 800 10732 2382
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 11808 800 11836 2382
rect 12912 800 12940 2382
rect 14016 800 14044 2994
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 15120 800 15148 2926
rect 754 0 810 800
rect 1858 0 1914 800
rect 2962 0 3018 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10690 0 10746 800
rect 11794 0 11850 800
rect 12898 0 12954 800
rect 14002 0 14058 800
rect 15106 0 15162 800
<< via2 >>
rect 2669 27770 2725 27772
rect 2749 27770 2805 27772
rect 2829 27770 2885 27772
rect 2909 27770 2965 27772
rect 2669 27718 2715 27770
rect 2715 27718 2725 27770
rect 2749 27718 2779 27770
rect 2779 27718 2791 27770
rect 2791 27718 2805 27770
rect 2829 27718 2843 27770
rect 2843 27718 2855 27770
rect 2855 27718 2885 27770
rect 2909 27718 2919 27770
rect 2919 27718 2965 27770
rect 2669 27716 2725 27718
rect 2749 27716 2805 27718
rect 2829 27716 2885 27718
rect 2909 27716 2965 27718
rect 2669 26682 2725 26684
rect 2749 26682 2805 26684
rect 2829 26682 2885 26684
rect 2909 26682 2965 26684
rect 2669 26630 2715 26682
rect 2715 26630 2725 26682
rect 2749 26630 2779 26682
rect 2779 26630 2791 26682
rect 2791 26630 2805 26682
rect 2829 26630 2843 26682
rect 2843 26630 2855 26682
rect 2855 26630 2885 26682
rect 2909 26630 2919 26682
rect 2919 26630 2965 26682
rect 2669 26628 2725 26630
rect 2749 26628 2805 26630
rect 2829 26628 2885 26630
rect 2909 26628 2965 26630
rect 2669 25594 2725 25596
rect 2749 25594 2805 25596
rect 2829 25594 2885 25596
rect 2909 25594 2965 25596
rect 2669 25542 2715 25594
rect 2715 25542 2725 25594
rect 2749 25542 2779 25594
rect 2779 25542 2791 25594
rect 2791 25542 2805 25594
rect 2829 25542 2843 25594
rect 2843 25542 2855 25594
rect 2855 25542 2885 25594
rect 2909 25542 2919 25594
rect 2919 25542 2965 25594
rect 2669 25540 2725 25542
rect 2749 25540 2805 25542
rect 2829 25540 2885 25542
rect 2909 25540 2965 25542
rect 2669 24506 2725 24508
rect 2749 24506 2805 24508
rect 2829 24506 2885 24508
rect 2909 24506 2965 24508
rect 2669 24454 2715 24506
rect 2715 24454 2725 24506
rect 2749 24454 2779 24506
rect 2779 24454 2791 24506
rect 2791 24454 2805 24506
rect 2829 24454 2843 24506
rect 2843 24454 2855 24506
rect 2855 24454 2885 24506
rect 2909 24454 2919 24506
rect 2919 24454 2965 24506
rect 2669 24452 2725 24454
rect 2749 24452 2805 24454
rect 2829 24452 2885 24454
rect 2909 24452 2965 24454
rect 2669 23418 2725 23420
rect 2749 23418 2805 23420
rect 2829 23418 2885 23420
rect 2909 23418 2965 23420
rect 2669 23366 2715 23418
rect 2715 23366 2725 23418
rect 2749 23366 2779 23418
rect 2779 23366 2791 23418
rect 2791 23366 2805 23418
rect 2829 23366 2843 23418
rect 2843 23366 2855 23418
rect 2855 23366 2885 23418
rect 2909 23366 2919 23418
rect 2919 23366 2965 23418
rect 2669 23364 2725 23366
rect 2749 23364 2805 23366
rect 2829 23364 2885 23366
rect 2909 23364 2965 23366
rect 2669 22330 2725 22332
rect 2749 22330 2805 22332
rect 2829 22330 2885 22332
rect 2909 22330 2965 22332
rect 2669 22278 2715 22330
rect 2715 22278 2725 22330
rect 2749 22278 2779 22330
rect 2779 22278 2791 22330
rect 2791 22278 2805 22330
rect 2829 22278 2843 22330
rect 2843 22278 2855 22330
rect 2855 22278 2885 22330
rect 2909 22278 2919 22330
rect 2919 22278 2965 22330
rect 2669 22276 2725 22278
rect 2749 22276 2805 22278
rect 2829 22276 2885 22278
rect 2909 22276 2965 22278
rect 2669 21242 2725 21244
rect 2749 21242 2805 21244
rect 2829 21242 2885 21244
rect 2909 21242 2965 21244
rect 2669 21190 2715 21242
rect 2715 21190 2725 21242
rect 2749 21190 2779 21242
rect 2779 21190 2791 21242
rect 2791 21190 2805 21242
rect 2829 21190 2843 21242
rect 2843 21190 2855 21242
rect 2855 21190 2885 21242
rect 2909 21190 2919 21242
rect 2919 21190 2965 21242
rect 2669 21188 2725 21190
rect 2749 21188 2805 21190
rect 2829 21188 2885 21190
rect 2909 21188 2965 21190
rect 2669 20154 2725 20156
rect 2749 20154 2805 20156
rect 2829 20154 2885 20156
rect 2909 20154 2965 20156
rect 2669 20102 2715 20154
rect 2715 20102 2725 20154
rect 2749 20102 2779 20154
rect 2779 20102 2791 20154
rect 2791 20102 2805 20154
rect 2829 20102 2843 20154
rect 2843 20102 2855 20154
rect 2855 20102 2885 20154
rect 2909 20102 2919 20154
rect 2919 20102 2965 20154
rect 2669 20100 2725 20102
rect 2749 20100 2805 20102
rect 2829 20100 2885 20102
rect 2909 20100 2965 20102
rect 2669 19066 2725 19068
rect 2749 19066 2805 19068
rect 2829 19066 2885 19068
rect 2909 19066 2965 19068
rect 2669 19014 2715 19066
rect 2715 19014 2725 19066
rect 2749 19014 2779 19066
rect 2779 19014 2791 19066
rect 2791 19014 2805 19066
rect 2829 19014 2843 19066
rect 2843 19014 2855 19066
rect 2855 19014 2885 19066
rect 2909 19014 2919 19066
rect 2919 19014 2965 19066
rect 2669 19012 2725 19014
rect 2749 19012 2805 19014
rect 2829 19012 2885 19014
rect 2909 19012 2965 19014
rect 2669 17978 2725 17980
rect 2749 17978 2805 17980
rect 2829 17978 2885 17980
rect 2909 17978 2965 17980
rect 2669 17926 2715 17978
rect 2715 17926 2725 17978
rect 2749 17926 2779 17978
rect 2779 17926 2791 17978
rect 2791 17926 2805 17978
rect 2829 17926 2843 17978
rect 2843 17926 2855 17978
rect 2855 17926 2885 17978
rect 2909 17926 2919 17978
rect 2919 17926 2965 17978
rect 2669 17924 2725 17926
rect 2749 17924 2805 17926
rect 2829 17924 2885 17926
rect 2909 17924 2965 17926
rect 4382 27226 4438 27228
rect 4462 27226 4518 27228
rect 4542 27226 4598 27228
rect 4622 27226 4678 27228
rect 4382 27174 4428 27226
rect 4428 27174 4438 27226
rect 4462 27174 4492 27226
rect 4492 27174 4504 27226
rect 4504 27174 4518 27226
rect 4542 27174 4556 27226
rect 4556 27174 4568 27226
rect 4568 27174 4598 27226
rect 4622 27174 4632 27226
rect 4632 27174 4678 27226
rect 4382 27172 4438 27174
rect 4462 27172 4518 27174
rect 4542 27172 4598 27174
rect 4622 27172 4678 27174
rect 4382 26138 4438 26140
rect 4462 26138 4518 26140
rect 4542 26138 4598 26140
rect 4622 26138 4678 26140
rect 4382 26086 4428 26138
rect 4428 26086 4438 26138
rect 4462 26086 4492 26138
rect 4492 26086 4504 26138
rect 4504 26086 4518 26138
rect 4542 26086 4556 26138
rect 4556 26086 4568 26138
rect 4568 26086 4598 26138
rect 4622 26086 4632 26138
rect 4632 26086 4678 26138
rect 4382 26084 4438 26086
rect 4462 26084 4518 26086
rect 4542 26084 4598 26086
rect 4622 26084 4678 26086
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 4382 25050 4438 25052
rect 4462 25050 4518 25052
rect 4542 25050 4598 25052
rect 4622 25050 4678 25052
rect 4382 24998 4428 25050
rect 4428 24998 4438 25050
rect 4462 24998 4492 25050
rect 4492 24998 4504 25050
rect 4504 24998 4518 25050
rect 4542 24998 4556 25050
rect 4556 24998 4568 25050
rect 4568 24998 4598 25050
rect 4622 24998 4632 25050
rect 4632 24998 4678 25050
rect 4382 24996 4438 24998
rect 4462 24996 4518 24998
rect 4542 24996 4598 24998
rect 4622 24996 4678 24998
rect 4382 23962 4438 23964
rect 4462 23962 4518 23964
rect 4542 23962 4598 23964
rect 4622 23962 4678 23964
rect 4382 23910 4428 23962
rect 4428 23910 4438 23962
rect 4462 23910 4492 23962
rect 4492 23910 4504 23962
rect 4504 23910 4518 23962
rect 4542 23910 4556 23962
rect 4556 23910 4568 23962
rect 4568 23910 4598 23962
rect 4622 23910 4632 23962
rect 4632 23910 4678 23962
rect 4382 23908 4438 23910
rect 4462 23908 4518 23910
rect 4542 23908 4598 23910
rect 4622 23908 4678 23910
rect 4382 22874 4438 22876
rect 4462 22874 4518 22876
rect 4542 22874 4598 22876
rect 4622 22874 4678 22876
rect 4382 22822 4428 22874
rect 4428 22822 4438 22874
rect 4462 22822 4492 22874
rect 4492 22822 4504 22874
rect 4504 22822 4518 22874
rect 4542 22822 4556 22874
rect 4556 22822 4568 22874
rect 4568 22822 4598 22874
rect 4622 22822 4632 22874
rect 4632 22822 4678 22874
rect 4382 22820 4438 22822
rect 4462 22820 4518 22822
rect 4542 22820 4598 22822
rect 4622 22820 4678 22822
rect 4382 21786 4438 21788
rect 4462 21786 4518 21788
rect 4542 21786 4598 21788
rect 4622 21786 4678 21788
rect 4382 21734 4428 21786
rect 4428 21734 4438 21786
rect 4462 21734 4492 21786
rect 4492 21734 4504 21786
rect 4504 21734 4518 21786
rect 4542 21734 4556 21786
rect 4556 21734 4568 21786
rect 4568 21734 4598 21786
rect 4622 21734 4632 21786
rect 4632 21734 4678 21786
rect 4382 21732 4438 21734
rect 4462 21732 4518 21734
rect 4542 21732 4598 21734
rect 4622 21732 4678 21734
rect 4382 20698 4438 20700
rect 4462 20698 4518 20700
rect 4542 20698 4598 20700
rect 4622 20698 4678 20700
rect 4382 20646 4428 20698
rect 4428 20646 4438 20698
rect 4462 20646 4492 20698
rect 4492 20646 4504 20698
rect 4504 20646 4518 20698
rect 4542 20646 4556 20698
rect 4556 20646 4568 20698
rect 4568 20646 4598 20698
rect 4622 20646 4632 20698
rect 4632 20646 4678 20698
rect 4382 20644 4438 20646
rect 4462 20644 4518 20646
rect 4542 20644 4598 20646
rect 4622 20644 4678 20646
rect 4382 19610 4438 19612
rect 4462 19610 4518 19612
rect 4542 19610 4598 19612
rect 4622 19610 4678 19612
rect 4382 19558 4428 19610
rect 4428 19558 4438 19610
rect 4462 19558 4492 19610
rect 4492 19558 4504 19610
rect 4504 19558 4518 19610
rect 4542 19558 4556 19610
rect 4556 19558 4568 19610
rect 4568 19558 4598 19610
rect 4622 19558 4632 19610
rect 4632 19558 4678 19610
rect 4382 19556 4438 19558
rect 4462 19556 4518 19558
rect 4542 19556 4598 19558
rect 4622 19556 4678 19558
rect 4382 18522 4438 18524
rect 4462 18522 4518 18524
rect 4542 18522 4598 18524
rect 4622 18522 4678 18524
rect 4382 18470 4428 18522
rect 4428 18470 4438 18522
rect 4462 18470 4492 18522
rect 4492 18470 4504 18522
rect 4504 18470 4518 18522
rect 4542 18470 4556 18522
rect 4556 18470 4568 18522
rect 4568 18470 4598 18522
rect 4622 18470 4632 18522
rect 4632 18470 4678 18522
rect 4382 18468 4438 18470
rect 4462 18468 4518 18470
rect 4542 18468 4598 18470
rect 4622 18468 4678 18470
rect 6096 27770 6152 27772
rect 6176 27770 6232 27772
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6096 27718 6142 27770
rect 6142 27718 6152 27770
rect 6176 27718 6206 27770
rect 6206 27718 6218 27770
rect 6218 27718 6232 27770
rect 6256 27718 6270 27770
rect 6270 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6096 27716 6152 27718
rect 6176 27716 6232 27718
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 6096 26682 6152 26684
rect 6176 26682 6232 26684
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6096 26630 6142 26682
rect 6142 26630 6152 26682
rect 6176 26630 6206 26682
rect 6206 26630 6218 26682
rect 6218 26630 6232 26682
rect 6256 26630 6270 26682
rect 6270 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6096 26628 6152 26630
rect 6176 26628 6232 26630
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 6096 25594 6152 25596
rect 6176 25594 6232 25596
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6096 25542 6142 25594
rect 6142 25542 6152 25594
rect 6176 25542 6206 25594
rect 6206 25542 6218 25594
rect 6218 25542 6232 25594
rect 6256 25542 6270 25594
rect 6270 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6096 25540 6152 25542
rect 6176 25540 6232 25542
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 6096 24506 6152 24508
rect 6176 24506 6232 24508
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6096 24454 6142 24506
rect 6142 24454 6152 24506
rect 6176 24454 6206 24506
rect 6206 24454 6218 24506
rect 6218 24454 6232 24506
rect 6256 24454 6270 24506
rect 6270 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6096 24452 6152 24454
rect 6176 24452 6232 24454
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 6096 23418 6152 23420
rect 6176 23418 6232 23420
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6096 23366 6142 23418
rect 6142 23366 6152 23418
rect 6176 23366 6206 23418
rect 6206 23366 6218 23418
rect 6218 23366 6232 23418
rect 6256 23366 6270 23418
rect 6270 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6096 23364 6152 23366
rect 6176 23364 6232 23366
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 6096 22330 6152 22332
rect 6176 22330 6232 22332
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6096 22278 6142 22330
rect 6142 22278 6152 22330
rect 6176 22278 6206 22330
rect 6206 22278 6218 22330
rect 6218 22278 6232 22330
rect 6256 22278 6270 22330
rect 6270 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6096 22276 6152 22278
rect 6176 22276 6232 22278
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 6096 21242 6152 21244
rect 6176 21242 6232 21244
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6096 21190 6142 21242
rect 6142 21190 6152 21242
rect 6176 21190 6206 21242
rect 6206 21190 6218 21242
rect 6218 21190 6232 21242
rect 6256 21190 6270 21242
rect 6270 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6096 21188 6152 21190
rect 6176 21188 6232 21190
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 7809 27226 7865 27228
rect 7889 27226 7945 27228
rect 7969 27226 8025 27228
rect 8049 27226 8105 27228
rect 7809 27174 7855 27226
rect 7855 27174 7865 27226
rect 7889 27174 7919 27226
rect 7919 27174 7931 27226
rect 7931 27174 7945 27226
rect 7969 27174 7983 27226
rect 7983 27174 7995 27226
rect 7995 27174 8025 27226
rect 8049 27174 8059 27226
rect 8059 27174 8105 27226
rect 7809 27172 7865 27174
rect 7889 27172 7945 27174
rect 7969 27172 8025 27174
rect 8049 27172 8105 27174
rect 6096 20154 6152 20156
rect 6176 20154 6232 20156
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6096 20102 6142 20154
rect 6142 20102 6152 20154
rect 6176 20102 6206 20154
rect 6206 20102 6218 20154
rect 6218 20102 6232 20154
rect 6256 20102 6270 20154
rect 6270 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6096 20100 6152 20102
rect 6176 20100 6232 20102
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 4618 2524 4620 2544
rect 4620 2524 4672 2544
rect 4672 2524 4674 2544
rect 4618 2488 4674 2524
rect 6096 19066 6152 19068
rect 6176 19066 6232 19068
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6096 19014 6142 19066
rect 6142 19014 6152 19066
rect 6176 19014 6206 19066
rect 6206 19014 6218 19066
rect 6218 19014 6232 19066
rect 6256 19014 6270 19066
rect 6270 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6096 19012 6152 19014
rect 6176 19012 6232 19014
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6096 17978 6152 17980
rect 6176 17978 6232 17980
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6096 17926 6142 17978
rect 6142 17926 6152 17978
rect 6176 17926 6206 17978
rect 6206 17926 6218 17978
rect 6218 17926 6232 17978
rect 6256 17926 6270 17978
rect 6270 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6096 17924 6152 17926
rect 6176 17924 6232 17926
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 7809 26138 7865 26140
rect 7889 26138 7945 26140
rect 7969 26138 8025 26140
rect 8049 26138 8105 26140
rect 7809 26086 7855 26138
rect 7855 26086 7865 26138
rect 7889 26086 7919 26138
rect 7919 26086 7931 26138
rect 7931 26086 7945 26138
rect 7969 26086 7983 26138
rect 7983 26086 7995 26138
rect 7995 26086 8025 26138
rect 8049 26086 8059 26138
rect 8059 26086 8105 26138
rect 7809 26084 7865 26086
rect 7889 26084 7945 26086
rect 7969 26084 8025 26086
rect 8049 26084 8105 26086
rect 7809 25050 7865 25052
rect 7889 25050 7945 25052
rect 7969 25050 8025 25052
rect 8049 25050 8105 25052
rect 7809 24998 7855 25050
rect 7855 24998 7865 25050
rect 7889 24998 7919 25050
rect 7919 24998 7931 25050
rect 7931 24998 7945 25050
rect 7969 24998 7983 25050
rect 7983 24998 7995 25050
rect 7995 24998 8025 25050
rect 8049 24998 8059 25050
rect 8059 24998 8105 25050
rect 7809 24996 7865 24998
rect 7889 24996 7945 24998
rect 7969 24996 8025 24998
rect 8049 24996 8105 24998
rect 7809 23962 7865 23964
rect 7889 23962 7945 23964
rect 7969 23962 8025 23964
rect 8049 23962 8105 23964
rect 7809 23910 7855 23962
rect 7855 23910 7865 23962
rect 7889 23910 7919 23962
rect 7919 23910 7931 23962
rect 7931 23910 7945 23962
rect 7969 23910 7983 23962
rect 7983 23910 7995 23962
rect 7995 23910 8025 23962
rect 8049 23910 8059 23962
rect 8059 23910 8105 23962
rect 7809 23908 7865 23910
rect 7889 23908 7945 23910
rect 7969 23908 8025 23910
rect 8049 23908 8105 23910
rect 7809 22874 7865 22876
rect 7889 22874 7945 22876
rect 7969 22874 8025 22876
rect 8049 22874 8105 22876
rect 7809 22822 7855 22874
rect 7855 22822 7865 22874
rect 7889 22822 7919 22874
rect 7919 22822 7931 22874
rect 7931 22822 7945 22874
rect 7969 22822 7983 22874
rect 7983 22822 7995 22874
rect 7995 22822 8025 22874
rect 8049 22822 8059 22874
rect 8059 22822 8105 22874
rect 7809 22820 7865 22822
rect 7889 22820 7945 22822
rect 7969 22820 8025 22822
rect 8049 22820 8105 22822
rect 7809 21786 7865 21788
rect 7889 21786 7945 21788
rect 7969 21786 8025 21788
rect 8049 21786 8105 21788
rect 7809 21734 7855 21786
rect 7855 21734 7865 21786
rect 7889 21734 7919 21786
rect 7919 21734 7931 21786
rect 7931 21734 7945 21786
rect 7969 21734 7983 21786
rect 7983 21734 7995 21786
rect 7995 21734 8025 21786
rect 8049 21734 8059 21786
rect 8059 21734 8105 21786
rect 7809 21732 7865 21734
rect 7889 21732 7945 21734
rect 7969 21732 8025 21734
rect 8049 21732 8105 21734
rect 7809 20698 7865 20700
rect 7889 20698 7945 20700
rect 7969 20698 8025 20700
rect 8049 20698 8105 20700
rect 7809 20646 7855 20698
rect 7855 20646 7865 20698
rect 7889 20646 7919 20698
rect 7919 20646 7931 20698
rect 7931 20646 7945 20698
rect 7969 20646 7983 20698
rect 7983 20646 7995 20698
rect 7995 20646 8025 20698
rect 8049 20646 8059 20698
rect 8059 20646 8105 20698
rect 7809 20644 7865 20646
rect 7889 20644 7945 20646
rect 7969 20644 8025 20646
rect 8049 20644 8105 20646
rect 7809 19610 7865 19612
rect 7889 19610 7945 19612
rect 7969 19610 8025 19612
rect 8049 19610 8105 19612
rect 7809 19558 7855 19610
rect 7855 19558 7865 19610
rect 7889 19558 7919 19610
rect 7919 19558 7931 19610
rect 7931 19558 7945 19610
rect 7969 19558 7983 19610
rect 7983 19558 7995 19610
rect 7995 19558 8025 19610
rect 8049 19558 8059 19610
rect 8059 19558 8105 19610
rect 7809 19556 7865 19558
rect 7889 19556 7945 19558
rect 7969 19556 8025 19558
rect 8049 19556 8105 19558
rect 7809 18522 7865 18524
rect 7889 18522 7945 18524
rect 7969 18522 8025 18524
rect 8049 18522 8105 18524
rect 7809 18470 7855 18522
rect 7855 18470 7865 18522
rect 7889 18470 7919 18522
rect 7919 18470 7931 18522
rect 7931 18470 7945 18522
rect 7969 18470 7983 18522
rect 7983 18470 7995 18522
rect 7995 18470 8025 18522
rect 8049 18470 8059 18522
rect 8059 18470 8105 18522
rect 7809 18468 7865 18470
rect 7889 18468 7945 18470
rect 7969 18468 8025 18470
rect 8049 18468 8105 18470
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 9523 27770 9579 27772
rect 9603 27770 9659 27772
rect 9683 27770 9739 27772
rect 9763 27770 9819 27772
rect 9523 27718 9569 27770
rect 9569 27718 9579 27770
rect 9603 27718 9633 27770
rect 9633 27718 9645 27770
rect 9645 27718 9659 27770
rect 9683 27718 9697 27770
rect 9697 27718 9709 27770
rect 9709 27718 9739 27770
rect 9763 27718 9773 27770
rect 9773 27718 9819 27770
rect 9523 27716 9579 27718
rect 9603 27716 9659 27718
rect 9683 27716 9739 27718
rect 9763 27716 9819 27718
rect 9523 26682 9579 26684
rect 9603 26682 9659 26684
rect 9683 26682 9739 26684
rect 9763 26682 9819 26684
rect 9523 26630 9569 26682
rect 9569 26630 9579 26682
rect 9603 26630 9633 26682
rect 9633 26630 9645 26682
rect 9645 26630 9659 26682
rect 9683 26630 9697 26682
rect 9697 26630 9709 26682
rect 9709 26630 9739 26682
rect 9763 26630 9773 26682
rect 9773 26630 9819 26682
rect 9523 26628 9579 26630
rect 9603 26628 9659 26630
rect 9683 26628 9739 26630
rect 9763 26628 9819 26630
rect 11236 27226 11292 27228
rect 11316 27226 11372 27228
rect 11396 27226 11452 27228
rect 11476 27226 11532 27228
rect 11236 27174 11282 27226
rect 11282 27174 11292 27226
rect 11316 27174 11346 27226
rect 11346 27174 11358 27226
rect 11358 27174 11372 27226
rect 11396 27174 11410 27226
rect 11410 27174 11422 27226
rect 11422 27174 11452 27226
rect 11476 27174 11486 27226
rect 11486 27174 11532 27226
rect 11236 27172 11292 27174
rect 11316 27172 11372 27174
rect 11396 27172 11452 27174
rect 11476 27172 11532 27174
rect 9523 25594 9579 25596
rect 9603 25594 9659 25596
rect 9683 25594 9739 25596
rect 9763 25594 9819 25596
rect 9523 25542 9569 25594
rect 9569 25542 9579 25594
rect 9603 25542 9633 25594
rect 9633 25542 9645 25594
rect 9645 25542 9659 25594
rect 9683 25542 9697 25594
rect 9697 25542 9709 25594
rect 9709 25542 9739 25594
rect 9763 25542 9773 25594
rect 9773 25542 9819 25594
rect 9523 25540 9579 25542
rect 9603 25540 9659 25542
rect 9683 25540 9739 25542
rect 9763 25540 9819 25542
rect 9523 24506 9579 24508
rect 9603 24506 9659 24508
rect 9683 24506 9739 24508
rect 9763 24506 9819 24508
rect 9523 24454 9569 24506
rect 9569 24454 9579 24506
rect 9603 24454 9633 24506
rect 9633 24454 9645 24506
rect 9645 24454 9659 24506
rect 9683 24454 9697 24506
rect 9697 24454 9709 24506
rect 9709 24454 9739 24506
rect 9763 24454 9773 24506
rect 9773 24454 9819 24506
rect 9523 24452 9579 24454
rect 9603 24452 9659 24454
rect 9683 24452 9739 24454
rect 9763 24452 9819 24454
rect 9523 23418 9579 23420
rect 9603 23418 9659 23420
rect 9683 23418 9739 23420
rect 9763 23418 9819 23420
rect 9523 23366 9569 23418
rect 9569 23366 9579 23418
rect 9603 23366 9633 23418
rect 9633 23366 9645 23418
rect 9645 23366 9659 23418
rect 9683 23366 9697 23418
rect 9697 23366 9709 23418
rect 9709 23366 9739 23418
rect 9763 23366 9773 23418
rect 9773 23366 9819 23418
rect 9523 23364 9579 23366
rect 9603 23364 9659 23366
rect 9683 23364 9739 23366
rect 9763 23364 9819 23366
rect 9523 22330 9579 22332
rect 9603 22330 9659 22332
rect 9683 22330 9739 22332
rect 9763 22330 9819 22332
rect 9523 22278 9569 22330
rect 9569 22278 9579 22330
rect 9603 22278 9633 22330
rect 9633 22278 9645 22330
rect 9645 22278 9659 22330
rect 9683 22278 9697 22330
rect 9697 22278 9709 22330
rect 9709 22278 9739 22330
rect 9763 22278 9773 22330
rect 9773 22278 9819 22330
rect 9523 22276 9579 22278
rect 9603 22276 9659 22278
rect 9683 22276 9739 22278
rect 9763 22276 9819 22278
rect 9523 21242 9579 21244
rect 9603 21242 9659 21244
rect 9683 21242 9739 21244
rect 9763 21242 9819 21244
rect 9523 21190 9569 21242
rect 9569 21190 9579 21242
rect 9603 21190 9633 21242
rect 9633 21190 9645 21242
rect 9645 21190 9659 21242
rect 9683 21190 9697 21242
rect 9697 21190 9709 21242
rect 9709 21190 9739 21242
rect 9763 21190 9773 21242
rect 9773 21190 9819 21242
rect 9523 21188 9579 21190
rect 9603 21188 9659 21190
rect 9683 21188 9739 21190
rect 9763 21188 9819 21190
rect 9523 20154 9579 20156
rect 9603 20154 9659 20156
rect 9683 20154 9739 20156
rect 9763 20154 9819 20156
rect 9523 20102 9569 20154
rect 9569 20102 9579 20154
rect 9603 20102 9633 20154
rect 9633 20102 9645 20154
rect 9645 20102 9659 20154
rect 9683 20102 9697 20154
rect 9697 20102 9709 20154
rect 9709 20102 9739 20154
rect 9763 20102 9773 20154
rect 9773 20102 9819 20154
rect 9523 20100 9579 20102
rect 9603 20100 9659 20102
rect 9683 20100 9739 20102
rect 9763 20100 9819 20102
rect 9523 19066 9579 19068
rect 9603 19066 9659 19068
rect 9683 19066 9739 19068
rect 9763 19066 9819 19068
rect 9523 19014 9569 19066
rect 9569 19014 9579 19066
rect 9603 19014 9633 19066
rect 9633 19014 9645 19066
rect 9645 19014 9659 19066
rect 9683 19014 9697 19066
rect 9697 19014 9709 19066
rect 9709 19014 9739 19066
rect 9763 19014 9773 19066
rect 9773 19014 9819 19066
rect 9523 19012 9579 19014
rect 9603 19012 9659 19014
rect 9683 19012 9739 19014
rect 9763 19012 9819 19014
rect 9523 17978 9579 17980
rect 9603 17978 9659 17980
rect 9683 17978 9739 17980
rect 9763 17978 9819 17980
rect 9523 17926 9569 17978
rect 9569 17926 9579 17978
rect 9603 17926 9633 17978
rect 9633 17926 9645 17978
rect 9645 17926 9659 17978
rect 9683 17926 9697 17978
rect 9697 17926 9709 17978
rect 9709 17926 9739 17978
rect 9763 17926 9773 17978
rect 9773 17926 9819 17978
rect 9523 17924 9579 17926
rect 9603 17924 9659 17926
rect 9683 17924 9739 17926
rect 9763 17924 9819 17926
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 7930 11076 7986 11112
rect 7930 11056 7932 11076
rect 7932 11056 7984 11076
rect 7984 11056 7986 11076
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7102 5072 7158 5128
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 7286 5072 7342 5128
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 11236 26138 11292 26140
rect 11316 26138 11372 26140
rect 11396 26138 11452 26140
rect 11476 26138 11532 26140
rect 11236 26086 11282 26138
rect 11282 26086 11292 26138
rect 11316 26086 11346 26138
rect 11346 26086 11358 26138
rect 11358 26086 11372 26138
rect 11396 26086 11410 26138
rect 11410 26086 11422 26138
rect 11422 26086 11452 26138
rect 11476 26086 11486 26138
rect 11486 26086 11532 26138
rect 11236 26084 11292 26086
rect 11316 26084 11372 26086
rect 11396 26084 11452 26086
rect 11476 26084 11532 26086
rect 10874 25200 10930 25256
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 25050 11292 25052
rect 11316 25050 11372 25052
rect 11396 25050 11452 25052
rect 11476 25050 11532 25052
rect 11236 24998 11282 25050
rect 11282 24998 11292 25050
rect 11316 24998 11346 25050
rect 11346 24998 11358 25050
rect 11358 24998 11372 25050
rect 11396 24998 11410 25050
rect 11410 24998 11422 25050
rect 11422 24998 11452 25050
rect 11476 24998 11486 25050
rect 11486 24998 11532 25050
rect 11236 24996 11292 24998
rect 11316 24996 11372 24998
rect 11396 24996 11452 24998
rect 11476 24996 11532 24998
rect 11236 23962 11292 23964
rect 11316 23962 11372 23964
rect 11396 23962 11452 23964
rect 11476 23962 11532 23964
rect 11236 23910 11282 23962
rect 11282 23910 11292 23962
rect 11316 23910 11346 23962
rect 11346 23910 11358 23962
rect 11358 23910 11372 23962
rect 11396 23910 11410 23962
rect 11410 23910 11422 23962
rect 11422 23910 11452 23962
rect 11476 23910 11486 23962
rect 11486 23910 11532 23962
rect 11236 23908 11292 23910
rect 11316 23908 11372 23910
rect 11396 23908 11452 23910
rect 11476 23908 11532 23910
rect 11236 22874 11292 22876
rect 11316 22874 11372 22876
rect 11396 22874 11452 22876
rect 11476 22874 11532 22876
rect 11236 22822 11282 22874
rect 11282 22822 11292 22874
rect 11316 22822 11346 22874
rect 11346 22822 11358 22874
rect 11358 22822 11372 22874
rect 11396 22822 11410 22874
rect 11410 22822 11422 22874
rect 11422 22822 11452 22874
rect 11476 22822 11486 22874
rect 11486 22822 11532 22874
rect 11236 22820 11292 22822
rect 11316 22820 11372 22822
rect 11396 22820 11452 22822
rect 11476 22820 11532 22822
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11396 21786 11452 21788
rect 11476 21786 11532 21788
rect 11236 21734 11282 21786
rect 11282 21734 11292 21786
rect 11316 21734 11346 21786
rect 11346 21734 11358 21786
rect 11358 21734 11372 21786
rect 11396 21734 11410 21786
rect 11410 21734 11422 21786
rect 11422 21734 11452 21786
rect 11476 21734 11486 21786
rect 11486 21734 11532 21786
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11396 21732 11452 21734
rect 11476 21732 11532 21734
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11396 20698 11452 20700
rect 11476 20698 11532 20700
rect 11236 20646 11282 20698
rect 11282 20646 11292 20698
rect 11316 20646 11346 20698
rect 11346 20646 11358 20698
rect 11358 20646 11372 20698
rect 11396 20646 11410 20698
rect 11410 20646 11422 20698
rect 11422 20646 11452 20698
rect 11476 20646 11486 20698
rect 11486 20646 11532 20698
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11396 20644 11452 20646
rect 11476 20644 11532 20646
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11396 19610 11452 19612
rect 11476 19610 11532 19612
rect 11236 19558 11282 19610
rect 11282 19558 11292 19610
rect 11316 19558 11346 19610
rect 11346 19558 11358 19610
rect 11358 19558 11372 19610
rect 11396 19558 11410 19610
rect 11410 19558 11422 19610
rect 11422 19558 11452 19610
rect 11476 19558 11486 19610
rect 11486 19558 11532 19610
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 11396 19556 11452 19558
rect 11476 19556 11532 19558
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11396 18522 11452 18524
rect 11476 18522 11532 18524
rect 11236 18470 11282 18522
rect 11282 18470 11292 18522
rect 11316 18470 11346 18522
rect 11346 18470 11358 18522
rect 11358 18470 11372 18522
rect 11396 18470 11410 18522
rect 11410 18470 11422 18522
rect 11422 18470 11452 18522
rect 11476 18470 11486 18522
rect 11486 18470 11532 18522
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11396 18468 11452 18470
rect 11476 18468 11532 18470
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 12530 25200 12586 25256
rect 12950 27770 13006 27772
rect 13030 27770 13086 27772
rect 13110 27770 13166 27772
rect 13190 27770 13246 27772
rect 12950 27718 12996 27770
rect 12996 27718 13006 27770
rect 13030 27718 13060 27770
rect 13060 27718 13072 27770
rect 13072 27718 13086 27770
rect 13110 27718 13124 27770
rect 13124 27718 13136 27770
rect 13136 27718 13166 27770
rect 13190 27718 13200 27770
rect 13200 27718 13246 27770
rect 12950 27716 13006 27718
rect 13030 27716 13086 27718
rect 13110 27716 13166 27718
rect 13190 27716 13246 27718
rect 12950 26682 13006 26684
rect 13030 26682 13086 26684
rect 13110 26682 13166 26684
rect 13190 26682 13246 26684
rect 12950 26630 12996 26682
rect 12996 26630 13006 26682
rect 13030 26630 13060 26682
rect 13060 26630 13072 26682
rect 13072 26630 13086 26682
rect 13110 26630 13124 26682
rect 13124 26630 13136 26682
rect 13136 26630 13166 26682
rect 13190 26630 13200 26682
rect 13200 26630 13246 26682
rect 12950 26628 13006 26630
rect 13030 26628 13086 26630
rect 13110 26628 13166 26630
rect 13190 26628 13246 26630
rect 12950 25594 13006 25596
rect 13030 25594 13086 25596
rect 13110 25594 13166 25596
rect 13190 25594 13246 25596
rect 12950 25542 12996 25594
rect 12996 25542 13006 25594
rect 13030 25542 13060 25594
rect 13060 25542 13072 25594
rect 13072 25542 13086 25594
rect 13110 25542 13124 25594
rect 13124 25542 13136 25594
rect 13136 25542 13166 25594
rect 13190 25542 13200 25594
rect 13200 25542 13246 25594
rect 12950 25540 13006 25542
rect 13030 25540 13086 25542
rect 13110 25540 13166 25542
rect 13190 25540 13246 25542
rect 12950 24506 13006 24508
rect 13030 24506 13086 24508
rect 13110 24506 13166 24508
rect 13190 24506 13246 24508
rect 12950 24454 12996 24506
rect 12996 24454 13006 24506
rect 13030 24454 13060 24506
rect 13060 24454 13072 24506
rect 13072 24454 13086 24506
rect 13110 24454 13124 24506
rect 13124 24454 13136 24506
rect 13136 24454 13166 24506
rect 13190 24454 13200 24506
rect 13200 24454 13246 24506
rect 12950 24452 13006 24454
rect 13030 24452 13086 24454
rect 13110 24452 13166 24454
rect 13190 24452 13246 24454
rect 14663 27226 14719 27228
rect 14743 27226 14799 27228
rect 14823 27226 14879 27228
rect 14903 27226 14959 27228
rect 14663 27174 14709 27226
rect 14709 27174 14719 27226
rect 14743 27174 14773 27226
rect 14773 27174 14785 27226
rect 14785 27174 14799 27226
rect 14823 27174 14837 27226
rect 14837 27174 14849 27226
rect 14849 27174 14879 27226
rect 14903 27174 14913 27226
rect 14913 27174 14959 27226
rect 14663 27172 14719 27174
rect 14743 27172 14799 27174
rect 14823 27172 14879 27174
rect 14903 27172 14959 27174
rect 14663 26138 14719 26140
rect 14743 26138 14799 26140
rect 14823 26138 14879 26140
rect 14903 26138 14959 26140
rect 14663 26086 14709 26138
rect 14709 26086 14719 26138
rect 14743 26086 14773 26138
rect 14773 26086 14785 26138
rect 14785 26086 14799 26138
rect 14823 26086 14837 26138
rect 14837 26086 14849 26138
rect 14849 26086 14879 26138
rect 14903 26086 14913 26138
rect 14913 26086 14959 26138
rect 14663 26084 14719 26086
rect 14743 26084 14799 26086
rect 14823 26084 14879 26086
rect 14903 26084 14959 26086
rect 14663 25050 14719 25052
rect 14743 25050 14799 25052
rect 14823 25050 14879 25052
rect 14903 25050 14959 25052
rect 14663 24998 14709 25050
rect 14709 24998 14719 25050
rect 14743 24998 14773 25050
rect 14773 24998 14785 25050
rect 14785 24998 14799 25050
rect 14823 24998 14837 25050
rect 14837 24998 14849 25050
rect 14849 24998 14879 25050
rect 14903 24998 14913 25050
rect 14913 24998 14959 25050
rect 14663 24996 14719 24998
rect 14743 24996 14799 24998
rect 14823 24996 14879 24998
rect 14903 24996 14959 24998
rect 14663 23962 14719 23964
rect 14743 23962 14799 23964
rect 14823 23962 14879 23964
rect 14903 23962 14959 23964
rect 14663 23910 14709 23962
rect 14709 23910 14719 23962
rect 14743 23910 14773 23962
rect 14773 23910 14785 23962
rect 14785 23910 14799 23962
rect 14823 23910 14837 23962
rect 14837 23910 14849 23962
rect 14849 23910 14879 23962
rect 14903 23910 14913 23962
rect 14913 23910 14959 23962
rect 14663 23908 14719 23910
rect 14743 23908 14799 23910
rect 14823 23908 14879 23910
rect 14903 23908 14959 23910
rect 12950 23418 13006 23420
rect 13030 23418 13086 23420
rect 13110 23418 13166 23420
rect 13190 23418 13246 23420
rect 12950 23366 12996 23418
rect 12996 23366 13006 23418
rect 13030 23366 13060 23418
rect 13060 23366 13072 23418
rect 13072 23366 13086 23418
rect 13110 23366 13124 23418
rect 13124 23366 13136 23418
rect 13136 23366 13166 23418
rect 13190 23366 13200 23418
rect 13200 23366 13246 23418
rect 12950 23364 13006 23366
rect 13030 23364 13086 23366
rect 13110 23364 13166 23366
rect 13190 23364 13246 23366
rect 14663 22874 14719 22876
rect 14743 22874 14799 22876
rect 14823 22874 14879 22876
rect 14903 22874 14959 22876
rect 14663 22822 14709 22874
rect 14709 22822 14719 22874
rect 14743 22822 14773 22874
rect 14773 22822 14785 22874
rect 14785 22822 14799 22874
rect 14823 22822 14837 22874
rect 14837 22822 14849 22874
rect 14849 22822 14879 22874
rect 14903 22822 14913 22874
rect 14913 22822 14959 22874
rect 14663 22820 14719 22822
rect 14743 22820 14799 22822
rect 14823 22820 14879 22822
rect 14903 22820 14959 22822
rect 12950 22330 13006 22332
rect 13030 22330 13086 22332
rect 13110 22330 13166 22332
rect 13190 22330 13246 22332
rect 12950 22278 12996 22330
rect 12996 22278 13006 22330
rect 13030 22278 13060 22330
rect 13060 22278 13072 22330
rect 13072 22278 13086 22330
rect 13110 22278 13124 22330
rect 13124 22278 13136 22330
rect 13136 22278 13166 22330
rect 13190 22278 13200 22330
rect 13200 22278 13246 22330
rect 12950 22276 13006 22278
rect 13030 22276 13086 22278
rect 13110 22276 13166 22278
rect 13190 22276 13246 22278
rect 14663 21786 14719 21788
rect 14743 21786 14799 21788
rect 14823 21786 14879 21788
rect 14903 21786 14959 21788
rect 14663 21734 14709 21786
rect 14709 21734 14719 21786
rect 14743 21734 14773 21786
rect 14773 21734 14785 21786
rect 14785 21734 14799 21786
rect 14823 21734 14837 21786
rect 14837 21734 14849 21786
rect 14849 21734 14879 21786
rect 14903 21734 14913 21786
rect 14913 21734 14959 21786
rect 14663 21732 14719 21734
rect 14743 21732 14799 21734
rect 14823 21732 14879 21734
rect 14903 21732 14959 21734
rect 12950 21242 13006 21244
rect 13030 21242 13086 21244
rect 13110 21242 13166 21244
rect 13190 21242 13246 21244
rect 12950 21190 12996 21242
rect 12996 21190 13006 21242
rect 13030 21190 13060 21242
rect 13060 21190 13072 21242
rect 13072 21190 13086 21242
rect 13110 21190 13124 21242
rect 13124 21190 13136 21242
rect 13136 21190 13166 21242
rect 13190 21190 13200 21242
rect 13200 21190 13246 21242
rect 12950 21188 13006 21190
rect 13030 21188 13086 21190
rect 13110 21188 13166 21190
rect 13190 21188 13246 21190
rect 14663 20698 14719 20700
rect 14743 20698 14799 20700
rect 14823 20698 14879 20700
rect 14903 20698 14959 20700
rect 14663 20646 14709 20698
rect 14709 20646 14719 20698
rect 14743 20646 14773 20698
rect 14773 20646 14785 20698
rect 14785 20646 14799 20698
rect 14823 20646 14837 20698
rect 14837 20646 14849 20698
rect 14849 20646 14879 20698
rect 14903 20646 14913 20698
rect 14913 20646 14959 20698
rect 14663 20644 14719 20646
rect 14743 20644 14799 20646
rect 14823 20644 14879 20646
rect 14903 20644 14959 20646
rect 12950 20154 13006 20156
rect 13030 20154 13086 20156
rect 13110 20154 13166 20156
rect 13190 20154 13246 20156
rect 12950 20102 12996 20154
rect 12996 20102 13006 20154
rect 13030 20102 13060 20154
rect 13060 20102 13072 20154
rect 13072 20102 13086 20154
rect 13110 20102 13124 20154
rect 13124 20102 13136 20154
rect 13136 20102 13166 20154
rect 13190 20102 13200 20154
rect 13200 20102 13246 20154
rect 12950 20100 13006 20102
rect 13030 20100 13086 20102
rect 13110 20100 13166 20102
rect 13190 20100 13246 20102
rect 14663 19610 14719 19612
rect 14743 19610 14799 19612
rect 14823 19610 14879 19612
rect 14903 19610 14959 19612
rect 14663 19558 14709 19610
rect 14709 19558 14719 19610
rect 14743 19558 14773 19610
rect 14773 19558 14785 19610
rect 14785 19558 14799 19610
rect 14823 19558 14837 19610
rect 14837 19558 14849 19610
rect 14849 19558 14879 19610
rect 14903 19558 14913 19610
rect 14913 19558 14959 19610
rect 14663 19556 14719 19558
rect 14743 19556 14799 19558
rect 14823 19556 14879 19558
rect 14903 19556 14959 19558
rect 12950 19066 13006 19068
rect 13030 19066 13086 19068
rect 13110 19066 13166 19068
rect 13190 19066 13246 19068
rect 12950 19014 12996 19066
rect 12996 19014 13006 19066
rect 13030 19014 13060 19066
rect 13060 19014 13072 19066
rect 13072 19014 13086 19066
rect 13110 19014 13124 19066
rect 13124 19014 13136 19066
rect 13136 19014 13166 19066
rect 13190 19014 13200 19066
rect 13200 19014 13246 19066
rect 12950 19012 13006 19014
rect 13030 19012 13086 19014
rect 13110 19012 13166 19014
rect 13190 19012 13246 19014
rect 14663 18522 14719 18524
rect 14743 18522 14799 18524
rect 14823 18522 14879 18524
rect 14903 18522 14959 18524
rect 14663 18470 14709 18522
rect 14709 18470 14719 18522
rect 14743 18470 14773 18522
rect 14773 18470 14785 18522
rect 14785 18470 14799 18522
rect 14823 18470 14837 18522
rect 14837 18470 14849 18522
rect 14849 18470 14879 18522
rect 14903 18470 14913 18522
rect 14913 18470 14959 18522
rect 14663 18468 14719 18470
rect 14743 18468 14799 18470
rect 14823 18468 14879 18470
rect 14903 18468 14959 18470
rect 12950 17978 13006 17980
rect 13030 17978 13086 17980
rect 13110 17978 13166 17980
rect 13190 17978 13246 17980
rect 12950 17926 12996 17978
rect 12996 17926 13006 17978
rect 13030 17926 13060 17978
rect 13060 17926 13072 17978
rect 13072 17926 13086 17978
rect 13110 17926 13124 17978
rect 13124 17926 13136 17978
rect 13136 17926 13166 17978
rect 13190 17926 13200 17978
rect 13200 17926 13246 17978
rect 12950 17924 13006 17926
rect 13030 17924 13086 17926
rect 13110 17924 13166 17926
rect 13190 17924 13246 17926
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
<< metal3 >>
rect 2659 27776 2975 27777
rect 2659 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2975 27776
rect 2659 27711 2975 27712
rect 6086 27776 6402 27777
rect 6086 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6402 27776
rect 6086 27711 6402 27712
rect 9513 27776 9829 27777
rect 9513 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9829 27776
rect 9513 27711 9829 27712
rect 12940 27776 13256 27777
rect 12940 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13256 27776
rect 12940 27711 13256 27712
rect 4372 27232 4688 27233
rect 4372 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4688 27232
rect 4372 27167 4688 27168
rect 7799 27232 8115 27233
rect 7799 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8115 27232
rect 7799 27167 8115 27168
rect 11226 27232 11542 27233
rect 11226 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11542 27232
rect 11226 27167 11542 27168
rect 14653 27232 14969 27233
rect 14653 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14969 27232
rect 14653 27167 14969 27168
rect 2659 26688 2975 26689
rect 2659 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2975 26688
rect 2659 26623 2975 26624
rect 6086 26688 6402 26689
rect 6086 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6402 26688
rect 6086 26623 6402 26624
rect 9513 26688 9829 26689
rect 9513 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9829 26688
rect 9513 26623 9829 26624
rect 12940 26688 13256 26689
rect 12940 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13256 26688
rect 12940 26623 13256 26624
rect 4372 26144 4688 26145
rect 4372 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4688 26144
rect 4372 26079 4688 26080
rect 7799 26144 8115 26145
rect 7799 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8115 26144
rect 7799 26079 8115 26080
rect 11226 26144 11542 26145
rect 11226 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11542 26144
rect 11226 26079 11542 26080
rect 14653 26144 14969 26145
rect 14653 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14969 26144
rect 14653 26079 14969 26080
rect 2659 25600 2975 25601
rect 2659 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2975 25600
rect 2659 25535 2975 25536
rect 6086 25600 6402 25601
rect 6086 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6402 25600
rect 6086 25535 6402 25536
rect 9513 25600 9829 25601
rect 9513 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9829 25600
rect 9513 25535 9829 25536
rect 12940 25600 13256 25601
rect 12940 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13256 25600
rect 12940 25535 13256 25536
rect 10869 25258 10935 25261
rect 12525 25258 12591 25261
rect 10869 25256 12591 25258
rect 10869 25200 10874 25256
rect 10930 25200 12530 25256
rect 12586 25200 12591 25256
rect 10869 25198 12591 25200
rect 10869 25195 10935 25198
rect 12525 25195 12591 25198
rect 4372 25056 4688 25057
rect 4372 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4688 25056
rect 4372 24991 4688 24992
rect 7799 25056 8115 25057
rect 7799 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8115 25056
rect 7799 24991 8115 24992
rect 11226 25056 11542 25057
rect 11226 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11542 25056
rect 11226 24991 11542 24992
rect 14653 25056 14969 25057
rect 14653 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14969 25056
rect 14653 24991 14969 24992
rect 2659 24512 2975 24513
rect 2659 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2975 24512
rect 2659 24447 2975 24448
rect 6086 24512 6402 24513
rect 6086 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6402 24512
rect 6086 24447 6402 24448
rect 9513 24512 9829 24513
rect 9513 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9829 24512
rect 9513 24447 9829 24448
rect 12940 24512 13256 24513
rect 12940 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13256 24512
rect 12940 24447 13256 24448
rect 4372 23968 4688 23969
rect 4372 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4688 23968
rect 4372 23903 4688 23904
rect 7799 23968 8115 23969
rect 7799 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8115 23968
rect 7799 23903 8115 23904
rect 11226 23968 11542 23969
rect 11226 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11542 23968
rect 11226 23903 11542 23904
rect 14653 23968 14969 23969
rect 14653 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14969 23968
rect 14653 23903 14969 23904
rect 2659 23424 2975 23425
rect 2659 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2975 23424
rect 2659 23359 2975 23360
rect 6086 23424 6402 23425
rect 6086 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6402 23424
rect 6086 23359 6402 23360
rect 9513 23424 9829 23425
rect 9513 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9829 23424
rect 9513 23359 9829 23360
rect 12940 23424 13256 23425
rect 12940 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13256 23424
rect 12940 23359 13256 23360
rect 4372 22880 4688 22881
rect 4372 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4688 22880
rect 4372 22815 4688 22816
rect 7799 22880 8115 22881
rect 7799 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8115 22880
rect 7799 22815 8115 22816
rect 11226 22880 11542 22881
rect 11226 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11542 22880
rect 11226 22815 11542 22816
rect 14653 22880 14969 22881
rect 14653 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14969 22880
rect 14653 22815 14969 22816
rect 2659 22336 2975 22337
rect 2659 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2975 22336
rect 2659 22271 2975 22272
rect 6086 22336 6402 22337
rect 6086 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6402 22336
rect 6086 22271 6402 22272
rect 9513 22336 9829 22337
rect 9513 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9829 22336
rect 9513 22271 9829 22272
rect 12940 22336 13256 22337
rect 12940 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13256 22336
rect 12940 22271 13256 22272
rect 4372 21792 4688 21793
rect 4372 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4688 21792
rect 4372 21727 4688 21728
rect 7799 21792 8115 21793
rect 7799 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8115 21792
rect 7799 21727 8115 21728
rect 11226 21792 11542 21793
rect 11226 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11542 21792
rect 11226 21727 11542 21728
rect 14653 21792 14969 21793
rect 14653 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14969 21792
rect 14653 21727 14969 21728
rect 2659 21248 2975 21249
rect 2659 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2975 21248
rect 2659 21183 2975 21184
rect 6086 21248 6402 21249
rect 6086 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6402 21248
rect 6086 21183 6402 21184
rect 9513 21248 9829 21249
rect 9513 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9829 21248
rect 9513 21183 9829 21184
rect 12940 21248 13256 21249
rect 12940 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13256 21248
rect 12940 21183 13256 21184
rect 4372 20704 4688 20705
rect 4372 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4688 20704
rect 4372 20639 4688 20640
rect 7799 20704 8115 20705
rect 7799 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8115 20704
rect 7799 20639 8115 20640
rect 11226 20704 11542 20705
rect 11226 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11542 20704
rect 11226 20639 11542 20640
rect 14653 20704 14969 20705
rect 14653 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14969 20704
rect 14653 20639 14969 20640
rect 2659 20160 2975 20161
rect 2659 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2975 20160
rect 2659 20095 2975 20096
rect 6086 20160 6402 20161
rect 6086 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6402 20160
rect 6086 20095 6402 20096
rect 9513 20160 9829 20161
rect 9513 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9829 20160
rect 9513 20095 9829 20096
rect 12940 20160 13256 20161
rect 12940 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13256 20160
rect 12940 20095 13256 20096
rect 4372 19616 4688 19617
rect 4372 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4688 19616
rect 4372 19551 4688 19552
rect 7799 19616 8115 19617
rect 7799 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8115 19616
rect 7799 19551 8115 19552
rect 11226 19616 11542 19617
rect 11226 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11542 19616
rect 11226 19551 11542 19552
rect 14653 19616 14969 19617
rect 14653 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14969 19616
rect 14653 19551 14969 19552
rect 2659 19072 2975 19073
rect 2659 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2975 19072
rect 2659 19007 2975 19008
rect 6086 19072 6402 19073
rect 6086 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6402 19072
rect 6086 19007 6402 19008
rect 9513 19072 9829 19073
rect 9513 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9829 19072
rect 9513 19007 9829 19008
rect 12940 19072 13256 19073
rect 12940 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13256 19072
rect 12940 19007 13256 19008
rect 4372 18528 4688 18529
rect 4372 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4688 18528
rect 4372 18463 4688 18464
rect 7799 18528 8115 18529
rect 7799 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8115 18528
rect 7799 18463 8115 18464
rect 11226 18528 11542 18529
rect 11226 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11542 18528
rect 11226 18463 11542 18464
rect 14653 18528 14969 18529
rect 14653 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14969 18528
rect 14653 18463 14969 18464
rect 2659 17984 2975 17985
rect 2659 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2975 17984
rect 2659 17919 2975 17920
rect 6086 17984 6402 17985
rect 6086 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6402 17984
rect 6086 17919 6402 17920
rect 9513 17984 9829 17985
rect 9513 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9829 17984
rect 9513 17919 9829 17920
rect 12940 17984 13256 17985
rect 12940 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13256 17984
rect 12940 17919 13256 17920
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 12940 16831 13256 16832
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 14653 15199 14969 15200
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 14653 11935 14969 11936
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 7414 11052 7420 11116
rect 7484 11114 7490 11116
rect 7925 11114 7991 11117
rect 7484 11112 7991 11114
rect 7484 11056 7930 11112
rect 7986 11056 7991 11112
rect 7484 11054 7991 11056
rect 7484 11052 7490 11054
rect 7925 11051 7991 11054
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 12940 7039 13256 7040
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 7097 5130 7163 5133
rect 7281 5130 7347 5133
rect 7097 5128 7347 5130
rect 7097 5072 7102 5128
rect 7158 5072 7286 5128
rect 7342 5072 7347 5128
rect 7097 5070 7347 5072
rect 7097 5067 7163 5070
rect 7281 5067 7347 5070
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 4613 2546 4679 2549
rect 7414 2546 7420 2548
rect 4613 2544 7420 2546
rect 4613 2488 4618 2544
rect 4674 2488 7420 2544
rect 4613 2486 7420 2488
rect 4613 2483 4679 2486
rect 7414 2484 7420 2486
rect 7484 2484 7490 2548
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
<< via3 >>
rect 2665 27772 2729 27776
rect 2665 27716 2669 27772
rect 2669 27716 2725 27772
rect 2725 27716 2729 27772
rect 2665 27712 2729 27716
rect 2745 27772 2809 27776
rect 2745 27716 2749 27772
rect 2749 27716 2805 27772
rect 2805 27716 2809 27772
rect 2745 27712 2809 27716
rect 2825 27772 2889 27776
rect 2825 27716 2829 27772
rect 2829 27716 2885 27772
rect 2885 27716 2889 27772
rect 2825 27712 2889 27716
rect 2905 27772 2969 27776
rect 2905 27716 2909 27772
rect 2909 27716 2965 27772
rect 2965 27716 2969 27772
rect 2905 27712 2969 27716
rect 6092 27772 6156 27776
rect 6092 27716 6096 27772
rect 6096 27716 6152 27772
rect 6152 27716 6156 27772
rect 6092 27712 6156 27716
rect 6172 27772 6236 27776
rect 6172 27716 6176 27772
rect 6176 27716 6232 27772
rect 6232 27716 6236 27772
rect 6172 27712 6236 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 9519 27772 9583 27776
rect 9519 27716 9523 27772
rect 9523 27716 9579 27772
rect 9579 27716 9583 27772
rect 9519 27712 9583 27716
rect 9599 27772 9663 27776
rect 9599 27716 9603 27772
rect 9603 27716 9659 27772
rect 9659 27716 9663 27772
rect 9599 27712 9663 27716
rect 9679 27772 9743 27776
rect 9679 27716 9683 27772
rect 9683 27716 9739 27772
rect 9739 27716 9743 27772
rect 9679 27712 9743 27716
rect 9759 27772 9823 27776
rect 9759 27716 9763 27772
rect 9763 27716 9819 27772
rect 9819 27716 9823 27772
rect 9759 27712 9823 27716
rect 12946 27772 13010 27776
rect 12946 27716 12950 27772
rect 12950 27716 13006 27772
rect 13006 27716 13010 27772
rect 12946 27712 13010 27716
rect 13026 27772 13090 27776
rect 13026 27716 13030 27772
rect 13030 27716 13086 27772
rect 13086 27716 13090 27772
rect 13026 27712 13090 27716
rect 13106 27772 13170 27776
rect 13106 27716 13110 27772
rect 13110 27716 13166 27772
rect 13166 27716 13170 27772
rect 13106 27712 13170 27716
rect 13186 27772 13250 27776
rect 13186 27716 13190 27772
rect 13190 27716 13246 27772
rect 13246 27716 13250 27772
rect 13186 27712 13250 27716
rect 4378 27228 4442 27232
rect 4378 27172 4382 27228
rect 4382 27172 4438 27228
rect 4438 27172 4442 27228
rect 4378 27168 4442 27172
rect 4458 27228 4522 27232
rect 4458 27172 4462 27228
rect 4462 27172 4518 27228
rect 4518 27172 4522 27228
rect 4458 27168 4522 27172
rect 4538 27228 4602 27232
rect 4538 27172 4542 27228
rect 4542 27172 4598 27228
rect 4598 27172 4602 27228
rect 4538 27168 4602 27172
rect 4618 27228 4682 27232
rect 4618 27172 4622 27228
rect 4622 27172 4678 27228
rect 4678 27172 4682 27228
rect 4618 27168 4682 27172
rect 7805 27228 7869 27232
rect 7805 27172 7809 27228
rect 7809 27172 7865 27228
rect 7865 27172 7869 27228
rect 7805 27168 7869 27172
rect 7885 27228 7949 27232
rect 7885 27172 7889 27228
rect 7889 27172 7945 27228
rect 7945 27172 7949 27228
rect 7885 27168 7949 27172
rect 7965 27228 8029 27232
rect 7965 27172 7969 27228
rect 7969 27172 8025 27228
rect 8025 27172 8029 27228
rect 7965 27168 8029 27172
rect 8045 27228 8109 27232
rect 8045 27172 8049 27228
rect 8049 27172 8105 27228
rect 8105 27172 8109 27228
rect 8045 27168 8109 27172
rect 11232 27228 11296 27232
rect 11232 27172 11236 27228
rect 11236 27172 11292 27228
rect 11292 27172 11296 27228
rect 11232 27168 11296 27172
rect 11312 27228 11376 27232
rect 11312 27172 11316 27228
rect 11316 27172 11372 27228
rect 11372 27172 11376 27228
rect 11312 27168 11376 27172
rect 11392 27228 11456 27232
rect 11392 27172 11396 27228
rect 11396 27172 11452 27228
rect 11452 27172 11456 27228
rect 11392 27168 11456 27172
rect 11472 27228 11536 27232
rect 11472 27172 11476 27228
rect 11476 27172 11532 27228
rect 11532 27172 11536 27228
rect 11472 27168 11536 27172
rect 14659 27228 14723 27232
rect 14659 27172 14663 27228
rect 14663 27172 14719 27228
rect 14719 27172 14723 27228
rect 14659 27168 14723 27172
rect 14739 27228 14803 27232
rect 14739 27172 14743 27228
rect 14743 27172 14799 27228
rect 14799 27172 14803 27228
rect 14739 27168 14803 27172
rect 14819 27228 14883 27232
rect 14819 27172 14823 27228
rect 14823 27172 14879 27228
rect 14879 27172 14883 27228
rect 14819 27168 14883 27172
rect 14899 27228 14963 27232
rect 14899 27172 14903 27228
rect 14903 27172 14959 27228
rect 14959 27172 14963 27228
rect 14899 27168 14963 27172
rect 2665 26684 2729 26688
rect 2665 26628 2669 26684
rect 2669 26628 2725 26684
rect 2725 26628 2729 26684
rect 2665 26624 2729 26628
rect 2745 26684 2809 26688
rect 2745 26628 2749 26684
rect 2749 26628 2805 26684
rect 2805 26628 2809 26684
rect 2745 26624 2809 26628
rect 2825 26684 2889 26688
rect 2825 26628 2829 26684
rect 2829 26628 2885 26684
rect 2885 26628 2889 26684
rect 2825 26624 2889 26628
rect 2905 26684 2969 26688
rect 2905 26628 2909 26684
rect 2909 26628 2965 26684
rect 2965 26628 2969 26684
rect 2905 26624 2969 26628
rect 6092 26684 6156 26688
rect 6092 26628 6096 26684
rect 6096 26628 6152 26684
rect 6152 26628 6156 26684
rect 6092 26624 6156 26628
rect 6172 26684 6236 26688
rect 6172 26628 6176 26684
rect 6176 26628 6232 26684
rect 6232 26628 6236 26684
rect 6172 26624 6236 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 9519 26684 9583 26688
rect 9519 26628 9523 26684
rect 9523 26628 9579 26684
rect 9579 26628 9583 26684
rect 9519 26624 9583 26628
rect 9599 26684 9663 26688
rect 9599 26628 9603 26684
rect 9603 26628 9659 26684
rect 9659 26628 9663 26684
rect 9599 26624 9663 26628
rect 9679 26684 9743 26688
rect 9679 26628 9683 26684
rect 9683 26628 9739 26684
rect 9739 26628 9743 26684
rect 9679 26624 9743 26628
rect 9759 26684 9823 26688
rect 9759 26628 9763 26684
rect 9763 26628 9819 26684
rect 9819 26628 9823 26684
rect 9759 26624 9823 26628
rect 12946 26684 13010 26688
rect 12946 26628 12950 26684
rect 12950 26628 13006 26684
rect 13006 26628 13010 26684
rect 12946 26624 13010 26628
rect 13026 26684 13090 26688
rect 13026 26628 13030 26684
rect 13030 26628 13086 26684
rect 13086 26628 13090 26684
rect 13026 26624 13090 26628
rect 13106 26684 13170 26688
rect 13106 26628 13110 26684
rect 13110 26628 13166 26684
rect 13166 26628 13170 26684
rect 13106 26624 13170 26628
rect 13186 26684 13250 26688
rect 13186 26628 13190 26684
rect 13190 26628 13246 26684
rect 13246 26628 13250 26684
rect 13186 26624 13250 26628
rect 4378 26140 4442 26144
rect 4378 26084 4382 26140
rect 4382 26084 4438 26140
rect 4438 26084 4442 26140
rect 4378 26080 4442 26084
rect 4458 26140 4522 26144
rect 4458 26084 4462 26140
rect 4462 26084 4518 26140
rect 4518 26084 4522 26140
rect 4458 26080 4522 26084
rect 4538 26140 4602 26144
rect 4538 26084 4542 26140
rect 4542 26084 4598 26140
rect 4598 26084 4602 26140
rect 4538 26080 4602 26084
rect 4618 26140 4682 26144
rect 4618 26084 4622 26140
rect 4622 26084 4678 26140
rect 4678 26084 4682 26140
rect 4618 26080 4682 26084
rect 7805 26140 7869 26144
rect 7805 26084 7809 26140
rect 7809 26084 7865 26140
rect 7865 26084 7869 26140
rect 7805 26080 7869 26084
rect 7885 26140 7949 26144
rect 7885 26084 7889 26140
rect 7889 26084 7945 26140
rect 7945 26084 7949 26140
rect 7885 26080 7949 26084
rect 7965 26140 8029 26144
rect 7965 26084 7969 26140
rect 7969 26084 8025 26140
rect 8025 26084 8029 26140
rect 7965 26080 8029 26084
rect 8045 26140 8109 26144
rect 8045 26084 8049 26140
rect 8049 26084 8105 26140
rect 8105 26084 8109 26140
rect 8045 26080 8109 26084
rect 11232 26140 11296 26144
rect 11232 26084 11236 26140
rect 11236 26084 11292 26140
rect 11292 26084 11296 26140
rect 11232 26080 11296 26084
rect 11312 26140 11376 26144
rect 11312 26084 11316 26140
rect 11316 26084 11372 26140
rect 11372 26084 11376 26140
rect 11312 26080 11376 26084
rect 11392 26140 11456 26144
rect 11392 26084 11396 26140
rect 11396 26084 11452 26140
rect 11452 26084 11456 26140
rect 11392 26080 11456 26084
rect 11472 26140 11536 26144
rect 11472 26084 11476 26140
rect 11476 26084 11532 26140
rect 11532 26084 11536 26140
rect 11472 26080 11536 26084
rect 14659 26140 14723 26144
rect 14659 26084 14663 26140
rect 14663 26084 14719 26140
rect 14719 26084 14723 26140
rect 14659 26080 14723 26084
rect 14739 26140 14803 26144
rect 14739 26084 14743 26140
rect 14743 26084 14799 26140
rect 14799 26084 14803 26140
rect 14739 26080 14803 26084
rect 14819 26140 14883 26144
rect 14819 26084 14823 26140
rect 14823 26084 14879 26140
rect 14879 26084 14883 26140
rect 14819 26080 14883 26084
rect 14899 26140 14963 26144
rect 14899 26084 14903 26140
rect 14903 26084 14959 26140
rect 14959 26084 14963 26140
rect 14899 26080 14963 26084
rect 2665 25596 2729 25600
rect 2665 25540 2669 25596
rect 2669 25540 2725 25596
rect 2725 25540 2729 25596
rect 2665 25536 2729 25540
rect 2745 25596 2809 25600
rect 2745 25540 2749 25596
rect 2749 25540 2805 25596
rect 2805 25540 2809 25596
rect 2745 25536 2809 25540
rect 2825 25596 2889 25600
rect 2825 25540 2829 25596
rect 2829 25540 2885 25596
rect 2885 25540 2889 25596
rect 2825 25536 2889 25540
rect 2905 25596 2969 25600
rect 2905 25540 2909 25596
rect 2909 25540 2965 25596
rect 2965 25540 2969 25596
rect 2905 25536 2969 25540
rect 6092 25596 6156 25600
rect 6092 25540 6096 25596
rect 6096 25540 6152 25596
rect 6152 25540 6156 25596
rect 6092 25536 6156 25540
rect 6172 25596 6236 25600
rect 6172 25540 6176 25596
rect 6176 25540 6232 25596
rect 6232 25540 6236 25596
rect 6172 25536 6236 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 9519 25596 9583 25600
rect 9519 25540 9523 25596
rect 9523 25540 9579 25596
rect 9579 25540 9583 25596
rect 9519 25536 9583 25540
rect 9599 25596 9663 25600
rect 9599 25540 9603 25596
rect 9603 25540 9659 25596
rect 9659 25540 9663 25596
rect 9599 25536 9663 25540
rect 9679 25596 9743 25600
rect 9679 25540 9683 25596
rect 9683 25540 9739 25596
rect 9739 25540 9743 25596
rect 9679 25536 9743 25540
rect 9759 25596 9823 25600
rect 9759 25540 9763 25596
rect 9763 25540 9819 25596
rect 9819 25540 9823 25596
rect 9759 25536 9823 25540
rect 12946 25596 13010 25600
rect 12946 25540 12950 25596
rect 12950 25540 13006 25596
rect 13006 25540 13010 25596
rect 12946 25536 13010 25540
rect 13026 25596 13090 25600
rect 13026 25540 13030 25596
rect 13030 25540 13086 25596
rect 13086 25540 13090 25596
rect 13026 25536 13090 25540
rect 13106 25596 13170 25600
rect 13106 25540 13110 25596
rect 13110 25540 13166 25596
rect 13166 25540 13170 25596
rect 13106 25536 13170 25540
rect 13186 25596 13250 25600
rect 13186 25540 13190 25596
rect 13190 25540 13246 25596
rect 13246 25540 13250 25596
rect 13186 25536 13250 25540
rect 4378 25052 4442 25056
rect 4378 24996 4382 25052
rect 4382 24996 4438 25052
rect 4438 24996 4442 25052
rect 4378 24992 4442 24996
rect 4458 25052 4522 25056
rect 4458 24996 4462 25052
rect 4462 24996 4518 25052
rect 4518 24996 4522 25052
rect 4458 24992 4522 24996
rect 4538 25052 4602 25056
rect 4538 24996 4542 25052
rect 4542 24996 4598 25052
rect 4598 24996 4602 25052
rect 4538 24992 4602 24996
rect 4618 25052 4682 25056
rect 4618 24996 4622 25052
rect 4622 24996 4678 25052
rect 4678 24996 4682 25052
rect 4618 24992 4682 24996
rect 7805 25052 7869 25056
rect 7805 24996 7809 25052
rect 7809 24996 7865 25052
rect 7865 24996 7869 25052
rect 7805 24992 7869 24996
rect 7885 25052 7949 25056
rect 7885 24996 7889 25052
rect 7889 24996 7945 25052
rect 7945 24996 7949 25052
rect 7885 24992 7949 24996
rect 7965 25052 8029 25056
rect 7965 24996 7969 25052
rect 7969 24996 8025 25052
rect 8025 24996 8029 25052
rect 7965 24992 8029 24996
rect 8045 25052 8109 25056
rect 8045 24996 8049 25052
rect 8049 24996 8105 25052
rect 8105 24996 8109 25052
rect 8045 24992 8109 24996
rect 11232 25052 11296 25056
rect 11232 24996 11236 25052
rect 11236 24996 11292 25052
rect 11292 24996 11296 25052
rect 11232 24992 11296 24996
rect 11312 25052 11376 25056
rect 11312 24996 11316 25052
rect 11316 24996 11372 25052
rect 11372 24996 11376 25052
rect 11312 24992 11376 24996
rect 11392 25052 11456 25056
rect 11392 24996 11396 25052
rect 11396 24996 11452 25052
rect 11452 24996 11456 25052
rect 11392 24992 11456 24996
rect 11472 25052 11536 25056
rect 11472 24996 11476 25052
rect 11476 24996 11532 25052
rect 11532 24996 11536 25052
rect 11472 24992 11536 24996
rect 14659 25052 14723 25056
rect 14659 24996 14663 25052
rect 14663 24996 14719 25052
rect 14719 24996 14723 25052
rect 14659 24992 14723 24996
rect 14739 25052 14803 25056
rect 14739 24996 14743 25052
rect 14743 24996 14799 25052
rect 14799 24996 14803 25052
rect 14739 24992 14803 24996
rect 14819 25052 14883 25056
rect 14819 24996 14823 25052
rect 14823 24996 14879 25052
rect 14879 24996 14883 25052
rect 14819 24992 14883 24996
rect 14899 25052 14963 25056
rect 14899 24996 14903 25052
rect 14903 24996 14959 25052
rect 14959 24996 14963 25052
rect 14899 24992 14963 24996
rect 2665 24508 2729 24512
rect 2665 24452 2669 24508
rect 2669 24452 2725 24508
rect 2725 24452 2729 24508
rect 2665 24448 2729 24452
rect 2745 24508 2809 24512
rect 2745 24452 2749 24508
rect 2749 24452 2805 24508
rect 2805 24452 2809 24508
rect 2745 24448 2809 24452
rect 2825 24508 2889 24512
rect 2825 24452 2829 24508
rect 2829 24452 2885 24508
rect 2885 24452 2889 24508
rect 2825 24448 2889 24452
rect 2905 24508 2969 24512
rect 2905 24452 2909 24508
rect 2909 24452 2965 24508
rect 2965 24452 2969 24508
rect 2905 24448 2969 24452
rect 6092 24508 6156 24512
rect 6092 24452 6096 24508
rect 6096 24452 6152 24508
rect 6152 24452 6156 24508
rect 6092 24448 6156 24452
rect 6172 24508 6236 24512
rect 6172 24452 6176 24508
rect 6176 24452 6232 24508
rect 6232 24452 6236 24508
rect 6172 24448 6236 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 9519 24508 9583 24512
rect 9519 24452 9523 24508
rect 9523 24452 9579 24508
rect 9579 24452 9583 24508
rect 9519 24448 9583 24452
rect 9599 24508 9663 24512
rect 9599 24452 9603 24508
rect 9603 24452 9659 24508
rect 9659 24452 9663 24508
rect 9599 24448 9663 24452
rect 9679 24508 9743 24512
rect 9679 24452 9683 24508
rect 9683 24452 9739 24508
rect 9739 24452 9743 24508
rect 9679 24448 9743 24452
rect 9759 24508 9823 24512
rect 9759 24452 9763 24508
rect 9763 24452 9819 24508
rect 9819 24452 9823 24508
rect 9759 24448 9823 24452
rect 12946 24508 13010 24512
rect 12946 24452 12950 24508
rect 12950 24452 13006 24508
rect 13006 24452 13010 24508
rect 12946 24448 13010 24452
rect 13026 24508 13090 24512
rect 13026 24452 13030 24508
rect 13030 24452 13086 24508
rect 13086 24452 13090 24508
rect 13026 24448 13090 24452
rect 13106 24508 13170 24512
rect 13106 24452 13110 24508
rect 13110 24452 13166 24508
rect 13166 24452 13170 24508
rect 13106 24448 13170 24452
rect 13186 24508 13250 24512
rect 13186 24452 13190 24508
rect 13190 24452 13246 24508
rect 13246 24452 13250 24508
rect 13186 24448 13250 24452
rect 4378 23964 4442 23968
rect 4378 23908 4382 23964
rect 4382 23908 4438 23964
rect 4438 23908 4442 23964
rect 4378 23904 4442 23908
rect 4458 23964 4522 23968
rect 4458 23908 4462 23964
rect 4462 23908 4518 23964
rect 4518 23908 4522 23964
rect 4458 23904 4522 23908
rect 4538 23964 4602 23968
rect 4538 23908 4542 23964
rect 4542 23908 4598 23964
rect 4598 23908 4602 23964
rect 4538 23904 4602 23908
rect 4618 23964 4682 23968
rect 4618 23908 4622 23964
rect 4622 23908 4678 23964
rect 4678 23908 4682 23964
rect 4618 23904 4682 23908
rect 7805 23964 7869 23968
rect 7805 23908 7809 23964
rect 7809 23908 7865 23964
rect 7865 23908 7869 23964
rect 7805 23904 7869 23908
rect 7885 23964 7949 23968
rect 7885 23908 7889 23964
rect 7889 23908 7945 23964
rect 7945 23908 7949 23964
rect 7885 23904 7949 23908
rect 7965 23964 8029 23968
rect 7965 23908 7969 23964
rect 7969 23908 8025 23964
rect 8025 23908 8029 23964
rect 7965 23904 8029 23908
rect 8045 23964 8109 23968
rect 8045 23908 8049 23964
rect 8049 23908 8105 23964
rect 8105 23908 8109 23964
rect 8045 23904 8109 23908
rect 11232 23964 11296 23968
rect 11232 23908 11236 23964
rect 11236 23908 11292 23964
rect 11292 23908 11296 23964
rect 11232 23904 11296 23908
rect 11312 23964 11376 23968
rect 11312 23908 11316 23964
rect 11316 23908 11372 23964
rect 11372 23908 11376 23964
rect 11312 23904 11376 23908
rect 11392 23964 11456 23968
rect 11392 23908 11396 23964
rect 11396 23908 11452 23964
rect 11452 23908 11456 23964
rect 11392 23904 11456 23908
rect 11472 23964 11536 23968
rect 11472 23908 11476 23964
rect 11476 23908 11532 23964
rect 11532 23908 11536 23964
rect 11472 23904 11536 23908
rect 14659 23964 14723 23968
rect 14659 23908 14663 23964
rect 14663 23908 14719 23964
rect 14719 23908 14723 23964
rect 14659 23904 14723 23908
rect 14739 23964 14803 23968
rect 14739 23908 14743 23964
rect 14743 23908 14799 23964
rect 14799 23908 14803 23964
rect 14739 23904 14803 23908
rect 14819 23964 14883 23968
rect 14819 23908 14823 23964
rect 14823 23908 14879 23964
rect 14879 23908 14883 23964
rect 14819 23904 14883 23908
rect 14899 23964 14963 23968
rect 14899 23908 14903 23964
rect 14903 23908 14959 23964
rect 14959 23908 14963 23964
rect 14899 23904 14963 23908
rect 2665 23420 2729 23424
rect 2665 23364 2669 23420
rect 2669 23364 2725 23420
rect 2725 23364 2729 23420
rect 2665 23360 2729 23364
rect 2745 23420 2809 23424
rect 2745 23364 2749 23420
rect 2749 23364 2805 23420
rect 2805 23364 2809 23420
rect 2745 23360 2809 23364
rect 2825 23420 2889 23424
rect 2825 23364 2829 23420
rect 2829 23364 2885 23420
rect 2885 23364 2889 23420
rect 2825 23360 2889 23364
rect 2905 23420 2969 23424
rect 2905 23364 2909 23420
rect 2909 23364 2965 23420
rect 2965 23364 2969 23420
rect 2905 23360 2969 23364
rect 6092 23420 6156 23424
rect 6092 23364 6096 23420
rect 6096 23364 6152 23420
rect 6152 23364 6156 23420
rect 6092 23360 6156 23364
rect 6172 23420 6236 23424
rect 6172 23364 6176 23420
rect 6176 23364 6232 23420
rect 6232 23364 6236 23420
rect 6172 23360 6236 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 9519 23420 9583 23424
rect 9519 23364 9523 23420
rect 9523 23364 9579 23420
rect 9579 23364 9583 23420
rect 9519 23360 9583 23364
rect 9599 23420 9663 23424
rect 9599 23364 9603 23420
rect 9603 23364 9659 23420
rect 9659 23364 9663 23420
rect 9599 23360 9663 23364
rect 9679 23420 9743 23424
rect 9679 23364 9683 23420
rect 9683 23364 9739 23420
rect 9739 23364 9743 23420
rect 9679 23360 9743 23364
rect 9759 23420 9823 23424
rect 9759 23364 9763 23420
rect 9763 23364 9819 23420
rect 9819 23364 9823 23420
rect 9759 23360 9823 23364
rect 12946 23420 13010 23424
rect 12946 23364 12950 23420
rect 12950 23364 13006 23420
rect 13006 23364 13010 23420
rect 12946 23360 13010 23364
rect 13026 23420 13090 23424
rect 13026 23364 13030 23420
rect 13030 23364 13086 23420
rect 13086 23364 13090 23420
rect 13026 23360 13090 23364
rect 13106 23420 13170 23424
rect 13106 23364 13110 23420
rect 13110 23364 13166 23420
rect 13166 23364 13170 23420
rect 13106 23360 13170 23364
rect 13186 23420 13250 23424
rect 13186 23364 13190 23420
rect 13190 23364 13246 23420
rect 13246 23364 13250 23420
rect 13186 23360 13250 23364
rect 4378 22876 4442 22880
rect 4378 22820 4382 22876
rect 4382 22820 4438 22876
rect 4438 22820 4442 22876
rect 4378 22816 4442 22820
rect 4458 22876 4522 22880
rect 4458 22820 4462 22876
rect 4462 22820 4518 22876
rect 4518 22820 4522 22876
rect 4458 22816 4522 22820
rect 4538 22876 4602 22880
rect 4538 22820 4542 22876
rect 4542 22820 4598 22876
rect 4598 22820 4602 22876
rect 4538 22816 4602 22820
rect 4618 22876 4682 22880
rect 4618 22820 4622 22876
rect 4622 22820 4678 22876
rect 4678 22820 4682 22876
rect 4618 22816 4682 22820
rect 7805 22876 7869 22880
rect 7805 22820 7809 22876
rect 7809 22820 7865 22876
rect 7865 22820 7869 22876
rect 7805 22816 7869 22820
rect 7885 22876 7949 22880
rect 7885 22820 7889 22876
rect 7889 22820 7945 22876
rect 7945 22820 7949 22876
rect 7885 22816 7949 22820
rect 7965 22876 8029 22880
rect 7965 22820 7969 22876
rect 7969 22820 8025 22876
rect 8025 22820 8029 22876
rect 7965 22816 8029 22820
rect 8045 22876 8109 22880
rect 8045 22820 8049 22876
rect 8049 22820 8105 22876
rect 8105 22820 8109 22876
rect 8045 22816 8109 22820
rect 11232 22876 11296 22880
rect 11232 22820 11236 22876
rect 11236 22820 11292 22876
rect 11292 22820 11296 22876
rect 11232 22816 11296 22820
rect 11312 22876 11376 22880
rect 11312 22820 11316 22876
rect 11316 22820 11372 22876
rect 11372 22820 11376 22876
rect 11312 22816 11376 22820
rect 11392 22876 11456 22880
rect 11392 22820 11396 22876
rect 11396 22820 11452 22876
rect 11452 22820 11456 22876
rect 11392 22816 11456 22820
rect 11472 22876 11536 22880
rect 11472 22820 11476 22876
rect 11476 22820 11532 22876
rect 11532 22820 11536 22876
rect 11472 22816 11536 22820
rect 14659 22876 14723 22880
rect 14659 22820 14663 22876
rect 14663 22820 14719 22876
rect 14719 22820 14723 22876
rect 14659 22816 14723 22820
rect 14739 22876 14803 22880
rect 14739 22820 14743 22876
rect 14743 22820 14799 22876
rect 14799 22820 14803 22876
rect 14739 22816 14803 22820
rect 14819 22876 14883 22880
rect 14819 22820 14823 22876
rect 14823 22820 14879 22876
rect 14879 22820 14883 22876
rect 14819 22816 14883 22820
rect 14899 22876 14963 22880
rect 14899 22820 14903 22876
rect 14903 22820 14959 22876
rect 14959 22820 14963 22876
rect 14899 22816 14963 22820
rect 2665 22332 2729 22336
rect 2665 22276 2669 22332
rect 2669 22276 2725 22332
rect 2725 22276 2729 22332
rect 2665 22272 2729 22276
rect 2745 22332 2809 22336
rect 2745 22276 2749 22332
rect 2749 22276 2805 22332
rect 2805 22276 2809 22332
rect 2745 22272 2809 22276
rect 2825 22332 2889 22336
rect 2825 22276 2829 22332
rect 2829 22276 2885 22332
rect 2885 22276 2889 22332
rect 2825 22272 2889 22276
rect 2905 22332 2969 22336
rect 2905 22276 2909 22332
rect 2909 22276 2965 22332
rect 2965 22276 2969 22332
rect 2905 22272 2969 22276
rect 6092 22332 6156 22336
rect 6092 22276 6096 22332
rect 6096 22276 6152 22332
rect 6152 22276 6156 22332
rect 6092 22272 6156 22276
rect 6172 22332 6236 22336
rect 6172 22276 6176 22332
rect 6176 22276 6232 22332
rect 6232 22276 6236 22332
rect 6172 22272 6236 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 9519 22332 9583 22336
rect 9519 22276 9523 22332
rect 9523 22276 9579 22332
rect 9579 22276 9583 22332
rect 9519 22272 9583 22276
rect 9599 22332 9663 22336
rect 9599 22276 9603 22332
rect 9603 22276 9659 22332
rect 9659 22276 9663 22332
rect 9599 22272 9663 22276
rect 9679 22332 9743 22336
rect 9679 22276 9683 22332
rect 9683 22276 9739 22332
rect 9739 22276 9743 22332
rect 9679 22272 9743 22276
rect 9759 22332 9823 22336
rect 9759 22276 9763 22332
rect 9763 22276 9819 22332
rect 9819 22276 9823 22332
rect 9759 22272 9823 22276
rect 12946 22332 13010 22336
rect 12946 22276 12950 22332
rect 12950 22276 13006 22332
rect 13006 22276 13010 22332
rect 12946 22272 13010 22276
rect 13026 22332 13090 22336
rect 13026 22276 13030 22332
rect 13030 22276 13086 22332
rect 13086 22276 13090 22332
rect 13026 22272 13090 22276
rect 13106 22332 13170 22336
rect 13106 22276 13110 22332
rect 13110 22276 13166 22332
rect 13166 22276 13170 22332
rect 13106 22272 13170 22276
rect 13186 22332 13250 22336
rect 13186 22276 13190 22332
rect 13190 22276 13246 22332
rect 13246 22276 13250 22332
rect 13186 22272 13250 22276
rect 4378 21788 4442 21792
rect 4378 21732 4382 21788
rect 4382 21732 4438 21788
rect 4438 21732 4442 21788
rect 4378 21728 4442 21732
rect 4458 21788 4522 21792
rect 4458 21732 4462 21788
rect 4462 21732 4518 21788
rect 4518 21732 4522 21788
rect 4458 21728 4522 21732
rect 4538 21788 4602 21792
rect 4538 21732 4542 21788
rect 4542 21732 4598 21788
rect 4598 21732 4602 21788
rect 4538 21728 4602 21732
rect 4618 21788 4682 21792
rect 4618 21732 4622 21788
rect 4622 21732 4678 21788
rect 4678 21732 4682 21788
rect 4618 21728 4682 21732
rect 7805 21788 7869 21792
rect 7805 21732 7809 21788
rect 7809 21732 7865 21788
rect 7865 21732 7869 21788
rect 7805 21728 7869 21732
rect 7885 21788 7949 21792
rect 7885 21732 7889 21788
rect 7889 21732 7945 21788
rect 7945 21732 7949 21788
rect 7885 21728 7949 21732
rect 7965 21788 8029 21792
rect 7965 21732 7969 21788
rect 7969 21732 8025 21788
rect 8025 21732 8029 21788
rect 7965 21728 8029 21732
rect 8045 21788 8109 21792
rect 8045 21732 8049 21788
rect 8049 21732 8105 21788
rect 8105 21732 8109 21788
rect 8045 21728 8109 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 11392 21788 11456 21792
rect 11392 21732 11396 21788
rect 11396 21732 11452 21788
rect 11452 21732 11456 21788
rect 11392 21728 11456 21732
rect 11472 21788 11536 21792
rect 11472 21732 11476 21788
rect 11476 21732 11532 21788
rect 11532 21732 11536 21788
rect 11472 21728 11536 21732
rect 14659 21788 14723 21792
rect 14659 21732 14663 21788
rect 14663 21732 14719 21788
rect 14719 21732 14723 21788
rect 14659 21728 14723 21732
rect 14739 21788 14803 21792
rect 14739 21732 14743 21788
rect 14743 21732 14799 21788
rect 14799 21732 14803 21788
rect 14739 21728 14803 21732
rect 14819 21788 14883 21792
rect 14819 21732 14823 21788
rect 14823 21732 14879 21788
rect 14879 21732 14883 21788
rect 14819 21728 14883 21732
rect 14899 21788 14963 21792
rect 14899 21732 14903 21788
rect 14903 21732 14959 21788
rect 14959 21732 14963 21788
rect 14899 21728 14963 21732
rect 2665 21244 2729 21248
rect 2665 21188 2669 21244
rect 2669 21188 2725 21244
rect 2725 21188 2729 21244
rect 2665 21184 2729 21188
rect 2745 21244 2809 21248
rect 2745 21188 2749 21244
rect 2749 21188 2805 21244
rect 2805 21188 2809 21244
rect 2745 21184 2809 21188
rect 2825 21244 2889 21248
rect 2825 21188 2829 21244
rect 2829 21188 2885 21244
rect 2885 21188 2889 21244
rect 2825 21184 2889 21188
rect 2905 21244 2969 21248
rect 2905 21188 2909 21244
rect 2909 21188 2965 21244
rect 2965 21188 2969 21244
rect 2905 21184 2969 21188
rect 6092 21244 6156 21248
rect 6092 21188 6096 21244
rect 6096 21188 6152 21244
rect 6152 21188 6156 21244
rect 6092 21184 6156 21188
rect 6172 21244 6236 21248
rect 6172 21188 6176 21244
rect 6176 21188 6232 21244
rect 6232 21188 6236 21244
rect 6172 21184 6236 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 9519 21244 9583 21248
rect 9519 21188 9523 21244
rect 9523 21188 9579 21244
rect 9579 21188 9583 21244
rect 9519 21184 9583 21188
rect 9599 21244 9663 21248
rect 9599 21188 9603 21244
rect 9603 21188 9659 21244
rect 9659 21188 9663 21244
rect 9599 21184 9663 21188
rect 9679 21244 9743 21248
rect 9679 21188 9683 21244
rect 9683 21188 9739 21244
rect 9739 21188 9743 21244
rect 9679 21184 9743 21188
rect 9759 21244 9823 21248
rect 9759 21188 9763 21244
rect 9763 21188 9819 21244
rect 9819 21188 9823 21244
rect 9759 21184 9823 21188
rect 12946 21244 13010 21248
rect 12946 21188 12950 21244
rect 12950 21188 13006 21244
rect 13006 21188 13010 21244
rect 12946 21184 13010 21188
rect 13026 21244 13090 21248
rect 13026 21188 13030 21244
rect 13030 21188 13086 21244
rect 13086 21188 13090 21244
rect 13026 21184 13090 21188
rect 13106 21244 13170 21248
rect 13106 21188 13110 21244
rect 13110 21188 13166 21244
rect 13166 21188 13170 21244
rect 13106 21184 13170 21188
rect 13186 21244 13250 21248
rect 13186 21188 13190 21244
rect 13190 21188 13246 21244
rect 13246 21188 13250 21244
rect 13186 21184 13250 21188
rect 4378 20700 4442 20704
rect 4378 20644 4382 20700
rect 4382 20644 4438 20700
rect 4438 20644 4442 20700
rect 4378 20640 4442 20644
rect 4458 20700 4522 20704
rect 4458 20644 4462 20700
rect 4462 20644 4518 20700
rect 4518 20644 4522 20700
rect 4458 20640 4522 20644
rect 4538 20700 4602 20704
rect 4538 20644 4542 20700
rect 4542 20644 4598 20700
rect 4598 20644 4602 20700
rect 4538 20640 4602 20644
rect 4618 20700 4682 20704
rect 4618 20644 4622 20700
rect 4622 20644 4678 20700
rect 4678 20644 4682 20700
rect 4618 20640 4682 20644
rect 7805 20700 7869 20704
rect 7805 20644 7809 20700
rect 7809 20644 7865 20700
rect 7865 20644 7869 20700
rect 7805 20640 7869 20644
rect 7885 20700 7949 20704
rect 7885 20644 7889 20700
rect 7889 20644 7945 20700
rect 7945 20644 7949 20700
rect 7885 20640 7949 20644
rect 7965 20700 8029 20704
rect 7965 20644 7969 20700
rect 7969 20644 8025 20700
rect 8025 20644 8029 20700
rect 7965 20640 8029 20644
rect 8045 20700 8109 20704
rect 8045 20644 8049 20700
rect 8049 20644 8105 20700
rect 8105 20644 8109 20700
rect 8045 20640 8109 20644
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 11392 20700 11456 20704
rect 11392 20644 11396 20700
rect 11396 20644 11452 20700
rect 11452 20644 11456 20700
rect 11392 20640 11456 20644
rect 11472 20700 11536 20704
rect 11472 20644 11476 20700
rect 11476 20644 11532 20700
rect 11532 20644 11536 20700
rect 11472 20640 11536 20644
rect 14659 20700 14723 20704
rect 14659 20644 14663 20700
rect 14663 20644 14719 20700
rect 14719 20644 14723 20700
rect 14659 20640 14723 20644
rect 14739 20700 14803 20704
rect 14739 20644 14743 20700
rect 14743 20644 14799 20700
rect 14799 20644 14803 20700
rect 14739 20640 14803 20644
rect 14819 20700 14883 20704
rect 14819 20644 14823 20700
rect 14823 20644 14879 20700
rect 14879 20644 14883 20700
rect 14819 20640 14883 20644
rect 14899 20700 14963 20704
rect 14899 20644 14903 20700
rect 14903 20644 14959 20700
rect 14959 20644 14963 20700
rect 14899 20640 14963 20644
rect 2665 20156 2729 20160
rect 2665 20100 2669 20156
rect 2669 20100 2725 20156
rect 2725 20100 2729 20156
rect 2665 20096 2729 20100
rect 2745 20156 2809 20160
rect 2745 20100 2749 20156
rect 2749 20100 2805 20156
rect 2805 20100 2809 20156
rect 2745 20096 2809 20100
rect 2825 20156 2889 20160
rect 2825 20100 2829 20156
rect 2829 20100 2885 20156
rect 2885 20100 2889 20156
rect 2825 20096 2889 20100
rect 2905 20156 2969 20160
rect 2905 20100 2909 20156
rect 2909 20100 2965 20156
rect 2965 20100 2969 20156
rect 2905 20096 2969 20100
rect 6092 20156 6156 20160
rect 6092 20100 6096 20156
rect 6096 20100 6152 20156
rect 6152 20100 6156 20156
rect 6092 20096 6156 20100
rect 6172 20156 6236 20160
rect 6172 20100 6176 20156
rect 6176 20100 6232 20156
rect 6232 20100 6236 20156
rect 6172 20096 6236 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 9519 20156 9583 20160
rect 9519 20100 9523 20156
rect 9523 20100 9579 20156
rect 9579 20100 9583 20156
rect 9519 20096 9583 20100
rect 9599 20156 9663 20160
rect 9599 20100 9603 20156
rect 9603 20100 9659 20156
rect 9659 20100 9663 20156
rect 9599 20096 9663 20100
rect 9679 20156 9743 20160
rect 9679 20100 9683 20156
rect 9683 20100 9739 20156
rect 9739 20100 9743 20156
rect 9679 20096 9743 20100
rect 9759 20156 9823 20160
rect 9759 20100 9763 20156
rect 9763 20100 9819 20156
rect 9819 20100 9823 20156
rect 9759 20096 9823 20100
rect 12946 20156 13010 20160
rect 12946 20100 12950 20156
rect 12950 20100 13006 20156
rect 13006 20100 13010 20156
rect 12946 20096 13010 20100
rect 13026 20156 13090 20160
rect 13026 20100 13030 20156
rect 13030 20100 13086 20156
rect 13086 20100 13090 20156
rect 13026 20096 13090 20100
rect 13106 20156 13170 20160
rect 13106 20100 13110 20156
rect 13110 20100 13166 20156
rect 13166 20100 13170 20156
rect 13106 20096 13170 20100
rect 13186 20156 13250 20160
rect 13186 20100 13190 20156
rect 13190 20100 13246 20156
rect 13246 20100 13250 20156
rect 13186 20096 13250 20100
rect 4378 19612 4442 19616
rect 4378 19556 4382 19612
rect 4382 19556 4438 19612
rect 4438 19556 4442 19612
rect 4378 19552 4442 19556
rect 4458 19612 4522 19616
rect 4458 19556 4462 19612
rect 4462 19556 4518 19612
rect 4518 19556 4522 19612
rect 4458 19552 4522 19556
rect 4538 19612 4602 19616
rect 4538 19556 4542 19612
rect 4542 19556 4598 19612
rect 4598 19556 4602 19612
rect 4538 19552 4602 19556
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 7805 19612 7869 19616
rect 7805 19556 7809 19612
rect 7809 19556 7865 19612
rect 7865 19556 7869 19612
rect 7805 19552 7869 19556
rect 7885 19612 7949 19616
rect 7885 19556 7889 19612
rect 7889 19556 7945 19612
rect 7945 19556 7949 19612
rect 7885 19552 7949 19556
rect 7965 19612 8029 19616
rect 7965 19556 7969 19612
rect 7969 19556 8025 19612
rect 8025 19556 8029 19612
rect 7965 19552 8029 19556
rect 8045 19612 8109 19616
rect 8045 19556 8049 19612
rect 8049 19556 8105 19612
rect 8105 19556 8109 19612
rect 8045 19552 8109 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 11392 19612 11456 19616
rect 11392 19556 11396 19612
rect 11396 19556 11452 19612
rect 11452 19556 11456 19612
rect 11392 19552 11456 19556
rect 11472 19612 11536 19616
rect 11472 19556 11476 19612
rect 11476 19556 11532 19612
rect 11532 19556 11536 19612
rect 11472 19552 11536 19556
rect 14659 19612 14723 19616
rect 14659 19556 14663 19612
rect 14663 19556 14719 19612
rect 14719 19556 14723 19612
rect 14659 19552 14723 19556
rect 14739 19612 14803 19616
rect 14739 19556 14743 19612
rect 14743 19556 14799 19612
rect 14799 19556 14803 19612
rect 14739 19552 14803 19556
rect 14819 19612 14883 19616
rect 14819 19556 14823 19612
rect 14823 19556 14879 19612
rect 14879 19556 14883 19612
rect 14819 19552 14883 19556
rect 14899 19612 14963 19616
rect 14899 19556 14903 19612
rect 14903 19556 14959 19612
rect 14959 19556 14963 19612
rect 14899 19552 14963 19556
rect 2665 19068 2729 19072
rect 2665 19012 2669 19068
rect 2669 19012 2725 19068
rect 2725 19012 2729 19068
rect 2665 19008 2729 19012
rect 2745 19068 2809 19072
rect 2745 19012 2749 19068
rect 2749 19012 2805 19068
rect 2805 19012 2809 19068
rect 2745 19008 2809 19012
rect 2825 19068 2889 19072
rect 2825 19012 2829 19068
rect 2829 19012 2885 19068
rect 2885 19012 2889 19068
rect 2825 19008 2889 19012
rect 2905 19068 2969 19072
rect 2905 19012 2909 19068
rect 2909 19012 2965 19068
rect 2965 19012 2969 19068
rect 2905 19008 2969 19012
rect 6092 19068 6156 19072
rect 6092 19012 6096 19068
rect 6096 19012 6152 19068
rect 6152 19012 6156 19068
rect 6092 19008 6156 19012
rect 6172 19068 6236 19072
rect 6172 19012 6176 19068
rect 6176 19012 6232 19068
rect 6232 19012 6236 19068
rect 6172 19008 6236 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 9519 19068 9583 19072
rect 9519 19012 9523 19068
rect 9523 19012 9579 19068
rect 9579 19012 9583 19068
rect 9519 19008 9583 19012
rect 9599 19068 9663 19072
rect 9599 19012 9603 19068
rect 9603 19012 9659 19068
rect 9659 19012 9663 19068
rect 9599 19008 9663 19012
rect 9679 19068 9743 19072
rect 9679 19012 9683 19068
rect 9683 19012 9739 19068
rect 9739 19012 9743 19068
rect 9679 19008 9743 19012
rect 9759 19068 9823 19072
rect 9759 19012 9763 19068
rect 9763 19012 9819 19068
rect 9819 19012 9823 19068
rect 9759 19008 9823 19012
rect 12946 19068 13010 19072
rect 12946 19012 12950 19068
rect 12950 19012 13006 19068
rect 13006 19012 13010 19068
rect 12946 19008 13010 19012
rect 13026 19068 13090 19072
rect 13026 19012 13030 19068
rect 13030 19012 13086 19068
rect 13086 19012 13090 19068
rect 13026 19008 13090 19012
rect 13106 19068 13170 19072
rect 13106 19012 13110 19068
rect 13110 19012 13166 19068
rect 13166 19012 13170 19068
rect 13106 19008 13170 19012
rect 13186 19068 13250 19072
rect 13186 19012 13190 19068
rect 13190 19012 13246 19068
rect 13246 19012 13250 19068
rect 13186 19008 13250 19012
rect 4378 18524 4442 18528
rect 4378 18468 4382 18524
rect 4382 18468 4438 18524
rect 4438 18468 4442 18524
rect 4378 18464 4442 18468
rect 4458 18524 4522 18528
rect 4458 18468 4462 18524
rect 4462 18468 4518 18524
rect 4518 18468 4522 18524
rect 4458 18464 4522 18468
rect 4538 18524 4602 18528
rect 4538 18468 4542 18524
rect 4542 18468 4598 18524
rect 4598 18468 4602 18524
rect 4538 18464 4602 18468
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 7805 18524 7869 18528
rect 7805 18468 7809 18524
rect 7809 18468 7865 18524
rect 7865 18468 7869 18524
rect 7805 18464 7869 18468
rect 7885 18524 7949 18528
rect 7885 18468 7889 18524
rect 7889 18468 7945 18524
rect 7945 18468 7949 18524
rect 7885 18464 7949 18468
rect 7965 18524 8029 18528
rect 7965 18468 7969 18524
rect 7969 18468 8025 18524
rect 8025 18468 8029 18524
rect 7965 18464 8029 18468
rect 8045 18524 8109 18528
rect 8045 18468 8049 18524
rect 8049 18468 8105 18524
rect 8105 18468 8109 18524
rect 8045 18464 8109 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 11392 18524 11456 18528
rect 11392 18468 11396 18524
rect 11396 18468 11452 18524
rect 11452 18468 11456 18524
rect 11392 18464 11456 18468
rect 11472 18524 11536 18528
rect 11472 18468 11476 18524
rect 11476 18468 11532 18524
rect 11532 18468 11536 18524
rect 11472 18464 11536 18468
rect 14659 18524 14723 18528
rect 14659 18468 14663 18524
rect 14663 18468 14719 18524
rect 14719 18468 14723 18524
rect 14659 18464 14723 18468
rect 14739 18524 14803 18528
rect 14739 18468 14743 18524
rect 14743 18468 14799 18524
rect 14799 18468 14803 18524
rect 14739 18464 14803 18468
rect 14819 18524 14883 18528
rect 14819 18468 14823 18524
rect 14823 18468 14879 18524
rect 14879 18468 14883 18524
rect 14819 18464 14883 18468
rect 14899 18524 14963 18528
rect 14899 18468 14903 18524
rect 14903 18468 14959 18524
rect 14959 18468 14963 18524
rect 14899 18464 14963 18468
rect 2665 17980 2729 17984
rect 2665 17924 2669 17980
rect 2669 17924 2725 17980
rect 2725 17924 2729 17980
rect 2665 17920 2729 17924
rect 2745 17980 2809 17984
rect 2745 17924 2749 17980
rect 2749 17924 2805 17980
rect 2805 17924 2809 17980
rect 2745 17920 2809 17924
rect 2825 17980 2889 17984
rect 2825 17924 2829 17980
rect 2829 17924 2885 17980
rect 2885 17924 2889 17980
rect 2825 17920 2889 17924
rect 2905 17980 2969 17984
rect 2905 17924 2909 17980
rect 2909 17924 2965 17980
rect 2965 17924 2969 17980
rect 2905 17920 2969 17924
rect 6092 17980 6156 17984
rect 6092 17924 6096 17980
rect 6096 17924 6152 17980
rect 6152 17924 6156 17980
rect 6092 17920 6156 17924
rect 6172 17980 6236 17984
rect 6172 17924 6176 17980
rect 6176 17924 6232 17980
rect 6232 17924 6236 17980
rect 6172 17920 6236 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 9519 17980 9583 17984
rect 9519 17924 9523 17980
rect 9523 17924 9579 17980
rect 9579 17924 9583 17980
rect 9519 17920 9583 17924
rect 9599 17980 9663 17984
rect 9599 17924 9603 17980
rect 9603 17924 9659 17980
rect 9659 17924 9663 17980
rect 9599 17920 9663 17924
rect 9679 17980 9743 17984
rect 9679 17924 9683 17980
rect 9683 17924 9739 17980
rect 9739 17924 9743 17980
rect 9679 17920 9743 17924
rect 9759 17980 9823 17984
rect 9759 17924 9763 17980
rect 9763 17924 9819 17980
rect 9819 17924 9823 17980
rect 9759 17920 9823 17924
rect 12946 17980 13010 17984
rect 12946 17924 12950 17980
rect 12950 17924 13006 17980
rect 13006 17924 13010 17980
rect 12946 17920 13010 17924
rect 13026 17980 13090 17984
rect 13026 17924 13030 17980
rect 13030 17924 13086 17980
rect 13086 17924 13090 17980
rect 13026 17920 13090 17924
rect 13106 17980 13170 17984
rect 13106 17924 13110 17980
rect 13110 17924 13166 17980
rect 13166 17924 13170 17980
rect 13106 17920 13170 17924
rect 13186 17980 13250 17984
rect 13186 17924 13190 17980
rect 13190 17924 13246 17980
rect 13246 17924 13250 17980
rect 13186 17920 13250 17924
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 7420 11052 7484 11116
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 7420 2484 7484 2548
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 27776 2977 27792
rect 2657 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2977 27776
rect 2657 26688 2977 27712
rect 2657 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2977 26688
rect 2657 25600 2977 26624
rect 2657 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2977 25600
rect 2657 24512 2977 25536
rect 2657 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2977 24512
rect 2657 23424 2977 24448
rect 2657 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2977 23424
rect 2657 22336 2977 23360
rect 2657 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2977 22336
rect 2657 21248 2977 22272
rect 2657 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2977 21248
rect 2657 20160 2977 21184
rect 2657 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2977 20160
rect 2657 19072 2977 20096
rect 2657 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2977 19072
rect 2657 17984 2977 19008
rect 2657 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2977 17984
rect 2657 16896 2977 17920
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 27232 4690 27792
rect 4370 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4690 27232
rect 4370 26144 4690 27168
rect 4370 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4690 26144
rect 4370 25056 4690 26080
rect 4370 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4690 25056
rect 4370 23968 4690 24992
rect 4370 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4690 23968
rect 4370 22880 4690 23904
rect 4370 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4690 22880
rect 4370 21792 4690 22816
rect 4370 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4690 21792
rect 4370 20704 4690 21728
rect 4370 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4690 20704
rect 4370 19616 4690 20640
rect 4370 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4690 19616
rect 4370 18528 4690 19552
rect 4370 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4690 18528
rect 4370 17440 4690 18464
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 27776 6404 27792
rect 6084 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6404 27776
rect 6084 26688 6404 27712
rect 6084 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6404 26688
rect 6084 25600 6404 26624
rect 6084 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6404 25600
rect 6084 24512 6404 25536
rect 6084 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6404 24512
rect 6084 23424 6404 24448
rect 6084 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6404 23424
rect 6084 22336 6404 23360
rect 6084 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6404 22336
rect 6084 21248 6404 22272
rect 6084 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6404 21248
rect 6084 20160 6404 21184
rect 6084 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6404 20160
rect 6084 19072 6404 20096
rect 6084 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6404 19072
rect 6084 17984 6404 19008
rect 6084 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6404 17984
rect 6084 16896 6404 17920
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 7797 27232 8117 27792
rect 7797 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8117 27232
rect 7797 26144 8117 27168
rect 7797 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8117 26144
rect 7797 25056 8117 26080
rect 7797 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8117 25056
rect 7797 23968 8117 24992
rect 7797 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8117 23968
rect 7797 22880 8117 23904
rect 7797 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8117 22880
rect 7797 21792 8117 22816
rect 7797 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8117 21792
rect 7797 20704 8117 21728
rect 7797 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8117 20704
rect 7797 19616 8117 20640
rect 7797 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8117 19616
rect 7797 18528 8117 19552
rect 7797 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8117 18528
rect 7797 17440 8117 18464
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7422 2549 7482 11051
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7419 2548 7485 2549
rect 7419 2484 7420 2548
rect 7484 2484 7485 2548
rect 7419 2483 7485 2484
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 27776 9831 27792
rect 9511 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9831 27776
rect 9511 26688 9831 27712
rect 9511 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9831 26688
rect 9511 25600 9831 26624
rect 9511 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9831 25600
rect 9511 24512 9831 25536
rect 9511 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9831 24512
rect 9511 23424 9831 24448
rect 9511 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9831 23424
rect 9511 22336 9831 23360
rect 9511 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9831 22336
rect 9511 21248 9831 22272
rect 9511 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9831 21248
rect 9511 20160 9831 21184
rect 9511 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9831 20160
rect 9511 19072 9831 20096
rect 9511 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9831 19072
rect 9511 17984 9831 19008
rect 9511 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9831 17984
rect 9511 16896 9831 17920
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 27232 11544 27792
rect 11224 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11544 27232
rect 11224 26144 11544 27168
rect 11224 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11544 26144
rect 11224 25056 11544 26080
rect 11224 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11544 25056
rect 11224 23968 11544 24992
rect 11224 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11544 23968
rect 11224 22880 11544 23904
rect 11224 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11544 22880
rect 11224 21792 11544 22816
rect 11224 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11544 21792
rect 11224 20704 11544 21728
rect 11224 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11544 20704
rect 11224 19616 11544 20640
rect 11224 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11544 19616
rect 11224 18528 11544 19552
rect 11224 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11544 18528
rect 11224 17440 11544 18464
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 27776 13258 27792
rect 12938 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13258 27776
rect 12938 26688 13258 27712
rect 12938 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13258 26688
rect 12938 25600 13258 26624
rect 12938 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13258 25600
rect 12938 24512 13258 25536
rect 12938 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13258 24512
rect 12938 23424 13258 24448
rect 12938 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13258 23424
rect 12938 22336 13258 23360
rect 12938 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13258 22336
rect 12938 21248 13258 22272
rect 12938 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13258 21248
rect 12938 20160 13258 21184
rect 12938 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13258 20160
rect 12938 19072 13258 20096
rect 12938 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13258 19072
rect 12938 17984 13258 19008
rect 12938 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13258 17984
rect 12938 16896 13258 17920
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 27232 14971 27792
rect 14651 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14971 27232
rect 14651 26144 14971 27168
rect 14651 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14971 26144
rect 14651 25056 14971 26080
rect 14651 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14971 25056
rect 14651 23968 14971 24992
rect 14651 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14971 23968
rect 14651 22880 14971 23904
rect 14651 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14971 22880
rect 14651 21792 14971 22816
rect 14651 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14971 21792
rect 14651 20704 14971 21728
rect 14651 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14971 20704
rect 14651 19616 14971 20640
rect 14651 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14971 19616
rect 14651 18528 14971 19552
rect 14651 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14971 18528
rect 14651 17440 14971 18464
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1670771148
transform -1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1670771148
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1670771148
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1670771148
transform -1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1670771148
transform -1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1670771148
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1670771148
transform -1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1670771148
transform -1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1670771148
transform -1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1670771148
transform -1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1670771148
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1670771148
transform -1 0 13064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1670771148
transform -1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1670771148
transform -1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output14_A
timestamp 1670771148
transform 1 0 10304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29
timestamp 1670771148
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1670771148
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1670771148
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1670771148
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1670771148
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62
timestamp 1670771148
transform 1 0 6808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68
timestamp 1670771148
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72
timestamp 1670771148
transform 1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1670771148
transform 1 0 8280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1670771148
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1670771148
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1670771148
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 9936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104
timestamp 1670771148
transform 1 0 10672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1670771148
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1670771148
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120
timestamp 1670771148
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128
timestamp 1670771148
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1670771148
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1670771148
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1670771148
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1670771148
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1670771148
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1670771148
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_14
timestamp 1670771148
transform 1 0 2392 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1670771148
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1670771148
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1670771148
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1670771148
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1670771148
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_72
timestamp 1670771148
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1670771148
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_84 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 8832 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_96
timestamp 1670771148
transform 1 0 9936 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_102
timestamp 1670771148
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1670771148
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1670771148
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1670771148
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_117
timestamp 1670771148
transform 1 0 11868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1670771148
transform 1 0 13064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1670771148
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1670771148
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1670771148
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1670771148
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1670771148
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1670771148
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1670771148
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1670771148
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1670771148
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1670771148
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1670771148
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1670771148
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1670771148
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1670771148
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp 1670771148
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1670771148
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1670771148
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1670771148
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1670771148
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1670771148
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1670771148
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_47
timestamp 1670771148
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1670771148
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1670771148
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1670771148
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_73
timestamp 1670771148
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_86
timestamp 1670771148
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_98
timestamp 1670771148
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1670771148
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1670771148
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1670771148
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1670771148
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1670771148
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1670771148
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1670771148
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1670771148
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1670771148
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1670771148
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1670771148
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1670771148
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp 1670771148
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1670771148
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1670771148
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1670771148
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_96
timestamp 1670771148
transform 1 0 9936 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_108
timestamp 1670771148
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_120
timestamp 1670771148
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1670771148
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1670771148
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1670771148
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1670771148
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1670771148
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1670771148
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1670771148
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1670771148
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1670771148
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1670771148
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1670771148
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_73
timestamp 1670771148
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_85
timestamp 1670771148
transform 1 0 8924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1670771148
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1670771148
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1670771148
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1670771148
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1670771148
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1670771148
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1670771148
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1670771148
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1670771148
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1670771148
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1670771148
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1670771148
transform 1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_50
timestamp 1670771148
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1670771148
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_71
timestamp 1670771148
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1670771148
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1670771148
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1670771148
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1670771148
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1670771148
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1670771148
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1670771148
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1670771148
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1670771148
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1670771148
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1670771148
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_23
timestamp 1670771148
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1670771148
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1670771148
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1670771148
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1670771148
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1670771148
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1670771148
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1670771148
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1670771148
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1670771148
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1670771148
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1670771148
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_137
timestamp 1670771148
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1670771148
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1670771148
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1670771148
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1670771148
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1670771148
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1670771148
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1670771148
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_64
timestamp 1670771148
transform 1 0 6992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1670771148
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1670771148
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1670771148
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1670771148
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1670771148
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1670771148
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1670771148
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1670771148
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1670771148
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1670771148
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_36
timestamp 1670771148
transform 1 0 4416 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_42
timestamp 1670771148
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1670771148
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1670771148
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1670771148
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1670771148
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1670771148
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1670771148
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1670771148
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1670771148
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1670771148
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1670771148
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp 1670771148
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_145
timestamp 1670771148
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1670771148
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1670771148
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1670771148
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1670771148
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1670771148
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1670771148
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1670771148
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1670771148
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1670771148
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1670771148
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_99
timestamp 1670771148
transform 1 0 10212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_111
timestamp 1670771148
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1670771148
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1670771148
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1670771148
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1670771148
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1670771148
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1670771148
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1670771148
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1670771148
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1670771148
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 1670771148
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1670771148
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1670771148
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1670771148
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp 1670771148
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_88
timestamp 1670771148
transform 1 0 9200 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_100
timestamp 1670771148
transform 1 0 10304 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1670771148
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1670771148
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1670771148
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1670771148
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1670771148
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1670771148
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1670771148
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1670771148
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_40
timestamp 1670771148
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_48
timestamp 1670771148
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_54
timestamp 1670771148
transform 1 0 6072 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1670771148
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1670771148
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1670771148
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1670771148
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1670771148
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1670771148
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1670771148
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1670771148
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1670771148
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1670771148
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1670771148
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1670771148
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1670771148
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1670771148
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1670771148
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1670771148
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1670771148
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_68
timestamp 1670771148
transform 1 0 7360 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_75
timestamp 1670771148
transform 1 0 8004 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_87
timestamp 1670771148
transform 1 0 9108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_99
timestamp 1670771148
transform 1 0 10212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1670771148
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1670771148
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1670771148
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1670771148
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_145
timestamp 1670771148
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1670771148
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1670771148
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1670771148
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1670771148
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1670771148
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1670771148
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1670771148
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1670771148
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1670771148
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_92
timestamp 1670771148
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_104
timestamp 1670771148
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_116
timestamp 1670771148
transform 1 0 11776 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_128
timestamp 1670771148
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1670771148
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1670771148
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1670771148
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1670771148
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_27
timestamp 1670771148
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1670771148
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1670771148
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1670771148
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1670771148
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1670771148
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_84
timestamp 1670771148
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_96
timestamp 1670771148
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1670771148
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1670771148
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1670771148
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1670771148
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_145
timestamp 1670771148
transform 1 0 14444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1670771148
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1670771148
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1670771148
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1670771148
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1670771148
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1670771148
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1670771148
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1670771148
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1670771148
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1670771148
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1670771148
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1670771148
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1670771148
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1670771148
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1670771148
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1670771148
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1670771148
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1670771148
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1670771148
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1670771148
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_35
timestamp 1670771148
transform 1 0 4324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1670771148
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1670771148
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1670771148
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1670771148
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1670771148
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1670771148
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1670771148
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1670771148
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1670771148
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1670771148
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1670771148
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1670771148
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1670771148
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1670771148
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1670771148
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1670771148
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1670771148
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_39
timestamp 1670771148
transform 1 0 4692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_67
timestamp 1670771148
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1670771148
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1670771148
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1670771148
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1670771148
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1670771148
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1670771148
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1670771148
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1670771148
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1670771148
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1670771148
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1670771148
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1670771148
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1670771148
transform 1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_44
timestamp 1670771148
transform 1 0 5152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1670771148
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1670771148
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1670771148
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 1670771148
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1670771148
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1670771148
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_99
timestamp 1670771148
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1670771148
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1670771148
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1670771148
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1670771148
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1670771148
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1670771148
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1670771148
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1670771148
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1670771148
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_37
timestamp 1670771148
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1670771148
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1670771148
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_68
timestamp 1670771148
transform 1 0 7360 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1670771148
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1670771148
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_90
timestamp 1670771148
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_102
timestamp 1670771148
transform 1 0 10488 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_114
timestamp 1670771148
transform 1 0 11592 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_126
timestamp 1670771148
transform 1 0 12696 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1670771148
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1670771148
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1670771148
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1670771148
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1670771148
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp 1670771148
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1670771148
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_50
timestamp 1670771148
transform 1 0 5704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1670771148
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1670771148
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_63
timestamp 1670771148
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_80
timestamp 1670771148
transform 1 0 8464 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_87
timestamp 1670771148
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1670771148
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1670771148
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1670771148
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1670771148
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_137
timestamp 1670771148
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_145
timestamp 1670771148
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1670771148
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1670771148
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1670771148
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1670771148
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1670771148
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1670771148
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1670771148
transform 1 0 5428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1670771148
transform 1 0 6992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1670771148
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1670771148
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1670771148
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_90
timestamp 1670771148
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_102
timestamp 1670771148
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_114
timestamp 1670771148
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_126
timestamp 1670771148
transform 1 0 12696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1670771148
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1670771148
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1670771148
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1670771148
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1670771148
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1670771148
transform 1 0 3588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1670771148
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1670771148
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1670771148
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1670771148
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1670771148
transform 1 0 8648 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_89
timestamp 1670771148
transform 1 0 9292 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1670771148
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1670771148
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1670771148
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1670771148
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1670771148
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_145
timestamp 1670771148
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1670771148
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1670771148
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1670771148
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1670771148
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1670771148
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1670771148
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1670771148
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1670771148
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1670771148
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1670771148
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1670771148
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1670771148
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1670771148
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1670771148
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1670771148
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1670771148
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1670771148
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1670771148
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_36
timestamp 1670771148
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1670771148
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1670771148
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1670771148
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1670771148
transform 1 0 7084 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1670771148
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1670771148
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1670771148
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1670771148
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1670771148
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1670771148
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1670771148
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1670771148
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1670771148
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1670771148
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1670771148
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1670771148
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_36
timestamp 1670771148
transform 1 0 4416 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1670771148
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1670771148
transform 1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1670771148
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1670771148
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1670771148
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_90
timestamp 1670771148
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_102
timestamp 1670771148
transform 1 0 10488 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_114
timestamp 1670771148
transform 1 0 11592 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_126
timestamp 1670771148
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1670771148
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1670771148
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1670771148
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1670771148
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1670771148
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1670771148
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_44
timestamp 1670771148
transform 1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1670771148
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1670771148
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1670771148
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_87
timestamp 1670771148
transform 1 0 9108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_99
timestamp 1670771148
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1670771148
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1670771148
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1670771148
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1670771148
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1670771148
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1670771148
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1670771148
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1670771148
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1670771148
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_41
timestamp 1670771148
transform 1 0 4876 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_47
timestamp 1670771148
transform 1 0 5428 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_55
timestamp 1670771148
transform 1 0 6164 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_63
timestamp 1670771148
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1670771148
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1670771148
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1670771148
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1670771148
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1670771148
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1670771148
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1670771148
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1670771148
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1670771148
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1670771148
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1670771148
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1670771148
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1670771148
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1670771148
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1670771148
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1670771148
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_65
timestamp 1670771148
transform 1 0 7084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_77
timestamp 1670771148
transform 1 0 8188 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_89
timestamp 1670771148
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1670771148
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1670771148
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1670771148
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1670771148
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_137
timestamp 1670771148
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_145
timestamp 1670771148
transform 1 0 14444 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1670771148
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1670771148
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1670771148
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1670771148
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1670771148
transform 1 0 4876 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_63
timestamp 1670771148
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_75
timestamp 1670771148
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1670771148
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1670771148
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1670771148
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1670771148
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1670771148
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1670771148
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1670771148
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1670771148
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1670771148
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1670771148
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1670771148
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1670771148
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_35
timestamp 1670771148
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1670771148
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1670771148
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_65
timestamp 1670771148
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_84
timestamp 1670771148
transform 1 0 8832 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_96
timestamp 1670771148
transform 1 0 9936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1670771148
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1670771148
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1670771148
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1670771148
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp 1670771148
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1670771148
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1670771148
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1670771148
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1670771148
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1670771148
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1670771148
transform 1 0 4968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp 1670771148
transform 1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1670771148
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1670771148
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1670771148
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1670771148
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1670771148
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1670771148
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1670771148
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1670771148
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1670771148
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1670771148
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_15
timestamp 1670771148
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1670771148
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1670771148
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1670771148
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_64
timestamp 1670771148
transform 1 0 6992 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_84
timestamp 1670771148
transform 1 0 8832 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_96
timestamp 1670771148
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1670771148
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1670771148
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1670771148
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_137
timestamp 1670771148
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_145
timestamp 1670771148
transform 1 0 14444 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1670771148
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_15
timestamp 1670771148
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1670771148
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1670771148
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1670771148
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_45
timestamp 1670771148
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_62
timestamp 1670771148
transform 1 0 6808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1670771148
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1670771148
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1670771148
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1670771148
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1670771148
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1670771148
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1670771148
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1670771148
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1670771148
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1670771148
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1670771148
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1670771148
transform 1 0 3588 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_31
timestamp 1670771148
transform 1 0 3956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1670771148
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1670771148
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1670771148
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1670771148
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1670771148
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1670771148
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1670771148
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1670771148
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1670771148
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1670771148
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_145
timestamp 1670771148
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1670771148
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1670771148
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1670771148
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1670771148
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_47
timestamp 1670771148
transform 1 0 5428 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_59
timestamp 1670771148
transform 1 0 6532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_71
timestamp 1670771148
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1670771148
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1670771148
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1670771148
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1670771148
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1670771148
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1670771148
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1670771148
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1670771148
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1670771148
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1670771148
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1670771148
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1670771148
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1670771148
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1670771148
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1670771148
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1670771148
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1670771148
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1670771148
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1670771148
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1670771148
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1670771148
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1670771148
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1670771148
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_137
timestamp 1670771148
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1670771148
transform 1 0 14444 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1670771148
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1670771148
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1670771148
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1670771148
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1670771148
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1670771148
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1670771148
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1670771148
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1670771148
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1670771148
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1670771148
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1670771148
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1670771148
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1670771148
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1670771148
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1670771148
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1670771148
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1670771148
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1670771148
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1670771148
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1670771148
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1670771148
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1670771148
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1670771148
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1670771148
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1670771148
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1670771148
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1670771148
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1670771148
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1670771148
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1670771148
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_137
timestamp 1670771148
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_144
timestamp 1670771148
transform 1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1670771148
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1670771148
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_12
timestamp 1670771148
transform 1 0 2208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1670771148
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1670771148
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1670771148
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1670771148
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1670771148
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1670771148
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1670771148
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1670771148
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1670771148
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1670771148
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1670771148
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_133
timestamp 1670771148
transform 1 0 13340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1670771148
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1670771148
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1670771148
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1670771148
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_10
timestamp 1670771148
transform 1 0 2024 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_18
timestamp 1670771148
transform 1 0 2760 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_30
timestamp 1670771148
transform 1 0 3864 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_42
timestamp 1670771148
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1670771148
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1670771148
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1670771148
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1670771148
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1670771148
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1670771148
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1670771148
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1670771148
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_121
timestamp 1670771148
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1670771148
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1670771148
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_142
timestamp 1670771148
transform 1 0 14168 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_3
timestamp 1670771148
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_11
timestamp 1670771148
transform 1 0 2116 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_16
timestamp 1670771148
transform 1 0 2576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1670771148
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_29
timestamp 1670771148
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_36
timestamp 1670771148
transform 1 0 4416 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1670771148
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_60
timestamp 1670771148
transform 1 0 6624 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_72
timestamp 1670771148
transform 1 0 7728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1670771148
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1670771148
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1670771148
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1670771148
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_129
timestamp 1670771148
transform 1 0 12972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1670771148
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1670771148
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1670771148
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1670771148
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_9
timestamp 1670771148
transform 1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_17
timestamp 1670771148
transform 1 0 2668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_25
timestamp 1670771148
transform 1 0 3404 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_33
timestamp 1670771148
transform 1 0 4140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_38
timestamp 1670771148
transform 1 0 4600 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_48
timestamp 1670771148
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1670771148
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_65
timestamp 1670771148
transform 1 0 7084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_77
timestamp 1670771148
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_82
timestamp 1670771148
transform 1 0 8648 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_94
timestamp 1670771148
transform 1 0 9752 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_102
timestamp 1670771148
transform 1 0 10488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1670771148
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1670771148
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1670771148
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_124
timestamp 1670771148
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1670771148
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_140
timestamp 1670771148
transform 1 0 13984 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1670771148
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_10
timestamp 1670771148
transform 1 0 2024 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_18
timestamp 1670771148
transform 1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1670771148
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_29
timestamp 1670771148
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_37
timestamp 1670771148
transform 1 0 4508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_42
timestamp 1670771148
transform 1 0 4968 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_50
timestamp 1670771148
transform 1 0 5704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1670771148
transform 1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_66
timestamp 1670771148
transform 1 0 7176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1670771148
transform 1 0 7912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1670771148
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1670771148
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1670771148
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_94
timestamp 1670771148
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1670771148
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_110
timestamp 1670771148
transform 1 0 11224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_118
timestamp 1670771148
transform 1 0 11960 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1670771148
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1670771148
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1670771148
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1670771148
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1670771148
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_9
timestamp 1670771148
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_14
timestamp 1670771148
transform 1 0 2392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_22
timestamp 1670771148
transform 1 0 3128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_30
timestamp 1670771148
transform 1 0 3864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_38
timestamp 1670771148
transform 1 0 4600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_46
timestamp 1670771148
transform 1 0 5336 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1670771148
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1670771148
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1670771148
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_68
timestamp 1670771148
transform 1 0 7360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp 1670771148
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_84
timestamp 1670771148
transform 1 0 8832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1670771148
transform 1 0 9936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1670771148
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1670771148
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_119
timestamp 1670771148
transform 1 0 12052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_127
timestamp 1670771148
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp 1670771148
transform 1 0 13524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1670771148
transform 1 0 14260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1670771148
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_10
timestamp 1670771148
transform 1 0 2024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_18
timestamp 1670771148
transform 1 0 2760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1670771148
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1670771148
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_33
timestamp 1670771148
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_38
timestamp 1670771148
transform 1 0 4600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_46
timestamp 1670771148
transform 1 0 5336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_54
timestamp 1670771148
transform 1 0 6072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_57
timestamp 1670771148
transform 1 0 6348 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_61
timestamp 1670771148
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_66
timestamp 1670771148
transform 1 0 7176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_74
timestamp 1670771148
transform 1 0 7912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1670771148
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1670771148
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_91
timestamp 1670771148
transform 1 0 9476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1670771148
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_107
timestamp 1670771148
transform 1 0 10948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_111
timestamp 1670771148
transform 1 0 11316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1670771148
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_119
timestamp 1670771148
transform 1 0 12052 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1670771148
transform 1 0 12788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1670771148
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1670771148
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1670771148
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1670771148
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1670771148
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1670771148
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1670771148
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1670771148
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1670771148
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1670771148
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1670771148
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1670771148
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1670771148
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1670771148
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1670771148
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1670771148
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1670771148
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1670771148
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1670771148
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1670771148
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1670771148
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1670771148
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1670771148
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1670771148
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1670771148
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1670771148
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1670771148
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1670771148
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1670771148
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1670771148
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1670771148
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1670771148
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1670771148
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1670771148
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1670771148
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1670771148
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1670771148
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1670771148
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1670771148
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1670771148
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1670771148
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1670771148
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1670771148
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1670771148
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1670771148
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1670771148
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1670771148
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1670771148
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1670771148
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1670771148
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1670771148
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1670771148
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1670771148
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1670771148
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1670771148
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1670771148
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1670771148
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1670771148
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1670771148
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1670771148
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1670771148
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1670771148
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1670771148
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1670771148
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1670771148
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1670771148
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1670771148
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1670771148
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1670771148
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1670771148
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1670771148
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1670771148
transform -1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1670771148
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1670771148
transform -1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1670771148
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1670771148
transform -1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1670771148
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1670771148
transform -1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1670771148
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1670771148
transform -1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1670771148
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1670771148
transform -1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1670771148
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1670771148
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1670771148
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1670771148
transform -1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1670771148
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1670771148
transform -1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1670771148
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1670771148
transform -1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1670771148
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1670771148
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1670771148
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1670771148
transform -1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1670771148
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1670771148
transform -1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1670771148
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1670771148
transform -1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1670771148
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1670771148
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1670771148
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1670771148
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1670771148
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1670771148
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1670771148
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1670771148
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1670771148
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1670771148
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1670771148
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1670771148
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1670771148
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1670771148
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1670771148
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1670771148
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1670771148
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1670771148
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1670771148
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1670771148
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1670771148
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1670771148
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1670771148
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1670771148
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1670771148
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1670771148
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1670771148
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1670771148
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1670771148
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1670771148
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1670771148
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1670771148
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1670771148
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1670771148
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1670771148
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1670771148
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1670771148
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1670771148
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1670771148
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1670771148
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1670771148
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1670771148
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1670771148
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1670771148
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1670771148
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1670771148
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1670771148
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1670771148
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1670771148
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1670771148
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1670771148
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1670771148
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1670771148
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1670771148
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1670771148
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1670771148
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1670771148
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1670771148
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1670771148
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1670771148
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1670771148
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1670771148
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1670771148
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1670771148
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1670771148
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1670771148
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1670771148
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1670771148
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1670771148
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1670771148
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1670771148
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1670771148
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1670771148
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1670771148
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1670771148
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1670771148
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1670771148
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1670771148
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1670771148
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1670771148
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1670771148
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1670771148
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1670771148
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1670771148
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1670771148
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1670771148
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1670771148
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1670771148
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1670771148
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1670771148
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1670771148
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1670771148
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1670771148
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1670771148
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1670771148
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1670771148
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1670771148
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1670771148
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1670771148
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1670771148
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1670771148
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1670771148
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1670771148
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1670771148
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1670771148
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1670771148
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1670771148
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1670771148
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1670771148
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1670771148
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1670771148
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1670771148
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1670771148
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1670771148
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1670771148
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1670771148
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1670771148
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1670771148
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1670771148
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1670771148
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1670771148
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _093_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _094_
timestamp 1670771148
transform 1 0 10120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _095_
timestamp 1670771148
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _096_
timestamp 1670771148
transform 1 0 8280 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _097_
timestamp 1670771148
transform 1 0 8280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _098_
timestamp 1670771148
transform 1 0 7544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _099_
timestamp 1670771148
transform 1 0 6808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _100_
timestamp 1670771148
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _101_
timestamp 1670771148
transform -1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _102_
timestamp 1670771148
transform 1 0 5336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _103_
timestamp 1670771148
transform -1 0 5520 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _104_
timestamp 1670771148
transform 1 0 4600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _105_
timestamp 1670771148
transform 1 0 4232 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _106_
timestamp 1670771148
transform 1 0 3128 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _107_
timestamp 1670771148
transform 1 0 3036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _108_
timestamp 1670771148
transform -1 0 2024 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _109_
timestamp 1670771148
transform 1 0 1564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _110_
timestamp 1670771148
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _111_
timestamp 1670771148
transform 1 0 13064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _112_
timestamp 1670771148
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _113_
timestamp 1670771148
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _114_
timestamp 1670771148
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _115_
timestamp 1670771148
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 6532 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1670771148
transform -1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1670771148
transform 1 0 9108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _120_
timestamp 1670771148
transform -1 0 8648 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _121_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _122_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1670771148
transform 1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _124_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _125_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _126_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1670771148
transform 1 0 6256 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _128_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _129_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 6900 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1670771148
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _131_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 8648 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1670771148
transform -1 0 7636 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _133_
timestamp 1670771148
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _134_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 7268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1670771148
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _136_
timestamp 1670771148
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _137_
timestamp 1670771148
transform 1 0 5336 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _138_
timestamp 1670771148
transform 1 0 5612 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _139_
timestamp 1670771148
transform -1 0 6808 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _140_
timestamp 1670771148
transform 1 0 6532 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1670771148
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _142_
timestamp 1670771148
transform -1 0 6072 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _143_
timestamp 1670771148
transform 1 0 6532 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _144_
timestamp 1670771148
transform 1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _145_
timestamp 1670771148
transform 1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1670771148
transform -1 0 6532 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _147_
timestamp 1670771148
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _148_
timestamp 1670771148
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _149_
timestamp 1670771148
transform 1 0 5060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _150_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _151_
timestamp 1670771148
transform 1 0 4232 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1670771148
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1670771148
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _154_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 4416 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _155_
timestamp 1670771148
transform -1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _156_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 9568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1670771148
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1670771148
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _159_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1670771148
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _161_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform -1 0 9384 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _162_
timestamp 1670771148
transform 1 0 8924 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1670771148
transform 1 0 9016 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 1670771148
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1670771148
transform 1 0 8096 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1670771148
transform 1 0 8280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1670771148
transform 1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _168_
timestamp 1670771148
transform 1 0 8096 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1670771148
transform 1 0 8372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 1670771148
transform 1 0 9108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _171_
timestamp 1670771148
transform 1 0 8004 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1670771148
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1670771148
transform -1 0 9016 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _174_
timestamp 1670771148
transform -1 0 10212 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1670771148
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _176_
timestamp 1670771148
transform -1 0 7728 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _177_
timestamp 1670771148
transform 1 0 7728 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1670771148
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1670771148
transform -1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _180_
timestamp 1670771148
transform 1 0 4692 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _181_
timestamp 1670771148
transform 1 0 7452 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 1670771148
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1670771148
transform 1 0 6532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _184_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 6900 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1670771148
transform 1 0 7544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 1670771148
transform 1 0 4232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1670771148
transform 1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _188_
timestamp 1670771148
transform 1 0 4324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _189_
timestamp 1670771148
transform -1 0 6532 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 1670771148
transform 1 0 4324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _191_
timestamp 1670771148
transform -1 0 5980 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 1670771148
transform -1 0 5244 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _193_
timestamp 1670771148
transform 1 0 4324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _194_
timestamp 1670771148
transform -1 0 6992 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1670771148
transform -1 0 3496 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 1670771148
transform -1 0 5980 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1670771148
transform -1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 1670771148
transform -1 0 5060 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1670771148
transform -1 0 4232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _200_
timestamp 1670771148
transform -1 0 5888 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _201_
timestamp 1670771148
transform -1 0 6072 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1670771148
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _203_
timestamp 1670771148
transform 1 0 4416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _204_
timestamp 1670771148
transform -1 0 7084 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1670771148
transform 1 0 7360 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _206_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 5520 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _207_
timestamp 1670771148
transform -1 0 5428 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _208_
timestamp 1670771148
transform 1 0 7452 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _209_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 7176 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1670771148
transform 1 0 6716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _211_
timestamp 1670771148
transform 1 0 6992 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1670771148
transform 1 0 6900 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1670771148
transform 1 0 7084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1670771148
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1670771148
transform -1 0 6716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1670771148
transform 1 0 5520 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1670771148
transform 1 0 4324 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1670771148
transform 1 0 3956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1670771148
transform 1 0 3956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1670771148
transform 1 0 7176 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1670771148
transform 1 0 7360 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1670771148
transform 1 0 7360 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1670771148
transform 1 0 7268 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1670771148
transform 1 0 7176 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1670771148
transform 1 0 7176 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1670771148
transform 1 0 6992 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1670771148
transform 1 0 4048 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1670771148
transform -1 0 3496 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1670771148
transform -1 0 5244 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1670771148
transform -1 0 4232 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1670771148
transform -1 0 5428 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1670771148
transform -1 0 5152 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1670771148
transform -1 0 5336 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1670771148
transform 1 0 5336 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1670771148
transform 1 0 6532 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1670771148
transform 1 0 6532 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1670771148
transform 1 0 5336 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1670771148
transform 1 0 4600 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1670771148
transform 1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1670771148
transform 1 0 5520 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1670771148
transform -1 0 6072 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 5428 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1670771148
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1670771148
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1670771148
transform 1 0 5244 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1670771148
transform 1 0 5244 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1670771148
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1670771148
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1670771148
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1670771148
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1670771148
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1670771148
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1670771148
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1670771148
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1670771148
transform -1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1670771148
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1670771148
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1670771148
transform 1 0 1932 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1670771148
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output14 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670771148
transform 1 0 10856 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1670771148
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1670771148
transform 1 0 11868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1670771148
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1670771148
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1670771148
transform 1 0 13892 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1670771148
transform 1 0 13156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1670771148
transform 1 0 11684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1670771148
transform -1 0 13800 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1670771148
transform 1 0 13340 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1670771148
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1670771148
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1670771148
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1670771148
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1670771148
transform 1 0 11684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1670771148
transform 1 0 2392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1670771148
transform -1 0 2024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1670771148
transform -1 0 2392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1670771148
transform -1 0 2668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1670771148
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1670771148
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1670771148
transform 1 0 10580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1670771148
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1670771148
transform 1 0 8280 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1670771148
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1670771148
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1670771148
transform -1 0 6072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1670771148
transform -1 0 6072 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1670771148
transform -1 0 4600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1670771148
transform -1 0 3496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1670771148
transform 1 0 10304 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1670771148
transform -1 0 3128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1670771148
transform -1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1670771148
transform -1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1670771148
transform -1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1670771148
transform 1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1670771148
transform 1 0 1840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1670771148
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1670771148
transform 1 0 9108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1670771148
transform 1 0 8464 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1670771148
transform 1 0 7728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1670771148
transform 1 0 6992 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1670771148
transform -1 0 5336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1670771148
transform -1 0 5336 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1670771148
transform -1 0 4600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1670771148
transform -1 0 3864 0 -1 27200
box -38 -48 406 592
<< labels >>
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 dac_in[0]
port 1 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 dac_in[1]
port 2 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 dac_in[2]
port 3 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 dac_in[3]
port 4 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 dac_in[4]
port 5 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 dac_in[5]
port 6 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 dac_in[6]
port 7 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 dac_in[7]
port 8 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 dac_in[8]
port 9 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 dac_in[9]
port 10 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 dummy
port 11 nsew signal input
flabel metal2 s 14186 29200 14242 30000 0 FreeSans 224 90 0 0 llsb
port 12 nsew signal tristate
flabel metal2 s 13910 29200 13966 30000 0 FreeSans 224 90 0 0 llsb_n
port 13 nsew signal tristate
flabel metal2 s 13634 29200 13690 30000 0 FreeSans 224 90 0 0 lsb[0]
port 14 nsew signal tristate
flabel metal2 s 13082 29200 13138 30000 0 FreeSans 224 90 0 0 lsb[1]
port 15 nsew signal tristate
flabel metal2 s 12530 29200 12586 30000 0 FreeSans 224 90 0 0 lsb[2]
port 16 nsew signal tristate
flabel metal2 s 11978 29200 12034 30000 0 FreeSans 224 90 0 0 lsb[3]
port 17 nsew signal tristate
flabel metal2 s 11426 29200 11482 30000 0 FreeSans 224 90 0 0 lsb[4]
port 18 nsew signal tristate
flabel metal2 s 10874 29200 10930 30000 0 FreeSans 224 90 0 0 lsb[5]
port 19 nsew signal tristate
flabel metal2 s 13358 29200 13414 30000 0 FreeSans 224 90 0 0 lsb_n[0]
port 20 nsew signal tristate
flabel metal2 s 12806 29200 12862 30000 0 FreeSans 224 90 0 0 lsb_n[1]
port 21 nsew signal tristate
flabel metal2 s 12254 29200 12310 30000 0 FreeSans 224 90 0 0 lsb_n[2]
port 22 nsew signal tristate
flabel metal2 s 11702 29200 11758 30000 0 FreeSans 224 90 0 0 lsb_n[3]
port 23 nsew signal tristate
flabel metal2 s 11150 29200 11206 30000 0 FreeSans 224 90 0 0 lsb_n[4]
port 24 nsew signal tristate
flabel metal2 s 10598 29200 10654 30000 0 FreeSans 224 90 0 0 lsb_n[5]
port 25 nsew signal tristate
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 msb[0]
port 26 nsew signal tristate
flabel metal2 s 4802 29200 4858 30000 0 FreeSans 224 90 0 0 msb[10]
port 27 nsew signal tristate
flabel metal2 s 4250 29200 4306 30000 0 FreeSans 224 90 0 0 msb[11]
port 28 nsew signal tristate
flabel metal2 s 3698 29200 3754 30000 0 FreeSans 224 90 0 0 msb[12]
port 29 nsew signal tristate
flabel metal2 s 3146 29200 3202 30000 0 FreeSans 224 90 0 0 msb[13]
port 30 nsew signal tristate
flabel metal2 s 2594 29200 2650 30000 0 FreeSans 224 90 0 0 msb[14]
port 31 nsew signal tristate
flabel metal2 s 2042 29200 2098 30000 0 FreeSans 224 90 0 0 msb[15]
port 32 nsew signal tristate
flabel metal2 s 9770 29200 9826 30000 0 FreeSans 224 90 0 0 msb[1]
port 33 nsew signal tristate
flabel metal2 s 9218 29200 9274 30000 0 FreeSans 224 90 0 0 msb[2]
port 34 nsew signal tristate
flabel metal2 s 8666 29200 8722 30000 0 FreeSans 224 90 0 0 msb[3]
port 35 nsew signal tristate
flabel metal2 s 8114 29200 8170 30000 0 FreeSans 224 90 0 0 msb[4]
port 36 nsew signal tristate
flabel metal2 s 7562 29200 7618 30000 0 FreeSans 224 90 0 0 msb[5]
port 37 nsew signal tristate
flabel metal2 s 7010 29200 7066 30000 0 FreeSans 224 90 0 0 msb[6]
port 38 nsew signal tristate
flabel metal2 s 6458 29200 6514 30000 0 FreeSans 224 90 0 0 msb[7]
port 39 nsew signal tristate
flabel metal2 s 5906 29200 5962 30000 0 FreeSans 224 90 0 0 msb[8]
port 40 nsew signal tristate
flabel metal2 s 5354 29200 5410 30000 0 FreeSans 224 90 0 0 msb[9]
port 41 nsew signal tristate
flabel metal2 s 10046 29200 10102 30000 0 FreeSans 224 90 0 0 msb_n[0]
port 42 nsew signal tristate
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 msb_n[10]
port 43 nsew signal tristate
flabel metal2 s 3974 29200 4030 30000 0 FreeSans 224 90 0 0 msb_n[11]
port 44 nsew signal tristate
flabel metal2 s 3422 29200 3478 30000 0 FreeSans 224 90 0 0 msb_n[12]
port 45 nsew signal tristate
flabel metal2 s 2870 29200 2926 30000 0 FreeSans 224 90 0 0 msb_n[13]
port 46 nsew signal tristate
flabel metal2 s 2318 29200 2374 30000 0 FreeSans 224 90 0 0 msb_n[14]
port 47 nsew signal tristate
flabel metal2 s 1766 29200 1822 30000 0 FreeSans 224 90 0 0 msb_n[15]
port 48 nsew signal tristate
flabel metal2 s 9494 29200 9550 30000 0 FreeSans 224 90 0 0 msb_n[1]
port 49 nsew signal tristate
flabel metal2 s 8942 29200 8998 30000 0 FreeSans 224 90 0 0 msb_n[2]
port 50 nsew signal tristate
flabel metal2 s 8390 29200 8446 30000 0 FreeSans 224 90 0 0 msb_n[3]
port 51 nsew signal tristate
flabel metal2 s 7838 29200 7894 30000 0 FreeSans 224 90 0 0 msb_n[4]
port 52 nsew signal tristate
flabel metal2 s 7286 29200 7342 30000 0 FreeSans 224 90 0 0 msb_n[5]
port 53 nsew signal tristate
flabel metal2 s 6734 29200 6790 30000 0 FreeSans 224 90 0 0 msb_n[6]
port 54 nsew signal tristate
flabel metal2 s 6182 29200 6238 30000 0 FreeSans 224 90 0 0 msb_n[7]
port 55 nsew signal tristate
flabel metal2 s 5630 29200 5686 30000 0 FreeSans 224 90 0 0 msb_n[8]
port 56 nsew signal tristate
flabel metal2 s 5078 29200 5134 30000 0 FreeSans 224 90 0 0 msb_n[9]
port 57 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 rst_n
port 58 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 test_mode
port 59 nsew signal input
flabel metal4 s 2657 2128 2977 27792 0 FreeSans 1920 90 0 0 vccd1
port 60 nsew power bidirectional
flabel metal4 s 6084 2128 6404 27792 0 FreeSans 1920 90 0 0 vccd1
port 60 nsew power bidirectional
flabel metal4 s 9511 2128 9831 27792 0 FreeSans 1920 90 0 0 vccd1
port 60 nsew power bidirectional
flabel metal4 s 12938 2128 13258 27792 0 FreeSans 1920 90 0 0 vccd1
port 60 nsew power bidirectional
flabel metal4 s 4370 2128 4690 27792 0 FreeSans 1920 90 0 0 vssd1
port 61 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 27792 0 FreeSans 1920 90 0 0 vssd1
port 61 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 27792 0 FreeSans 1920 90 0 0 vssd1
port 61 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 27792 0 FreeSans 1920 90 0 0 vssd1
port 61 nsew ground bidirectional
rlabel metal1 7958 27744 7958 27744 0 vccd1
rlabel via1 8037 27200 8037 27200 0 vssd1
rlabel metal1 8321 20842 8321 20842 0 _000_
rlabel metal1 6486 5882 6486 5882 0 _001_
rlabel metal1 7355 8534 7355 8534 0 _002_
rlabel metal1 7728 9690 7728 9690 0 _003_
rlabel via1 7401 3502 7401 3502 0 _004_
rlabel metal1 5147 3094 5147 3094 0 _005_
rlabel metal1 6501 3434 6501 3434 0 _006_
rlabel metal1 5883 6698 5883 6698 0 _007_
rlabel metal1 4324 8058 4324 8058 0 _008_
rlabel metal2 4554 9350 4554 9350 0 _009_
rlabel via1 4273 4114 4273 4114 0 _010_
rlabel metal2 8602 11118 8602 11118 0 _011_
rlabel metal1 8367 19346 8367 19346 0 _012_
rlabel metal1 7999 20502 7999 20502 0 _013_
rlabel metal2 8418 15606 8418 15606 0 _014_
rlabel metal1 8183 19754 8183 19754 0 _015_
rlabel metal1 8367 17578 8367 17578 0 _016_
rlabel metal1 8045 13906 8045 13906 0 _017_
rlabel metal2 4370 21318 4370 21318 0 _018_
rlabel metal1 4324 17850 4324 17850 0 _019_
rlabel via1 4926 15062 4926 15062 0 _020_
rlabel metal1 4370 17646 4370 17646 0 _021_
rlabel metal2 3450 21522 3450 21522 0 _022_
rlabel metal2 4370 16966 4370 16966 0 _023_
rlabel metal1 4604 13974 4604 13974 0 _024_
rlabel metal1 5014 20026 5014 20026 0 _025_
rlabel metal1 7038 17204 7038 17204 0 _026_
rlabel metal2 7406 14790 7406 14790 0 _027_
rlabel metal1 6205 19754 6205 19754 0 _028_
rlabel metal1 5612 17850 5612 17850 0 _029_
rlabel metal1 5550 18666 5550 18666 0 _030_
rlabel metal2 7498 14858 7498 14858 0 _031_
rlabel via1 5754 19414 5754 19414 0 _032_
rlabel metal1 5842 12852 5842 12852 0 _033_
rlabel metal1 6854 12716 6854 12716 0 _034_
rlabel metal2 9338 15572 9338 15572 0 _035_
rlabel metal2 8326 6290 8326 6290 0 _036_
rlabel metal1 7728 5202 7728 5202 0 _037_
rlabel metal1 8280 7854 8280 7854 0 _038_
rlabel metal2 9154 8738 9154 8738 0 _039_
rlabel metal1 9108 7990 9108 7990 0 _040_
rlabel metal1 6946 5032 6946 5032 0 _041_
rlabel metal1 7544 8058 7544 8058 0 _042_
rlabel metal2 7498 9350 7498 9350 0 _043_
rlabel metal1 6624 5746 6624 5746 0 _044_
rlabel metal1 7452 5202 7452 5202 0 _045_
rlabel metal2 7498 4556 7498 4556 0 _046_
rlabel metal1 6762 4080 6762 4080 0 _047_
rlabel metal1 6072 3978 6072 3978 0 _048_
rlabel metal1 5888 5338 5888 5338 0 _049_
rlabel metal1 6854 4794 6854 4794 0 _050_
rlabel metal1 6946 2414 6946 2414 0 _051_
rlabel metal2 5566 6902 5566 6902 0 _052_
rlabel metal1 5152 6766 5152 6766 0 _053_
rlabel metal1 5934 8602 5934 8602 0 _054_
rlabel metal1 5428 7514 5428 7514 0 _055_
rlabel metal1 7774 7242 7774 7242 0 _056_
rlabel metal1 4784 6086 4784 6086 0 _057_
rlabel metal1 4662 6358 4662 6358 0 _058_
rlabel metal1 4692 6426 4692 6426 0 _059_
rlabel metal2 5566 6018 5566 6018 0 _060_
rlabel metal2 3818 6494 3818 6494 0 _061_
rlabel metal2 9154 10438 9154 10438 0 _062_
rlabel metal1 7912 12750 7912 12750 0 _063_
rlabel metal1 6210 2482 6210 2482 0 _064_
rlabel metal1 8234 4522 8234 4522 0 _065_
rlabel metal1 9246 12818 9246 12818 0 _066_
rlabel metal1 9292 12954 9292 12954 0 _067_
rlabel metal1 8602 12818 8602 12818 0 _068_
rlabel metal2 8510 13668 8510 13668 0 _069_
rlabel metal1 8510 13294 8510 13294 0 _070_
rlabel metal1 8556 13498 8556 13498 0 _071_
rlabel metal1 8694 4794 8694 4794 0 _072_
rlabel metal1 8740 12410 8740 12410 0 _073_
rlabel metal1 10028 12818 10028 12818 0 _074_
rlabel metal2 9798 13124 9798 13124 0 _075_
rlabel metal1 7636 3162 7636 3162 0 _076_
rlabel metal1 8694 10778 8694 10778 0 _077_
rlabel metal1 5244 12818 5244 12818 0 _078_
rlabel metal1 4922 15980 4922 15980 0 _079_
rlabel metal1 5198 13260 5198 13260 0 _080_
rlabel metal1 6532 13294 6532 13294 0 _081_
rlabel metal1 5750 17714 5750 17714 0 _082_
rlabel metal2 5934 11492 5934 11492 0 _083_
rlabel metal1 4876 14450 4876 14450 0 _084_
rlabel metal2 5750 17714 5750 17714 0 _085_
rlabel metal1 5336 15470 5336 15470 0 _086_
rlabel metal2 4830 14994 4830 14994 0 _087_
rlabel metal1 6394 20434 6394 20434 0 _088_
rlabel metal2 5658 16796 5658 16796 0 _089_
rlabel metal1 4324 14382 4324 14382 0 _090_
rlabel metal2 5934 18700 5934 18700 0 _091_
rlabel metal2 6026 13430 6026 13430 0 _092_
rlabel metal2 2990 1690 2990 1690 0 clk
rlabel metal1 5474 15402 5474 15402 0 clknet_0_clk
rlabel metal2 5290 14144 5290 14144 0 clknet_2_0__leaf_clk
rlabel metal1 7130 11730 7130 11730 0 clknet_2_1__leaf_clk
rlabel metal1 5520 18734 5520 18734 0 clknet_2_2__leaf_clk
rlabel metal1 6210 17170 6210 17170 0 clknet_2_3__leaf_clk
rlabel metal2 8602 7276 8602 7276 0 cnt_r\[0\]
rlabel metal1 8418 8568 8418 8568 0 cnt_r\[1\]
rlabel metal1 7958 7888 7958 7888 0 cnt_r\[2\]
rlabel metal1 8050 4114 8050 4114 0 cnt_r\[3\]
rlabel metal2 6026 5134 6026 5134 0 cnt_r\[4\]
rlabel metal1 6532 4590 6532 4590 0 cnt_r\[5\]
rlabel metal1 5750 8500 5750 8500 0 cnt_r\[6\]
rlabel metal2 6486 10268 6486 10268 0 cnt_r\[7\]
rlabel metal1 5290 9418 5290 9418 0 cnt_r\[8\]
rlabel metal1 4876 3910 4876 3910 0 cnt_r\[9\]
rlabel metal1 14168 3026 14168 3026 0 dac_in[0]
rlabel metal1 13064 2414 13064 2414 0 dac_in[1]
rlabel metal1 11960 2414 11960 2414 0 dac_in[2]
rlabel metal1 10856 2414 10856 2414 0 dac_in[3]
rlabel metal1 9430 2278 9430 2278 0 dac_in[4]
rlabel metal1 8556 2414 8556 2414 0 dac_in[5]
rlabel metal1 7544 2414 7544 2414 0 dac_in[6]
rlabel metal1 6072 2414 6072 2414 0 dac_in[7]
rlabel metal1 4784 2414 4784 2414 0 dac_in[8]
rlabel metal1 3680 2414 3680 2414 0 dac_in[9]
rlabel metal1 13662 2992 13662 2992 0 dummy
rlabel metal1 12650 25738 12650 25738 0 llsb
rlabel metal1 14076 23834 14076 23834 0 llsb_n
rlabel metal1 12880 25126 12880 25126 0 lsb[0]
rlabel metal2 13209 29308 13209 29308 0 lsb[1]
rlabel metal1 12788 25466 12788 25466 0 lsb[2]
rlabel metal1 13156 27098 13156 27098 0 lsb[3]
rlabel metal1 12834 27574 12834 27574 0 lsb[4]
rlabel metal1 11500 27098 11500 27098 0 lsb[5]
rlabel metal1 13524 24378 13524 24378 0 lsb_n[0]
rlabel metal1 13248 25398 13248 25398 0 lsb_n[1]
rlabel metal1 12696 26010 12696 26010 0 lsb_n[2]
rlabel metal1 12558 26758 12558 26758 0 lsb_n[3]
rlabel metal1 11914 26826 11914 26826 0 lsb_n[4]
rlabel metal1 11638 27302 11638 27302 0 lsb_n[5]
rlabel metal1 11408 27574 11408 27574 0 msb[0]
rlabel metal1 3634 27302 3634 27302 0 msb[10]
rlabel metal1 1794 27336 1794 27336 0 msb[11]
rlabel metal1 2852 27098 2852 27098 0 msb[12]
rlabel metal1 2806 26010 2806 26010 0 msb[13]
rlabel metal1 2484 25466 2484 25466 0 msb[14]
rlabel metal2 1971 29308 1971 29308 0 msb[15]
rlabel metal1 10396 27574 10396 27574 0 msb[1]
rlabel metal1 9706 26010 9706 26010 0 msb[2]
rlabel metal2 8510 28441 8510 28441 0 msb[3]
rlabel metal1 7958 27574 7958 27574 0 msb[4]
rlabel metal1 7268 27302 7268 27302 0 msb[5]
rlabel metal2 7038 28434 7038 28434 0 msb[6]
rlabel metal1 6164 27098 6164 27098 0 msb[7]
rlabel metal1 5060 27574 5060 27574 0 msb[8]
rlabel metal1 3266 27540 3266 27540 0 msb[9]
rlabel metal1 10304 27098 10304 27098 0 msb_n[0]
rlabel metal1 3588 26826 3588 26826 0 msb_n[10]
rlabel metal1 4094 25466 4094 25466 0 msb_n[11]
rlabel metal1 2990 26554 2990 26554 0 msb_n[12]
rlabel metal2 2997 29308 2997 29308 0 msb_n[13]
rlabel metal1 2484 24650 2484 24650 0 msb_n[14]
rlabel metal1 1886 24378 1886 24378 0 msb_n[15]
rlabel metal1 9660 26214 9660 26214 0 msb_n[1]
rlabel metal1 9154 27574 9154 27574 0 msb_n[2]
rlabel metal1 8556 27098 8556 27098 0 msb_n[3]
rlabel metal1 7820 27098 7820 27098 0 msb_n[4]
rlabel metal2 7222 28203 7222 28203 0 msb_n[5]
rlabel metal1 5842 27302 5842 27302 0 msb_n[6]
rlabel metal1 5566 26826 5566 26826 0 msb_n[7]
rlabel metal1 5014 27098 5014 27098 0 msb_n[8]
rlabel metal1 3634 27064 3634 27064 0 msb_n[9]
rlabel metal2 14122 5270 14122 5270 0 net1
rlabel metal1 3818 2618 3818 2618 0 net10
rlabel metal2 13478 6562 13478 6562 0 net11
rlabel metal1 3496 2482 3496 2482 0 net12
rlabel metal1 4738 2346 4738 2346 0 net13
rlabel metal1 10672 25874 10672 25874 0 net14
rlabel metal2 14030 24140 14030 24140 0 net15
rlabel metal1 10350 25262 10350 25262 0 net16
rlabel metal1 12972 24786 12972 24786 0 net17
rlabel metal1 12420 25262 12420 25262 0 net18
rlabel metal1 10534 20026 10534 20026 0 net19
rlabel metal1 12742 2618 12742 2618 0 net2
rlabel metal1 10120 17850 10120 17850 0 net20
rlabel metal1 8418 14008 8418 14008 0 net21
rlabel metal2 13754 24922 13754 24922 0 net22
rlabel metal2 13386 25772 13386 25772 0 net23
rlabel metal1 12696 25874 12696 25874 0 net24
rlabel metal1 12880 26962 12880 26962 0 net25
rlabel metal1 12144 26962 12144 26962 0 net26
rlabel metal1 12466 27404 12466 27404 0 net27
rlabel metal2 10258 26860 10258 26860 0 net28
rlabel metal2 2438 26860 2438 26860 0 net29
rlabel metal1 11454 2618 11454 2618 0 net3
rlabel metal2 4278 22848 4278 22848 0 net30
rlabel metal1 2990 20570 2990 20570 0 net31
rlabel metal1 3312 25874 3312 25874 0 net32
rlabel metal1 2668 25262 2668 25262 0 net33
rlabel metal1 1702 24752 1702 24752 0 net34
rlabel metal1 6716 21114 6716 21114 0 net35
rlabel metal1 8464 17306 8464 17306 0 net36
rlabel metal1 8602 25874 8602 25874 0 net37
rlabel metal1 7176 20026 7176 20026 0 net38
rlabel metal1 6302 20570 6302 20570 0 net39
rlabel metal1 10166 4522 10166 4522 0 net4
rlabel metal2 6854 22406 6854 22406 0 net40
rlabel metal1 6394 26316 6394 26316 0 net41
rlabel metal1 4738 19482 4738 19482 0 net42
rlabel metal2 5382 23766 5382 23766 0 net43
rlabel metal2 10350 26758 10350 26758 0 net44
rlabel metal1 4186 26554 4186 26554 0 net45
rlabel metal2 4370 25466 4370 25466 0 net46
rlabel metal1 2714 26384 2714 26384 0 net47
rlabel metal2 3266 25466 3266 25466 0 net48
rlabel metal1 2208 24786 2208 24786 0 net49
rlabel metal1 9798 2618 9798 2618 0 net5
rlabel metal1 1840 24174 1840 24174 0 net50
rlabel metal2 9430 26758 9430 26758 0 net51
rlabel metal2 9154 26996 9154 26996 0 net52
rlabel metal2 8510 26486 8510 26486 0 net53
rlabel metal2 7774 26758 7774 26758 0 net54
rlabel metal2 7038 26758 7038 26758 0 net55
rlabel metal1 5566 27438 5566 27438 0 net56
rlabel metal2 5290 26758 5290 26758 0 net57
rlabel metal1 4968 26486 4968 26486 0 net58
rlabel metal1 4692 25942 4692 25942 0 net59
rlabel metal1 7866 3026 7866 3026 0 net6
rlabel metal1 7360 2618 7360 2618 0 net7
rlabel metal1 6670 2550 6670 2550 0 net8
rlabel via2 4646 2533 4646 2533 0 net9
rlabel metal1 1932 2414 1932 2414 0 rst_n
rlabel metal1 1196 3026 1196 3026 0 test_mode
<< properties >>
string FIXED_BBOX 0 0 16000 30000
<< end >>
