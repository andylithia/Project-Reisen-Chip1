* NGSPICE file created from gated_iref.ext - technology: sky130A

X0 IN_GATED S IN VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X3 IN S IN_GATED VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X1 VSUB SBAR IN_GATED VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X4 IN_GATED SBAR VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X2 IN_GATED OUT VSUB sky130_fd_pr__res_xhigh_po w=350000u l=1.49e+06u
X5 VSUB OUT sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=2.7e+07u
X6 OUT VSUB sky130_fd_pr__cap_mim_m3_2 l=7e+06u w=2.7e+07u
C0 OUT VSUB 45.88fF $ **FLOATING
C1 IN_GATED VSUB 2.05fF $ **FLOATING
