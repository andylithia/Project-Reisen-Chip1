magic
tech sky130A
timestamp 1671631703
<< pwell >>
rect -176 -342 176 342
<< psubdiff >>
rect -158 307 -110 324
rect 110 307 158 324
rect -158 276 -141 307
rect 141 276 158 307
rect -158 -307 -141 -276
rect 141 -307 158 -276
rect -158 -324 -110 -307
rect 110 -324 158 -307
<< psubdiffcont >>
rect -110 307 110 324
rect -158 -276 -141 276
rect 141 -276 158 276
rect -110 -324 110 -307
<< xpolycontact >>
rect -93 -259 -24 -43
rect 24 -259 93 -43
<< ppolyres >>
rect -93 190 93 259
rect -93 -43 -24 190
rect 24 -43 93 190
<< locali >>
rect -158 307 -110 324
rect 110 307 158 324
rect -158 276 -141 307
rect 141 276 158 307
rect -158 -307 -141 -276
rect 141 -307 158 -276
rect -158 -324 -110 -307
rect 110 -324 158 -307
<< properties >>
string FIXED_BBOX -149 -315 149 315
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 2.5 m 1 nx 2 wmin 0.690 lmin 0.50 rho 319.8 val 3.201k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 1 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
