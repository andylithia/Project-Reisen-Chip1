magic
tech sky130A
magscale 1 2
timestamp 1670863211
<< nwell >>
rect 1066 6789 18898 7355
rect 1066 5701 18898 6267
rect 1066 4613 18898 5179
rect 1066 3525 18898 4091
rect 1066 2437 18898 3003
<< obsli1 >>
rect 1104 2159 18860 7633
<< obsm1 >>
rect 1104 2048 19019 7664
<< metal2 >>
rect 1122 9200 1178 10000
rect 3330 9200 3386 10000
rect 5538 9200 5594 10000
rect 7746 9200 7802 10000
rect 9954 9200 10010 10000
rect 12162 9200 12218 10000
rect 14370 9200 14426 10000
rect 16578 9200 16634 10000
rect 18786 9200 18842 10000
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< obsm2 >>
rect 1234 9144 3274 9330
rect 3442 9144 5482 9330
rect 5650 9144 7690 9330
rect 7858 9144 9898 9330
rect 10066 9144 12106 9330
rect 12274 9144 14314 9330
rect 14482 9144 16522 9330
rect 16690 9144 18730 9330
rect 18898 9144 19013 9330
rect 1124 856 19013 9144
rect 1124 800 2446 856
rect 2614 800 7414 856
rect 7582 800 12382 856
rect 12550 800 17350 856
rect 17518 800 19013 856
<< obsm3 >>
rect 3165 2143 19017 7649
<< metal4 >>
rect 3163 2128 3483 7664
rect 5382 2128 5702 7664
rect 7602 2128 7922 7664
rect 9821 2128 10141 7664
rect 12041 2128 12361 7664
rect 14260 2128 14580 7664
rect 16480 2128 16800 7664
rect 18699 2128 19019 7664
<< labels >>
rlabel metal2 s 7470 0 7526 800 6 clk
port 1 nsew signal input
rlabel metal2 s 9954 9200 10010 10000 6 comp
port 2 nsew signal input
rlabel metal2 s 1122 9200 1178 10000 6 dq[0]
port 3 nsew signal output
rlabel metal2 s 3330 9200 3386 10000 6 dq[1]
port 4 nsew signal output
rlabel metal2 s 5538 9200 5594 10000 6 dq[2]
port 5 nsew signal output
rlabel metal2 s 7746 9200 7802 10000 6 dq[3]
port 6 nsew signal output
rlabel metal2 s 12162 9200 12218 10000 6 dq[4]
port 7 nsew signal output
rlabel metal2 s 14370 9200 14426 10000 6 dq[5]
port 8 nsew signal output
rlabel metal2 s 16578 9200 16634 10000 6 dq[6]
port 9 nsew signal output
rlabel metal2 s 18786 9200 18842 10000 6 dq[7]
port 10 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 last_cycle
port 11 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 rst_n
port 12 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 valid
port 13 nsew signal output
rlabel metal4 s 3163 2128 3483 7664 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 7664 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 7664 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 7664 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 7664 6 vssd1
port 15 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 7664 6 vssd1
port 15 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 7664 6 vssd1
port 15 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 7664 6 vssd1
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 297544
string GDS_FILE /home/andylithia/openmpw/Project-Reisen-Chip1_digital/openlane/sarcon_sync/runs/22_12_12_11_39/results/signoff/sarcon_sync.magic.gds
string GDS_START 106056
<< end >>

