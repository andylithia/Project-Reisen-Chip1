magic
tech sky130A
timestamp 1672102605
<< metal1 >>
rect -250 10200 10250 10250
rect -250 -200 -200 10200
rect -50 10000 300 10050
rect -50 0 0 10000
rect 250 0 300 10000
rect -50 -50 300 0
rect 450 10000 800 10050
rect 450 0 500 10000
rect 750 0 800 10000
rect 450 -50 800 0
rect 950 10000 1300 10050
rect 950 0 1000 10000
rect 1250 0 1300 10000
rect 950 -50 1300 0
rect 1450 10000 1800 10050
rect 1450 0 1500 10000
rect 1750 0 1800 10000
rect 1450 -50 1800 0
rect 1950 10000 2300 10050
rect 1950 0 2000 10000
rect 2250 0 2300 10000
rect 1950 -50 2300 0
rect 2450 10000 2800 10050
rect 2450 0 2500 10000
rect 2750 0 2800 10000
rect 2450 -50 2800 0
rect 2950 10000 3300 10050
rect 2950 0 3000 10000
rect 3250 0 3300 10000
rect 2950 -50 3300 0
rect 3450 10000 3800 10050
rect 3450 0 3500 10000
rect 3750 0 3800 10000
rect 3450 -50 3800 0
rect 3950 10000 4300 10050
rect 3950 0 4000 10000
rect 4250 0 4300 10000
rect 3950 -50 4300 0
rect 4450 10000 4800 10050
rect 4450 0 4500 10000
rect 4750 0 4800 10000
rect 4450 -50 4800 0
rect 4950 10000 5300 10050
rect 4950 0 5000 10000
rect 5250 0 5300 10000
rect 4950 -50 5300 0
rect 5450 10000 5800 10050
rect 5450 0 5500 10000
rect 5750 0 5800 10000
rect 5450 -50 5800 0
rect 5950 10000 6300 10050
rect 5950 0 6000 10000
rect 6250 0 6300 10000
rect 5950 -50 6300 0
rect 6450 10000 6800 10050
rect 6450 0 6500 10000
rect 6750 0 6800 10000
rect 6450 -50 6800 0
rect 6950 10000 7300 10050
rect 6950 0 7000 10000
rect 7250 0 7300 10000
rect 6950 -50 7300 0
rect 7450 10000 7800 10050
rect 7450 0 7500 10000
rect 7750 0 7800 10000
rect 7450 -50 7800 0
rect 7950 10000 8300 10050
rect 7950 0 8000 10000
rect 8250 0 8300 10000
rect 7950 -50 8300 0
rect 8450 10000 8800 10050
rect 8450 0 8500 10000
rect 8750 0 8800 10000
rect 8450 -50 8800 0
rect 8950 10000 9300 10050
rect 8950 0 9000 10000
rect 9250 0 9300 10000
rect 8950 -50 9300 0
rect 9450 10000 9800 10050
rect 9450 0 9500 10000
rect 9750 0 9800 10000
rect 9450 -50 9800 0
rect 9950 -50 10050 10050
rect 10200 -200 10250 10200
rect -250 -250 10250 -200
<< via1 >>
rect -200 10050 10200 10200
rect -200 -50 -50 10050
rect 300 -50 450 10050
rect 800 -50 950 10050
rect 1300 -50 1450 10050
rect 1800 -50 1950 10050
rect 2300 -50 2450 10050
rect 2800 -50 2950 10050
rect 3300 -50 3450 10050
rect 3800 -50 3950 10050
rect 4300 -50 4450 10050
rect 4800 -50 4950 10050
rect 5300 -50 5450 10050
rect 5800 -50 5950 10050
rect 6300 -50 6450 10050
rect 6800 -50 6950 10050
rect 7300 -50 7450 10050
rect 7800 -50 7950 10050
rect 8300 -50 8450 10050
rect 8800 -50 8950 10050
rect 9300 -50 9450 10050
rect 9800 -50 9950 10050
rect 10050 -50 10200 10050
rect -200 -200 10200 -50
<< metal2 >>
rect -250 10200 10250 10250
rect -250 -200 -200 10200
rect -50 10000 300 10050
rect -50 0 0 10000
rect 250 0 300 10000
rect -50 -50 300 0
rect 450 10000 800 10050
rect 450 0 500 10000
rect 750 0 800 10000
rect 450 -50 800 0
rect 950 10000 1300 10050
rect 950 0 1000 10000
rect 1250 0 1300 10000
rect 950 -50 1300 0
rect 1450 10000 1800 10050
rect 1450 0 1500 10000
rect 1750 0 1800 10000
rect 1450 -50 1800 0
rect 1950 10000 2300 10050
rect 1950 0 2000 10000
rect 2250 0 2300 10000
rect 1950 -50 2300 0
rect 2450 10000 2800 10050
rect 2450 0 2500 10000
rect 2750 0 2800 10000
rect 2450 -50 2800 0
rect 2950 10000 3300 10050
rect 2950 0 3000 10000
rect 3250 0 3300 10000
rect 2950 -50 3300 0
rect 3450 10000 3800 10050
rect 3450 0 3500 10000
rect 3750 0 3800 10000
rect 3450 -50 3800 0
rect 3950 10000 4300 10050
rect 3950 0 4000 10000
rect 4250 0 4300 10000
rect 3950 -50 4300 0
rect 4450 10000 4800 10050
rect 4450 0 4500 10000
rect 4750 0 4800 10000
rect 4450 -50 4800 0
rect 4950 10000 5300 10050
rect 4950 0 5000 10000
rect 5250 0 5300 10000
rect 4950 -50 5300 0
rect 5450 10000 5800 10050
rect 5450 0 5500 10000
rect 5750 0 5800 10000
rect 5450 -50 5800 0
rect 5950 10000 6300 10050
rect 5950 0 6000 10000
rect 6250 0 6300 10000
rect 5950 -50 6300 0
rect 6450 10000 6800 10050
rect 6450 0 6500 10000
rect 6750 0 6800 10000
rect 6450 -50 6800 0
rect 6950 10000 7300 10050
rect 6950 0 7000 10000
rect 7250 0 7300 10000
rect 6950 -50 7300 0
rect 7450 10000 7800 10050
rect 7450 0 7500 10000
rect 7750 0 7800 10000
rect 7450 -50 7800 0
rect 7950 10000 8300 10050
rect 7950 0 8000 10000
rect 8250 0 8300 10000
rect 7950 -50 8300 0
rect 8450 10000 8800 10050
rect 8450 0 8500 10000
rect 8750 0 8800 10000
rect 8450 -50 8800 0
rect 8950 10000 9300 10050
rect 8950 0 9000 10000
rect 9250 0 9300 10000
rect 8950 -50 9300 0
rect 9450 10000 9800 10050
rect 9450 0 9500 10000
rect 9750 0 9800 10000
rect 9450 -50 9800 0
rect 9950 -50 10050 10050
rect 10200 -200 10250 10200
rect -250 -250 10250 -200
<< via2 >>
rect -200 10050 10200 10200
rect -200 -50 -50 10050
rect 300 -50 450 10050
rect 800 -50 950 10050
rect 1300 -50 1450 10050
rect 1800 -50 1950 10050
rect 2300 -50 2450 10050
rect 2800 -50 2950 10050
rect 3300 -50 3450 10050
rect 3800 -50 3950 10050
rect 4300 -50 4450 10050
rect 4800 -50 4950 10050
rect 5300 -50 5450 10050
rect 5800 -50 5950 10050
rect 6300 -50 6450 10050
rect 6800 -50 6950 10050
rect 7300 -50 7450 10050
rect 7800 -50 7950 10050
rect 8300 -50 8450 10050
rect 8800 -50 8950 10050
rect 9300 -50 9450 10050
rect 9800 -50 9950 10050
rect 10050 -50 10200 10050
rect -200 -200 10200 -50
<< metal3 >>
rect -250 10200 400 10250
rect 9600 10200 10250 10250
rect -250 9600 -200 10200
rect -50 10000 300 10050
rect -250 -200 -200 400
rect -50 0 0 10000
rect 250 0 300 10000
rect 450 10000 800 10050
rect -50 -50 300 0
rect 450 0 500 10000
rect 750 0 800 10000
rect 450 -50 800 0
rect 950 10000 1300 10050
rect 950 0 1000 10000
rect 1250 0 1300 10000
rect 950 -50 1300 0
rect 1450 10000 1800 10050
rect 1450 0 1500 10000
rect 1750 0 1800 10000
rect 1450 -50 1800 0
rect 1950 10000 2300 10050
rect 1950 0 2000 10000
rect 2250 0 2300 10000
rect 1950 -50 2300 0
rect 2450 10000 2800 10050
rect 2450 0 2500 10000
rect 2750 0 2800 10000
rect 2450 -50 2800 0
rect 2950 10000 3300 10050
rect 2950 0 3000 10000
rect 3250 0 3300 10000
rect 2950 -50 3300 0
rect 3450 10000 3800 10050
rect 3450 0 3500 10000
rect 3750 0 3800 10000
rect 3450 -50 3800 0
rect 3950 10000 4300 10050
rect 3950 0 4000 10000
rect 4250 0 4300 10000
rect 3950 -50 4300 0
rect 4450 10000 4800 10050
rect 4450 0 4500 10000
rect 4750 0 4800 10000
rect 4450 -50 4800 0
rect 4950 10000 5300 10050
rect 4950 0 5000 10000
rect 5250 0 5300 10000
rect 4950 -50 5300 0
rect 5450 10000 5800 10050
rect 5450 0 5500 10000
rect 5750 0 5800 10000
rect 5450 -50 5800 0
rect 5950 10000 6300 10050
rect 5950 0 6000 10000
rect 6250 0 6300 10000
rect 5950 -50 6300 0
rect 6450 10000 6800 10050
rect 6450 0 6500 10000
rect 6750 0 6800 10000
rect 6450 -50 6800 0
rect 6950 10000 7300 10050
rect 6950 0 7000 10000
rect 7250 0 7300 10000
rect 6950 -50 7300 0
rect 7450 10000 7800 10050
rect 7450 0 7500 10000
rect 7750 0 7800 10000
rect 7450 -50 7800 0
rect 7950 10000 8300 10050
rect 7950 0 8000 10000
rect 8250 0 8300 10000
rect 7950 -50 8300 0
rect 8450 10000 8800 10050
rect 8450 0 8500 10000
rect 8750 0 8800 10000
rect 8450 -50 8800 0
rect 8950 10000 9300 10050
rect 8950 0 9000 10000
rect 9250 0 9300 10000
rect 8950 -50 9300 0
rect 9450 10000 9800 10050
rect 9450 0 9500 10000
rect 9750 0 9800 10000
rect 9450 -50 9800 0
rect 9950 -50 10050 10050
rect 10200 9600 10250 10200
rect 10200 -200 10250 400
rect -250 -250 400 -200
rect 9600 -250 10250 -200
<< via3 >>
rect 400 10200 9600 10250
rect 400 10050 9600 10200
rect -250 400 -200 9600
rect -200 400 -50 9600
rect 300 150 450 9850
rect 800 -50 950 10050
rect 1300 -50 1450 10050
rect 1800 -50 1950 10050
rect 2300 -50 2450 10050
rect 2800 -50 2950 10050
rect 3300 -50 3450 10050
rect 3800 -50 3950 10050
rect 4300 -50 4450 10050
rect 4800 -50 4950 10050
rect 5300 -50 5450 10050
rect 5800 -50 5950 10050
rect 6300 -50 6450 10050
rect 6800 -50 6950 10050
rect 7300 -50 7450 10050
rect 7800 -50 7950 10050
rect 8300 -50 8450 10050
rect 8800 -50 8950 10050
rect 9300 -50 9450 10050
rect 10050 400 10200 9600
rect 10200 400 10250 9600
rect 400 -200 9600 -50
rect 400 -250 9600 -200
<< metal4 >>
tri 269 10179 360 10270 se
rect 360 10250 9640 10270
rect 360 10179 400 10250
rect 9600 10179 9640 10250
tri 9640 10179 9731 10270 sw
tri 135 10045 269 10179 se
rect 269 10061 301 10179
rect 9699 10061 9731 10179
rect 269 10050 400 10061
rect 9600 10050 9731 10061
rect 269 10045 800 10050
tri -51 9859 135 10045 se
rect 135 10019 800 10045
rect 135 9901 141 10019
rect 259 10000 800 10019
rect 950 10000 1300 10050
rect 1450 10000 1800 10050
rect 1950 10000 2300 10050
rect 2450 10000 2800 10050
rect 2950 10000 3300 10050
rect 3450 10000 3800 10050
rect 3950 10000 4300 10050
rect 4450 10000 4800 10050
rect 4950 10000 5300 10050
rect 5450 10000 5800 10050
rect 5950 10000 6300 10050
rect 6450 10000 6800 10050
rect 6950 10000 7300 10050
rect 7450 10000 7800 10050
rect 7950 10000 8300 10050
rect 8450 10000 8800 10050
rect 8950 10000 9300 10050
rect 9450 10045 9731 10050
tri 9731 10045 9865 10179 sw
rect 9450 10019 9865 10045
rect 259 9901 500 10000
rect 135 9859 500 9901
tri -211 9699 -51 9859 se
rect -51 9741 -19 9859
rect 99 9850 500 9859
rect 99 9741 300 9850
rect -51 9699 300 9741
tri -270 9640 -211 9699 se
rect -211 9640 -179 9699
rect -270 9600 -179 9640
rect -61 9600 300 9699
rect -270 400 -250 9600
rect -50 400 0 9600
tri 0 9505 95 9600 nw
tri 0 400 95 495 sw
rect 250 400 300 9600
rect -270 360 -179 400
tri -270 301 -211 360 ne
rect -211 301 -179 360
rect -61 301 300 400
tri -211 135 -45 301 ne
rect -45 259 300 301
rect -45 141 -19 259
rect 99 150 300 259
rect 450 150 500 9850
rect 99 141 500 150
rect -45 135 500 141
tri -45 -19 109 135 ne
rect 109 99 500 135
rect 109 -19 141 99
rect 259 0 500 99
rect 750 0 800 10000
rect 950 0 1000 10000
rect 1250 0 1300 10000
rect 1450 0 1500 10000
rect 1750 0 1800 10000
rect 1950 0 2000 10000
rect 2250 0 2300 10000
rect 2450 0 2500 10000
rect 2750 0 2800 10000
rect 2950 0 3000 10000
rect 3250 0 3300 10000
rect 3450 0 3500 10000
rect 3750 0 3800 10000
rect 3950 0 4000 10000
rect 4250 0 4300 10000
rect 4450 0 4500 10000
rect 4750 0 4800 10000
rect 4950 0 5000 10000
rect 5250 0 5300 10000
rect 5450 0 5500 10000
rect 5750 0 5800 10000
rect 5950 0 6000 10000
rect 6250 0 6300 10000
rect 6450 0 6500 10000
rect 6750 0 6800 10000
rect 6950 0 7000 10000
rect 7250 0 7300 10000
rect 7450 0 7500 10000
rect 7750 0 7800 10000
rect 7950 0 8000 10000
rect 8250 0 8300 10000
rect 8450 0 8500 10000
rect 8750 0 8800 10000
rect 8950 0 9000 10000
rect 9250 0 9300 10000
rect 9450 9901 9741 10019
rect 9859 9901 9865 10019
rect 9450 9859 9865 9901
tri 9865 9859 10051 10045 sw
rect 9450 9850 9901 9859
rect 9450 200 9500 9850
tri 9655 9640 9865 9850 ne
rect 9865 9741 9901 9850
rect 10019 9741 10051 9859
rect 9865 9699 10051 9741
tri 10051 9699 10211 9859 sw
rect 9865 9640 10061 9699
tri 9865 9505 10000 9640 ne
rect 10000 9600 10061 9640
rect 10179 9640 10211 9699
tri 10211 9640 10270 9699 sw
rect 10179 9600 10270 9640
tri 9865 360 10000 495 se
rect 10000 400 10050 9600
rect 10250 400 10270 9600
rect 10000 360 10061 400
tri 9705 200 9865 360 se
rect 9865 301 10061 360
rect 10179 360 10270 400
rect 10179 301 10211 360
tri 10211 301 10270 360 nw
rect 9865 259 10051 301
rect 9865 200 9901 259
rect 9450 141 9901 200
rect 10019 141 10051 259
tri 10051 141 10211 301 nw
rect 9450 99 9891 141
rect 259 -19 800 0
tri 109 -179 269 -19 ne
rect 269 -50 800 -19
rect 950 -50 1300 0
rect 1450 -50 1800 0
rect 1950 -50 2300 0
rect 2450 -50 2800 0
rect 2950 -50 3300 0
rect 3450 -50 3800 0
rect 3950 -50 4300 0
rect 4450 -50 4800 0
rect 4950 -50 5300 0
rect 5450 -50 5800 0
rect 5950 -50 6300 0
rect 6450 -50 6800 0
rect 6950 -50 7300 0
rect 7450 -50 7800 0
rect 7950 -50 8300 0
rect 8450 -50 8800 0
rect 8950 -50 9300 0
rect 9450 -19 9741 99
rect 9859 -19 9891 99
tri 9891 -19 10051 141 nw
rect 9450 -50 9731 -19
rect 269 -61 400 -50
rect 9600 -61 9731 -50
rect 269 -179 301 -61
rect 9699 -179 9731 -61
tri 9731 -179 9891 -19 nw
tri 269 -270 360 -179 ne
rect 360 -250 400 -179
rect 9600 -250 9640 -179
rect 360 -270 9640 -250
tri 9640 -270 9731 -179 nw
<< via4 >>
rect 301 10061 400 10179
rect 400 10061 419 10179
rect 461 10061 579 10179
rect 621 10061 739 10179
rect 781 10061 899 10179
rect 941 10061 1059 10179
rect 1101 10061 1219 10179
rect 1261 10061 1379 10179
rect 1421 10061 1539 10179
rect 1581 10061 1699 10179
rect 1741 10061 1859 10179
rect 1901 10061 2019 10179
rect 2061 10061 2179 10179
rect 2221 10061 2339 10179
rect 2381 10061 2499 10179
rect 2541 10061 2659 10179
rect 2701 10061 2819 10179
rect 2861 10061 2979 10179
rect 3021 10061 3139 10179
rect 3181 10061 3299 10179
rect 3341 10061 3459 10179
rect 3501 10061 3619 10179
rect 3661 10061 3779 10179
rect 3821 10061 3939 10179
rect 3981 10061 4099 10179
rect 4141 10061 4259 10179
rect 4301 10061 4419 10179
rect 4461 10061 4579 10179
rect 4621 10061 4739 10179
rect 4781 10061 4899 10179
rect 4941 10061 5059 10179
rect 5101 10061 5219 10179
rect 5261 10061 5379 10179
rect 5421 10061 5539 10179
rect 5581 10061 5699 10179
rect 5741 10061 5859 10179
rect 5901 10061 6019 10179
rect 6061 10061 6179 10179
rect 6221 10061 6339 10179
rect 6381 10061 6499 10179
rect 6541 10061 6659 10179
rect 6701 10061 6819 10179
rect 6861 10061 6979 10179
rect 7021 10061 7139 10179
rect 7181 10061 7299 10179
rect 7341 10061 7459 10179
rect 7501 10061 7619 10179
rect 7661 10061 7779 10179
rect 7821 10061 7939 10179
rect 7981 10061 8099 10179
rect 8141 10061 8259 10179
rect 8301 10061 8419 10179
rect 8461 10061 8579 10179
rect 8621 10061 8739 10179
rect 8781 10061 8899 10179
rect 8941 10061 9059 10179
rect 9101 10061 9219 10179
rect 9261 10061 9379 10179
rect 9421 10061 9539 10179
rect 9581 10061 9600 10179
rect 9600 10061 9699 10179
rect 141 9901 259 10019
rect -19 9741 99 9859
rect -179 9600 -61 9699
rect -179 9581 -61 9600
rect -179 9421 -61 9539
rect -179 9261 -61 9379
rect -179 9101 -61 9219
rect -179 8941 -61 9059
rect -179 8781 -61 8899
rect -179 8621 -61 8739
rect -179 8461 -61 8579
rect -179 8301 -61 8419
rect -179 8141 -61 8259
rect -179 7981 -61 8099
rect -179 7821 -61 7939
rect -179 7661 -61 7779
rect -179 7501 -61 7619
rect -179 7341 -61 7459
rect -179 7181 -61 7299
rect -179 7021 -61 7139
rect -179 6861 -61 6979
rect -179 6701 -61 6819
rect -179 6541 -61 6659
rect -179 6381 -61 6499
rect -179 6221 -61 6339
rect -179 6061 -61 6179
rect -179 5901 -61 6019
rect -179 5741 -61 5859
rect -179 5581 -61 5699
rect -179 5421 -61 5539
rect -179 5261 -61 5379
rect -179 5101 -61 5219
rect -179 4941 -61 5059
rect -179 4781 -61 4899
rect -179 4621 -61 4739
rect -179 4461 -61 4579
rect -179 4301 -61 4419
rect -179 4141 -61 4259
rect -179 3981 -61 4099
rect -179 3821 -61 3939
rect -179 3661 -61 3779
rect -179 3501 -61 3619
rect -179 3341 -61 3459
rect -179 3181 -61 3299
rect -179 3021 -61 3139
rect -179 2861 -61 2979
rect -179 2701 -61 2819
rect -179 2541 -61 2659
rect -179 2381 -61 2499
rect -179 2221 -61 2339
rect -179 2061 -61 2179
rect -179 1901 -61 2019
rect -179 1741 -61 1859
rect -179 1581 -61 1699
rect -179 1421 -61 1539
rect -179 1261 -61 1379
rect -179 1101 -61 1219
rect -179 941 -61 1059
rect -179 781 -61 899
rect -179 621 -61 739
rect -179 461 -61 579
rect -179 400 -61 419
rect -179 301 -61 400
rect -19 141 99 259
rect 300 150 450 9850
rect 141 -19 259 99
rect 800 0 950 10000
rect 1300 0 1450 10000
rect 1800 0 1950 10000
rect 2300 0 2450 10000
rect 2800 0 2950 10000
rect 3300 0 3450 10000
rect 3800 0 3950 10000
rect 4300 0 4450 10000
rect 4800 0 4950 10000
rect 5300 0 5450 10000
rect 5800 0 5950 10000
rect 6300 0 6450 10000
rect 6800 0 6950 10000
rect 7300 0 7450 10000
rect 7800 0 7950 10000
rect 8300 0 8450 10000
rect 8800 0 8950 10000
rect 9300 0 9450 10000
rect 9741 9901 9859 10019
rect 9901 9741 10019 9859
rect 10061 9600 10179 9699
rect 10061 9581 10179 9600
rect 10061 9421 10179 9539
rect 10061 9261 10179 9379
rect 10061 9101 10179 9219
rect 10061 8941 10179 9059
rect 10061 8781 10179 8899
rect 10061 8621 10179 8739
rect 10061 8461 10179 8579
rect 10061 8301 10179 8419
rect 10061 8141 10179 8259
rect 10061 7981 10179 8099
rect 10061 7821 10179 7939
rect 10061 7661 10179 7779
rect 10061 7501 10179 7619
rect 10061 7341 10179 7459
rect 10061 7181 10179 7299
rect 10061 7021 10179 7139
rect 10061 6861 10179 6979
rect 10061 6701 10179 6819
rect 10061 6541 10179 6659
rect 10061 6381 10179 6499
rect 10061 6221 10179 6339
rect 10061 6061 10179 6179
rect 10061 5901 10179 6019
rect 10061 5741 10179 5859
rect 10061 5581 10179 5699
rect 10061 5421 10179 5539
rect 10061 5261 10179 5379
rect 10061 5101 10179 5219
rect 10061 4941 10179 5059
rect 10061 4781 10179 4899
rect 10061 4621 10179 4739
rect 10061 4461 10179 4579
rect 10061 4301 10179 4419
rect 10061 4141 10179 4259
rect 10061 3981 10179 4099
rect 10061 3821 10179 3939
rect 10061 3661 10179 3779
rect 10061 3501 10179 3619
rect 10061 3341 10179 3459
rect 10061 3181 10179 3299
rect 10061 3021 10179 3139
rect 10061 2861 10179 2979
rect 10061 2701 10179 2819
rect 10061 2541 10179 2659
rect 10061 2381 10179 2499
rect 10061 2221 10179 2339
rect 10061 2061 10179 2179
rect 10061 1901 10179 2019
rect 10061 1741 10179 1859
rect 10061 1581 10179 1699
rect 10061 1421 10179 1539
rect 10061 1261 10179 1379
rect 10061 1101 10179 1219
rect 10061 941 10179 1059
rect 10061 781 10179 899
rect 10061 621 10179 739
rect 10061 461 10179 579
rect 10061 400 10179 419
rect 10061 301 10179 400
rect 9901 141 10019 259
rect 9741 -19 9859 99
rect 301 -179 400 -61
rect 400 -179 419 -61
rect 461 -179 579 -61
rect 621 -179 739 -61
rect 781 -179 899 -61
rect 941 -179 1059 -61
rect 1101 -179 1219 -61
rect 1261 -179 1379 -61
rect 1421 -179 1539 -61
rect 1581 -179 1699 -61
rect 1741 -179 1859 -61
rect 1901 -179 2019 -61
rect 2061 -179 2179 -61
rect 2221 -179 2339 -61
rect 2381 -179 2499 -61
rect 2541 -179 2659 -61
rect 2701 -179 2819 -61
rect 2861 -179 2979 -61
rect 3021 -179 3139 -61
rect 3181 -179 3299 -61
rect 3341 -179 3459 -61
rect 3501 -179 3619 -61
rect 3661 -179 3779 -61
rect 3821 -179 3939 -61
rect 3981 -179 4099 -61
rect 4141 -179 4259 -61
rect 4301 -179 4419 -61
rect 4461 -179 4579 -61
rect 4621 -179 4739 -61
rect 4781 -179 4899 -61
rect 4941 -179 5059 -61
rect 5101 -179 5219 -61
rect 5261 -179 5379 -61
rect 5421 -179 5539 -61
rect 5581 -179 5699 -61
rect 5741 -179 5859 -61
rect 5901 -179 6019 -61
rect 6061 -179 6179 -61
rect 6221 -179 6339 -61
rect 6381 -179 6499 -61
rect 6541 -179 6659 -61
rect 6701 -179 6819 -61
rect 6861 -179 6979 -61
rect 7021 -179 7139 -61
rect 7181 -179 7299 -61
rect 7341 -179 7459 -61
rect 7501 -179 7619 -61
rect 7661 -179 7779 -61
rect 7821 -179 7939 -61
rect 7981 -179 8099 -61
rect 8141 -179 8259 -61
rect 8301 -179 8419 -61
rect 8461 -179 8579 -61
rect 8621 -179 8739 -61
rect 8781 -179 8899 -61
rect 8941 -179 9059 -61
rect 9101 -179 9219 -61
rect 9261 -179 9379 -61
rect 9421 -179 9539 -61
rect 9581 -179 9600 -61
rect 9600 -179 9699 -61
<< metal5 >>
tri 269 10179 360 10270 se
rect 360 10179 9640 10270
tri 9640 10179 9731 10270 sw
tri 109 10019 269 10179 se
rect 269 10061 301 10179
rect 419 10061 461 10179
rect 579 10061 621 10179
rect 739 10061 781 10179
rect 899 10061 941 10179
rect 1059 10061 1101 10179
rect 1219 10061 1261 10179
rect 1379 10061 1421 10179
rect 1539 10061 1581 10179
rect 1699 10061 1741 10179
rect 1859 10061 1901 10179
rect 2019 10061 2061 10179
rect 2179 10061 2221 10179
rect 2339 10061 2381 10179
rect 2499 10061 2541 10179
rect 2659 10061 2701 10179
rect 2819 10061 2861 10179
rect 2979 10061 3021 10179
rect 3139 10061 3181 10179
rect 3299 10061 3341 10179
rect 3459 10061 3501 10179
rect 3619 10061 3661 10179
rect 3779 10061 3821 10179
rect 3939 10061 3981 10179
rect 4099 10061 4141 10179
rect 4259 10061 4301 10179
rect 4419 10061 4461 10179
rect 4579 10061 4621 10179
rect 4739 10061 4781 10179
rect 4899 10061 4941 10179
rect 5059 10061 5101 10179
rect 5219 10061 5261 10179
rect 5379 10061 5421 10179
rect 5539 10061 5581 10179
rect 5699 10061 5741 10179
rect 5859 10061 5901 10179
rect 6019 10061 6061 10179
rect 6179 10061 6221 10179
rect 6339 10061 6381 10179
rect 6499 10061 6541 10179
rect 6659 10061 6701 10179
rect 6819 10061 6861 10179
rect 6979 10061 7021 10179
rect 7139 10061 7181 10179
rect 7299 10061 7341 10179
rect 7459 10061 7501 10179
rect 7619 10061 7661 10179
rect 7779 10061 7821 10179
rect 7939 10061 7981 10179
rect 8099 10061 8141 10179
rect 8259 10061 8301 10179
rect 8419 10061 8461 10179
rect 8579 10061 8621 10179
rect 8739 10061 8781 10179
rect 8899 10061 8941 10179
rect 9059 10061 9101 10179
rect 9219 10061 9261 10179
rect 9379 10061 9421 10179
rect 9539 10061 9581 10179
rect 9699 10061 9731 10179
rect 269 10019 9731 10061
tri 9731 10019 9891 10179 sw
tri 0 9910 109 10019 se
rect 109 9910 141 10019
tri -51 9859 0 9910 se
rect 0 9901 141 9910
rect 259 10000 9741 10019
rect 259 9901 800 10000
rect 0 9859 800 9901
tri -211 9699 -51 9859 se
rect -51 9741 -19 9859
rect 99 9850 800 9859
rect 99 9741 300 9850
rect -51 9699 300 9741
tri -270 9640 -211 9699 se
rect -211 9640 -179 9699
rect -270 9581 -179 9640
rect -61 9581 300 9699
rect -270 9539 300 9581
rect -270 9421 -179 9539
rect -61 9421 300 9539
rect -270 9379 300 9421
rect -270 9261 -179 9379
rect -61 9261 300 9379
rect -270 9219 300 9261
rect -270 9101 -179 9219
rect -61 9101 300 9219
rect -270 9059 300 9101
rect -270 8941 -179 9059
rect -61 8941 300 9059
rect -270 8899 300 8941
rect -270 8781 -179 8899
rect -61 8781 300 8899
rect -270 8739 300 8781
rect -270 8621 -179 8739
rect -61 8621 300 8739
rect -270 8579 300 8621
rect -270 8461 -179 8579
rect -61 8461 300 8579
rect -270 8419 300 8461
rect -270 8301 -179 8419
rect -61 8301 300 8419
rect -270 8259 300 8301
rect -270 8141 -179 8259
rect -61 8141 300 8259
rect -270 8099 300 8141
rect -270 7981 -179 8099
rect -61 7981 300 8099
rect -270 7939 300 7981
rect -270 7821 -179 7939
rect -61 7821 300 7939
rect -270 7779 300 7821
rect -270 7661 -179 7779
rect -61 7661 300 7779
rect -270 7619 300 7661
rect -270 7501 -179 7619
rect -61 7501 300 7619
rect -270 7459 300 7501
rect -270 7341 -179 7459
rect -61 7341 300 7459
rect -270 7299 300 7341
rect -270 7181 -179 7299
rect -61 7181 300 7299
rect -270 7139 300 7181
rect -270 7021 -179 7139
rect -61 7021 300 7139
rect -270 6979 300 7021
rect -270 6861 -179 6979
rect -61 6861 300 6979
rect -270 6819 300 6861
rect -270 6701 -179 6819
rect -61 6701 300 6819
rect -270 6659 300 6701
rect -270 6541 -179 6659
rect -61 6541 300 6659
rect -270 6499 300 6541
rect -270 6381 -179 6499
rect -61 6381 300 6499
rect -270 6339 300 6381
rect -270 6221 -179 6339
rect -61 6221 300 6339
rect -270 6179 300 6221
rect -270 6061 -179 6179
rect -61 6061 300 6179
rect -270 6019 300 6061
rect -270 5901 -179 6019
rect -61 5901 300 6019
rect -270 5859 300 5901
rect -270 5741 -179 5859
rect -61 5741 300 5859
rect -270 5699 300 5741
rect -270 5581 -179 5699
rect -61 5581 300 5699
rect -270 5539 300 5581
rect -270 5421 -179 5539
rect -61 5421 300 5539
rect -270 5379 300 5421
rect -270 5261 -179 5379
rect -61 5261 300 5379
rect -270 5219 300 5261
rect -270 5101 -179 5219
rect -61 5101 300 5219
rect -270 5059 300 5101
rect -270 4941 -179 5059
rect -61 4941 300 5059
rect -270 4899 300 4941
rect -270 4781 -179 4899
rect -61 4781 300 4899
rect -270 4739 300 4781
rect -270 4621 -179 4739
rect -61 4621 300 4739
rect -270 4579 300 4621
rect -270 4461 -179 4579
rect -61 4461 300 4579
rect -270 4419 300 4461
rect -270 4301 -179 4419
rect -61 4301 300 4419
rect -270 4259 300 4301
rect -270 4141 -179 4259
rect -61 4141 300 4259
rect -270 4099 300 4141
rect -270 3981 -179 4099
rect -61 3981 300 4099
rect -270 3939 300 3981
rect -270 3821 -179 3939
rect -61 3821 300 3939
rect -270 3779 300 3821
rect -270 3661 -179 3779
rect -61 3661 300 3779
rect -270 3619 300 3661
rect -270 3501 -179 3619
rect -61 3501 300 3619
rect -270 3459 300 3501
rect -270 3341 -179 3459
rect -61 3341 300 3459
rect -270 3299 300 3341
rect -270 3181 -179 3299
rect -61 3181 300 3299
rect -270 3139 300 3181
rect -270 3021 -179 3139
rect -61 3021 300 3139
rect -270 2979 300 3021
rect -270 2861 -179 2979
rect -61 2861 300 2979
rect -270 2819 300 2861
rect -270 2701 -179 2819
rect -61 2701 300 2819
rect -270 2659 300 2701
rect -270 2541 -179 2659
rect -61 2541 300 2659
rect -270 2499 300 2541
rect -270 2381 -179 2499
rect -61 2381 300 2499
rect -270 2339 300 2381
rect -270 2221 -179 2339
rect -61 2221 300 2339
rect -270 2179 300 2221
rect -270 2061 -179 2179
rect -61 2061 300 2179
rect -270 2019 300 2061
rect -270 1901 -179 2019
rect -61 1901 300 2019
rect -270 1859 300 1901
rect -270 1741 -179 1859
rect -61 1741 300 1859
rect -270 1699 300 1741
rect -270 1581 -179 1699
rect -61 1581 300 1699
rect -270 1539 300 1581
rect -270 1421 -179 1539
rect -61 1421 300 1539
rect -270 1379 300 1421
rect -270 1261 -179 1379
rect -61 1261 300 1379
rect -270 1219 300 1261
rect -270 1101 -179 1219
rect -61 1101 300 1219
rect -270 1059 300 1101
rect -270 941 -179 1059
rect -61 941 300 1059
rect -270 899 300 941
rect -270 781 -179 899
rect -61 781 300 899
rect -270 739 300 781
rect -270 621 -179 739
rect -61 621 300 739
rect -270 579 300 621
rect -270 461 -179 579
rect -61 461 300 579
rect -270 419 300 461
rect -270 360 -179 419
tri -270 301 -211 360 ne
rect -211 301 -179 360
rect -61 301 300 419
tri -211 141 -51 301 ne
rect -51 259 300 301
rect -51 141 -19 259
rect 99 150 300 259
rect 450 150 800 9850
rect 99 141 800 150
tri -51 -19 109 141 ne
rect 109 99 800 141
rect 109 -19 141 99
rect 259 0 800 99
rect 950 0 1300 10000
rect 1450 0 1800 10000
rect 1950 0 2300 10000
rect 2450 0 2800 10000
rect 2950 0 3300 10000
rect 3450 0 3800 10000
rect 3950 0 4300 10000
rect 4450 0 4800 10000
rect 4950 0 5300 10000
rect 5450 0 5800 10000
rect 5950 0 6300 10000
rect 6450 0 6800 10000
rect 6950 0 7300 10000
rect 7450 0 7800 10000
rect 7950 0 8300 10000
rect 8450 0 8800 10000
rect 8950 0 9300 10000
rect 9450 9901 9741 10000
rect 9859 9901 9891 10019
rect 9450 9859 9891 9901
tri 9891 9859 10051 10019 sw
rect 9450 9741 9901 9859
rect 10019 9741 10051 9859
rect 9450 9699 10051 9741
tri 10051 9699 10211 9859 sw
rect 9450 9581 10061 9699
rect 10179 9640 10211 9699
tri 10211 9640 10270 9699 sw
rect 10179 9581 10270 9640
rect 9450 9539 10270 9581
rect 9450 9421 10061 9539
rect 10179 9421 10270 9539
rect 9450 9379 10270 9421
rect 9450 9261 10061 9379
rect 10179 9261 10270 9379
rect 9450 9219 10270 9261
rect 9450 9101 10061 9219
rect 10179 9101 10270 9219
rect 9450 9059 10270 9101
rect 9450 8941 10061 9059
rect 10179 8941 10270 9059
rect 9450 8899 10270 8941
rect 9450 8781 10061 8899
rect 10179 8781 10270 8899
rect 9450 8739 10270 8781
rect 9450 8621 10061 8739
rect 10179 8621 10270 8739
rect 9450 8579 10270 8621
rect 9450 8461 10061 8579
rect 10179 8461 10270 8579
rect 9450 8419 10270 8461
rect 9450 8301 10061 8419
rect 10179 8301 10270 8419
rect 9450 8259 10270 8301
rect 9450 8141 10061 8259
rect 10179 8141 10270 8259
rect 9450 8099 10270 8141
rect 9450 7981 10061 8099
rect 10179 7981 10270 8099
rect 9450 7939 10270 7981
rect 9450 7821 10061 7939
rect 10179 7821 10270 7939
rect 9450 7779 10270 7821
rect 9450 7661 10061 7779
rect 10179 7661 10270 7779
rect 9450 7619 10270 7661
rect 9450 7501 10061 7619
rect 10179 7501 10270 7619
rect 9450 7459 10270 7501
rect 9450 7341 10061 7459
rect 10179 7341 10270 7459
rect 9450 7299 10270 7341
rect 9450 7181 10061 7299
rect 10179 7181 10270 7299
rect 9450 7139 10270 7181
rect 9450 7021 10061 7139
rect 10179 7021 10270 7139
rect 9450 6979 10270 7021
rect 9450 6861 10061 6979
rect 10179 6861 10270 6979
rect 9450 6819 10270 6861
rect 9450 6701 10061 6819
rect 10179 6701 10270 6819
rect 9450 6659 10270 6701
rect 9450 6541 10061 6659
rect 10179 6541 10270 6659
rect 9450 6499 10270 6541
rect 9450 6381 10061 6499
rect 10179 6381 10270 6499
rect 9450 6339 10270 6381
rect 9450 6221 10061 6339
rect 10179 6221 10270 6339
rect 9450 6179 10270 6221
rect 9450 6061 10061 6179
rect 10179 6061 10270 6179
rect 9450 6019 10270 6061
rect 9450 5901 10061 6019
rect 10179 5901 10270 6019
rect 9450 5859 10270 5901
rect 9450 5741 10061 5859
rect 10179 5741 10270 5859
rect 9450 5699 10270 5741
rect 9450 5581 10061 5699
rect 10179 5581 10270 5699
rect 9450 5539 10270 5581
rect 9450 5421 10061 5539
rect 10179 5421 10270 5539
rect 9450 5379 10270 5421
rect 9450 5261 10061 5379
rect 10179 5261 10270 5379
rect 9450 5219 10270 5261
rect 9450 5101 10061 5219
rect 10179 5101 10270 5219
rect 9450 5059 10270 5101
rect 9450 4941 10061 5059
rect 10179 4941 10270 5059
rect 9450 4899 10270 4941
rect 9450 4781 10061 4899
rect 10179 4781 10270 4899
rect 9450 4739 10270 4781
rect 9450 4621 10061 4739
rect 10179 4621 10270 4739
rect 9450 4579 10270 4621
rect 9450 4461 10061 4579
rect 10179 4461 10270 4579
rect 9450 4419 10270 4461
rect 9450 4301 10061 4419
rect 10179 4301 10270 4419
rect 9450 4259 10270 4301
rect 9450 4141 10061 4259
rect 10179 4141 10270 4259
rect 9450 4099 10270 4141
rect 9450 3981 10061 4099
rect 10179 3981 10270 4099
rect 9450 3939 10270 3981
rect 9450 3821 10061 3939
rect 10179 3821 10270 3939
rect 9450 3779 10270 3821
rect 9450 3661 10061 3779
rect 10179 3661 10270 3779
rect 9450 3619 10270 3661
rect 9450 3501 10061 3619
rect 10179 3501 10270 3619
rect 9450 3459 10270 3501
rect 9450 3341 10061 3459
rect 10179 3341 10270 3459
rect 9450 3299 10270 3341
rect 9450 3181 10061 3299
rect 10179 3181 10270 3299
rect 9450 3139 10270 3181
rect 9450 3021 10061 3139
rect 10179 3021 10270 3139
rect 9450 2979 10270 3021
rect 9450 2861 10061 2979
rect 10179 2861 10270 2979
rect 9450 2819 10270 2861
rect 9450 2701 10061 2819
rect 10179 2701 10270 2819
rect 9450 2659 10270 2701
rect 9450 2541 10061 2659
rect 10179 2541 10270 2659
rect 9450 2499 10270 2541
rect 9450 2381 10061 2499
rect 10179 2381 10270 2499
rect 9450 2339 10270 2381
rect 9450 2221 10061 2339
rect 10179 2221 10270 2339
rect 9450 2179 10270 2221
rect 9450 2061 10061 2179
rect 10179 2061 10270 2179
rect 9450 2019 10270 2061
rect 9450 1901 10061 2019
rect 10179 1901 10270 2019
rect 9450 1859 10270 1901
rect 9450 1741 10061 1859
rect 10179 1741 10270 1859
rect 9450 1699 10270 1741
rect 9450 1581 10061 1699
rect 10179 1581 10270 1699
rect 9450 1539 10270 1581
rect 9450 1421 10061 1539
rect 10179 1421 10270 1539
rect 9450 1379 10270 1421
rect 9450 1261 10061 1379
rect 10179 1261 10270 1379
rect 9450 1219 10270 1261
rect 9450 1101 10061 1219
rect 10179 1101 10270 1219
rect 9450 1059 10270 1101
rect 9450 941 10061 1059
rect 10179 941 10270 1059
rect 9450 899 10270 941
rect 9450 781 10061 899
rect 10179 781 10270 899
rect 9450 739 10270 781
rect 9450 621 10061 739
rect 10179 621 10270 739
rect 9450 579 10270 621
rect 9450 461 10061 579
rect 10179 461 10270 579
rect 9450 419 10270 461
rect 9450 301 10061 419
rect 10179 360 10270 419
rect 10179 301 10211 360
tri 10211 301 10270 360 nw
rect 9450 259 10051 301
rect 9450 141 9901 259
rect 10019 141 10051 259
tri 10051 141 10211 301 nw
rect 9450 99 9891 141
rect 9450 0 9741 99
rect 259 -19 9741 0
rect 9859 -19 9891 99
tri 9891 -19 10051 141 nw
tri 109 -179 269 -19 ne
rect 269 -61 9731 -19
rect 269 -179 301 -61
rect 419 -179 461 -61
rect 579 -179 621 -61
rect 739 -179 781 -61
rect 899 -179 941 -61
rect 1059 -179 1101 -61
rect 1219 -179 1261 -61
rect 1379 -179 1421 -61
rect 1539 -179 1581 -61
rect 1699 -179 1741 -61
rect 1859 -179 1901 -61
rect 2019 -179 2061 -61
rect 2179 -179 2221 -61
rect 2339 -179 2381 -61
rect 2499 -179 2541 -61
rect 2659 -179 2701 -61
rect 2819 -179 2861 -61
rect 2979 -179 3021 -61
rect 3139 -179 3181 -61
rect 3299 -179 3341 -61
rect 3459 -179 3501 -61
rect 3619 -179 3661 -61
rect 3779 -179 3821 -61
rect 3939 -179 3981 -61
rect 4099 -179 4141 -61
rect 4259 -179 4301 -61
rect 4419 -179 4461 -61
rect 4579 -179 4621 -61
rect 4739 -179 4781 -61
rect 4899 -179 4941 -61
rect 5059 -179 5101 -61
rect 5219 -179 5261 -61
rect 5379 -179 5421 -61
rect 5539 -179 5581 -61
rect 5699 -179 5741 -61
rect 5859 -179 5901 -61
rect 6019 -179 6061 -61
rect 6179 -179 6221 -61
rect 6339 -179 6381 -61
rect 6499 -179 6541 -61
rect 6659 -179 6701 -61
rect 6819 -179 6861 -61
rect 6979 -179 7021 -61
rect 7139 -179 7181 -61
rect 7299 -179 7341 -61
rect 7459 -179 7501 -61
rect 7619 -179 7661 -61
rect 7779 -179 7821 -61
rect 7939 -179 7981 -61
rect 8099 -179 8141 -61
rect 8259 -179 8301 -61
rect 8419 -179 8461 -61
rect 8579 -179 8621 -61
rect 8739 -179 8781 -61
rect 8899 -179 8941 -61
rect 9059 -179 9101 -61
rect 9219 -179 9261 -61
rect 9379 -179 9421 -61
rect 9539 -179 9581 -61
rect 9699 -179 9731 -61
tri 9731 -179 9891 -19 nw
tri 269 -270 360 -179 ne
rect 360 -270 9640 -179
tri 9640 -270 9731 -179 nw
<< glass >>
tri 0 9505 495 10000 se
rect 495 9505 9505 10000
tri 9505 9505 10000 10000 sw
rect 0 495 10000 9505
tri 0 0 495 495 ne
rect 495 0 9505 495
tri 9505 0 10000 495 nw
<< labels >>
flabel metal5 s 5000 5000 5000 5000 0 FreeSans 10000 0 0 0 PAD
port 1 nsew
<< end >>
