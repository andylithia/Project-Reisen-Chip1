magic
tech sky130A
magscale 1 2
timestamp 1671855415
<< nwell >>
rect -2253 -3134 1857 -696
<< pwell >>
rect -2490 -5634 -1448 -3214
rect -1325 -4310 929 -3390
rect 1051 -3582 2093 -3214
rect -3760 -6214 -2840 -5748
rect -3760 -6218 -3002 -6214
rect -2956 -6218 -2840 -6214
rect -3760 -6534 -2840 -6218
rect -3760 -6640 -2928 -6534
rect -2919 -6640 -2840 -6534
rect -3760 -6882 -2840 -6640
rect -1281 -6750 885 -4330
rect 1051 -4950 2796 -3582
rect 1051 -5634 2093 -4950
<< nmos >>
rect -2294 -5424 -2234 -3424
rect -2176 -5424 -2116 -3424
rect -2058 -5424 -1998 -3424
rect -1940 -5424 -1880 -3424
rect -1822 -5424 -1762 -3424
rect -1704 -5424 -1644 -3424
rect -3550 -5978 -3050 -5948
rect -3550 -6074 -3050 -6044
rect -3550 -6170 -3050 -6140
rect -3550 -6266 -3050 -6236
rect -1085 -6540 -685 -4540
rect -627 -6540 -227 -4540
rect -169 -6540 231 -4540
rect 289 -6540 689 -4540
rect 1247 -5424 1307 -3424
rect 1365 -5424 1425 -3424
rect 1483 -5424 1543 -3424
rect 1601 -5424 1661 -3424
rect 1719 -5424 1779 -3424
rect 1837 -5424 1897 -3424
<< pmos >>
rect -2057 -2915 -1997 -915
rect -1939 -2915 -1879 -915
rect -1821 -2915 -1761 -915
rect -1703 -2915 -1643 -915
rect -1585 -2915 -1525 -915
rect -1467 -2915 -1407 -915
rect -1349 -2915 -1289 -915
rect -1231 -2915 -1171 -915
rect -1113 -2915 -1053 -915
rect -995 -2915 -935 -915
rect -877 -2915 -817 -915
rect -759 -2915 -699 -915
rect -641 -2915 -581 -915
rect -523 -2915 -463 -915
rect -405 -2915 -345 -915
rect -287 -2915 -227 -915
rect -169 -2915 -109 -915
rect -51 -2915 9 -915
rect 67 -2915 127 -915
rect 185 -2915 245 -915
rect 303 -2915 363 -915
rect 421 -2915 481 -915
rect 539 -2915 599 -915
rect 657 -2915 717 -915
rect 775 -2915 835 -915
rect 893 -2915 953 -915
rect 1011 -2915 1071 -915
rect 1129 -2915 1189 -915
rect 1247 -2915 1307 -915
rect 1365 -2915 1425 -915
rect 1483 -2915 1543 -915
rect 1601 -2915 1661 -915
<< nmoslvt >>
rect -1125 -4100 -1095 -3600
rect -1029 -4100 -999 -3600
rect -933 -4100 -903 -3600
rect -837 -4100 -807 -3600
rect -741 -4100 -711 -3600
rect -645 -4100 -615 -3600
rect -549 -4100 -519 -3600
rect -453 -4100 -423 -3600
rect -357 -4100 -327 -3600
rect -261 -4100 -231 -3600
rect -165 -4100 -135 -3600
rect -69 -4100 -39 -3600
rect 27 -4100 57 -3600
rect 123 -4100 153 -3600
rect 219 -4100 249 -3600
rect 315 -4100 345 -3600
rect 411 -4100 441 -3600
rect 507 -4100 537 -3600
rect 603 -4100 633 -3600
rect 699 -4100 729 -3600
<< ndiff >>
rect -2352 -3436 -2294 -3424
rect -2352 -5412 -2340 -3436
rect -2306 -5412 -2294 -3436
rect -2352 -5424 -2294 -5412
rect -2234 -3436 -2176 -3424
rect -2234 -5412 -2222 -3436
rect -2188 -5412 -2176 -3436
rect -2234 -5424 -2176 -5412
rect -2116 -3436 -2058 -3424
rect -2116 -5412 -2104 -3436
rect -2070 -5412 -2058 -3436
rect -2116 -5424 -2058 -5412
rect -1998 -3436 -1940 -3424
rect -1998 -5412 -1986 -3436
rect -1952 -5412 -1940 -3436
rect -1998 -5424 -1940 -5412
rect -1880 -3436 -1822 -3424
rect -1880 -5412 -1868 -3436
rect -1834 -5412 -1822 -3436
rect -1880 -5424 -1822 -5412
rect -1762 -3436 -1704 -3424
rect -1762 -5412 -1750 -3436
rect -1716 -5412 -1704 -3436
rect -1762 -5424 -1704 -5412
rect -1644 -3436 -1586 -3424
rect -1644 -5412 -1632 -3436
rect -1598 -5412 -1586 -3436
rect -1644 -5424 -1586 -5412
rect -1187 -3612 -1125 -3600
rect -1187 -4088 -1175 -3612
rect -1141 -4088 -1125 -3612
rect -1187 -4100 -1125 -4088
rect -1095 -3612 -1029 -3600
rect -1095 -4088 -1079 -3612
rect -1045 -4088 -1029 -3612
rect -1095 -4100 -1029 -4088
rect -999 -3612 -933 -3600
rect -999 -4088 -983 -3612
rect -949 -4088 -933 -3612
rect -999 -4100 -933 -4088
rect -903 -3612 -837 -3600
rect -903 -4088 -887 -3612
rect -853 -4088 -837 -3612
rect -903 -4100 -837 -4088
rect -807 -3612 -741 -3600
rect -807 -4088 -791 -3612
rect -757 -4088 -741 -3612
rect -807 -4100 -741 -4088
rect -711 -3612 -645 -3600
rect -711 -4088 -695 -3612
rect -661 -4088 -645 -3612
rect -711 -4100 -645 -4088
rect -615 -3612 -549 -3600
rect -615 -4088 -599 -3612
rect -565 -4088 -549 -3612
rect -615 -4100 -549 -4088
rect -519 -3612 -453 -3600
rect -519 -4088 -503 -3612
rect -469 -4088 -453 -3612
rect -519 -4100 -453 -4088
rect -423 -3612 -357 -3600
rect -423 -4088 -407 -3612
rect -373 -4088 -357 -3612
rect -423 -4100 -357 -4088
rect -327 -3612 -261 -3600
rect -327 -4088 -311 -3612
rect -277 -4088 -261 -3612
rect -327 -4100 -261 -4088
rect -231 -3612 -165 -3600
rect -231 -4088 -215 -3612
rect -181 -4088 -165 -3612
rect -231 -4100 -165 -4088
rect -135 -3612 -69 -3600
rect -135 -4088 -119 -3612
rect -85 -4088 -69 -3612
rect -135 -4100 -69 -4088
rect -39 -3612 27 -3600
rect -39 -4088 -23 -3612
rect 11 -4088 27 -3612
rect -39 -4100 27 -4088
rect 57 -3612 123 -3600
rect 57 -4088 73 -3612
rect 107 -4088 123 -3612
rect 57 -4100 123 -4088
rect 153 -3612 219 -3600
rect 153 -4088 169 -3612
rect 203 -4088 219 -3612
rect 153 -4100 219 -4088
rect 249 -3612 315 -3600
rect 249 -4088 265 -3612
rect 299 -4088 315 -3612
rect 249 -4100 315 -4088
rect 345 -3612 411 -3600
rect 345 -4088 361 -3612
rect 395 -4088 411 -3612
rect 345 -4100 411 -4088
rect 441 -3612 507 -3600
rect 441 -4088 457 -3612
rect 491 -4088 507 -3612
rect 441 -4100 507 -4088
rect 537 -3612 603 -3600
rect 537 -4088 553 -3612
rect 587 -4088 603 -3612
rect 537 -4100 603 -4088
rect 633 -3612 699 -3600
rect 633 -4088 649 -3612
rect 683 -4088 699 -3612
rect 633 -4100 699 -4088
rect 729 -3612 791 -3600
rect 729 -4088 745 -3612
rect 779 -4088 791 -3612
rect 729 -4100 791 -4088
rect -3550 -5898 -3050 -5886
rect -3550 -5932 -3538 -5898
rect -3062 -5932 -3050 -5898
rect -3550 -5948 -3050 -5932
rect -3550 -5994 -3050 -5978
rect -3550 -6028 -3538 -5994
rect -3062 -6028 -3050 -5994
rect -3550 -6044 -3050 -6028
rect -3550 -6090 -3050 -6074
rect -3550 -6124 -3538 -6090
rect -3062 -6124 -3050 -6090
rect -3550 -6140 -3050 -6124
rect -3550 -6186 -3050 -6170
rect -3550 -6220 -3538 -6186
rect -3062 -6220 -3050 -6186
rect -3550 -6236 -3050 -6220
rect -3550 -6282 -3050 -6266
rect -3550 -6316 -3538 -6282
rect -3062 -6316 -3050 -6282
rect -3550 -6328 -3050 -6316
rect -1143 -4552 -1085 -4540
rect -1143 -6528 -1131 -4552
rect -1097 -6528 -1085 -4552
rect -1143 -6540 -1085 -6528
rect -685 -4552 -627 -4540
rect -685 -6528 -673 -4552
rect -639 -6528 -627 -4552
rect -685 -6540 -627 -6528
rect -227 -4552 -169 -4540
rect -227 -6528 -215 -4552
rect -181 -6528 -169 -4552
rect -227 -6540 -169 -6528
rect 231 -4552 289 -4540
rect 231 -6528 243 -4552
rect 277 -6528 289 -4552
rect 231 -6540 289 -6528
rect 689 -4552 747 -4540
rect 689 -6528 701 -4552
rect 735 -6528 747 -4552
rect 689 -6540 747 -6528
rect 1189 -3436 1247 -3424
rect 1189 -5412 1201 -3436
rect 1235 -5412 1247 -3436
rect 1189 -5424 1247 -5412
rect 1307 -3436 1365 -3424
rect 1307 -5412 1319 -3436
rect 1353 -5412 1365 -3436
rect 1307 -5424 1365 -5412
rect 1425 -3436 1483 -3424
rect 1425 -5412 1437 -3436
rect 1471 -5412 1483 -3436
rect 1425 -5424 1483 -5412
rect 1543 -3436 1601 -3424
rect 1543 -5412 1555 -3436
rect 1589 -5412 1601 -3436
rect 1543 -5424 1601 -5412
rect 1661 -3436 1719 -3424
rect 1661 -5412 1673 -3436
rect 1707 -5412 1719 -3436
rect 1661 -5424 1719 -5412
rect 1779 -3436 1837 -3424
rect 1779 -5412 1791 -3436
rect 1825 -5412 1837 -3436
rect 1779 -5424 1837 -5412
rect 1897 -3436 1955 -3424
rect 1897 -5412 1909 -3436
rect 1943 -5412 1955 -3436
rect 1897 -5424 1955 -5412
<< pdiff >>
rect -2115 -927 -2057 -915
rect -2115 -2903 -2103 -927
rect -2069 -2903 -2057 -927
rect -2115 -2915 -2057 -2903
rect -1997 -927 -1939 -915
rect -1997 -2903 -1985 -927
rect -1951 -2903 -1939 -927
rect -1997 -2915 -1939 -2903
rect -1879 -927 -1821 -915
rect -1879 -2903 -1867 -927
rect -1833 -2903 -1821 -927
rect -1879 -2915 -1821 -2903
rect -1761 -927 -1703 -915
rect -1761 -2903 -1749 -927
rect -1715 -2903 -1703 -927
rect -1761 -2915 -1703 -2903
rect -1643 -927 -1585 -915
rect -1643 -2903 -1631 -927
rect -1597 -2903 -1585 -927
rect -1643 -2915 -1585 -2903
rect -1525 -927 -1467 -915
rect -1525 -2903 -1513 -927
rect -1479 -2903 -1467 -927
rect -1525 -2915 -1467 -2903
rect -1407 -927 -1349 -915
rect -1407 -2903 -1395 -927
rect -1361 -2903 -1349 -927
rect -1407 -2915 -1349 -2903
rect -1289 -927 -1231 -915
rect -1289 -2903 -1277 -927
rect -1243 -2903 -1231 -927
rect -1289 -2915 -1231 -2903
rect -1171 -927 -1113 -915
rect -1171 -2903 -1159 -927
rect -1125 -2903 -1113 -927
rect -1171 -2915 -1113 -2903
rect -1053 -927 -995 -915
rect -1053 -2903 -1041 -927
rect -1007 -2903 -995 -927
rect -1053 -2915 -995 -2903
rect -935 -927 -877 -915
rect -935 -2903 -923 -927
rect -889 -2903 -877 -927
rect -935 -2915 -877 -2903
rect -817 -927 -759 -915
rect -817 -2903 -805 -927
rect -771 -2903 -759 -927
rect -817 -2915 -759 -2903
rect -699 -927 -641 -915
rect -699 -2903 -687 -927
rect -653 -2903 -641 -927
rect -699 -2915 -641 -2903
rect -581 -927 -523 -915
rect -581 -2903 -569 -927
rect -535 -2903 -523 -927
rect -581 -2915 -523 -2903
rect -463 -927 -405 -915
rect -463 -2903 -451 -927
rect -417 -2903 -405 -927
rect -463 -2915 -405 -2903
rect -345 -927 -287 -915
rect -345 -2903 -333 -927
rect -299 -2903 -287 -927
rect -345 -2915 -287 -2903
rect -227 -927 -169 -915
rect -227 -2903 -215 -927
rect -181 -2903 -169 -927
rect -227 -2915 -169 -2903
rect -109 -927 -51 -915
rect -109 -2903 -97 -927
rect -63 -2903 -51 -927
rect -109 -2915 -51 -2903
rect 9 -927 67 -915
rect 9 -2903 21 -927
rect 55 -2903 67 -927
rect 9 -2915 67 -2903
rect 127 -927 185 -915
rect 127 -2903 139 -927
rect 173 -2903 185 -927
rect 127 -2915 185 -2903
rect 245 -927 303 -915
rect 245 -2903 257 -927
rect 291 -2903 303 -927
rect 245 -2915 303 -2903
rect 363 -927 421 -915
rect 363 -2903 375 -927
rect 409 -2903 421 -927
rect 363 -2915 421 -2903
rect 481 -927 539 -915
rect 481 -2903 493 -927
rect 527 -2903 539 -927
rect 481 -2915 539 -2903
rect 599 -927 657 -915
rect 599 -2903 611 -927
rect 645 -2903 657 -927
rect 599 -2915 657 -2903
rect 717 -927 775 -915
rect 717 -2903 729 -927
rect 763 -2903 775 -927
rect 717 -2915 775 -2903
rect 835 -927 893 -915
rect 835 -2903 847 -927
rect 881 -2903 893 -927
rect 835 -2915 893 -2903
rect 953 -927 1011 -915
rect 953 -2903 965 -927
rect 999 -2903 1011 -927
rect 953 -2915 1011 -2903
rect 1071 -927 1129 -915
rect 1071 -2903 1083 -927
rect 1117 -2903 1129 -927
rect 1071 -2915 1129 -2903
rect 1189 -927 1247 -915
rect 1189 -2903 1201 -927
rect 1235 -2903 1247 -927
rect 1189 -2915 1247 -2903
rect 1307 -927 1365 -915
rect 1307 -2903 1319 -927
rect 1353 -2903 1365 -927
rect 1307 -2915 1365 -2903
rect 1425 -927 1483 -915
rect 1425 -2903 1437 -927
rect 1471 -2903 1483 -927
rect 1425 -2915 1483 -2903
rect 1543 -927 1601 -915
rect 1543 -2903 1555 -927
rect 1589 -2903 1601 -927
rect 1543 -2915 1601 -2903
rect 1661 -927 1719 -915
rect 1661 -2903 1673 -927
rect 1707 -2903 1719 -927
rect 1661 -2915 1719 -2903
<< ndiffc >>
rect -2340 -5412 -2306 -3436
rect -2222 -5412 -2188 -3436
rect -2104 -5412 -2070 -3436
rect -1986 -5412 -1952 -3436
rect -1868 -5412 -1834 -3436
rect -1750 -5412 -1716 -3436
rect -1632 -5412 -1598 -3436
rect -1175 -4088 -1141 -3612
rect -1079 -4088 -1045 -3612
rect -983 -4088 -949 -3612
rect -887 -4088 -853 -3612
rect -791 -4088 -757 -3612
rect -695 -4088 -661 -3612
rect -599 -4088 -565 -3612
rect -503 -4088 -469 -3612
rect -407 -4088 -373 -3612
rect -311 -4088 -277 -3612
rect -215 -4088 -181 -3612
rect -119 -4088 -85 -3612
rect -23 -4088 11 -3612
rect 73 -4088 107 -3612
rect 169 -4088 203 -3612
rect 265 -4088 299 -3612
rect 361 -4088 395 -3612
rect 457 -4088 491 -3612
rect 553 -4088 587 -3612
rect 649 -4088 683 -3612
rect 745 -4088 779 -3612
rect -3538 -5932 -3062 -5898
rect -3538 -6028 -3062 -5994
rect -3538 -6124 -3062 -6090
rect -3538 -6220 -3062 -6186
rect -3538 -6316 -3062 -6282
rect -1131 -6528 -1097 -4552
rect -673 -6528 -639 -4552
rect -215 -6528 -181 -4552
rect 243 -6528 277 -4552
rect 701 -6528 735 -4552
rect 1201 -5412 1235 -3436
rect 1319 -5412 1353 -3436
rect 1437 -5412 1471 -3436
rect 1555 -5412 1589 -3436
rect 1673 -5412 1707 -3436
rect 1791 -5412 1825 -3436
rect 1909 -5412 1943 -3436
<< pdiffc >>
rect -2103 -2903 -2069 -927
rect -1985 -2903 -1951 -927
rect -1867 -2903 -1833 -927
rect -1749 -2903 -1715 -927
rect -1631 -2903 -1597 -927
rect -1513 -2903 -1479 -927
rect -1395 -2903 -1361 -927
rect -1277 -2903 -1243 -927
rect -1159 -2903 -1125 -927
rect -1041 -2903 -1007 -927
rect -923 -2903 -889 -927
rect -805 -2903 -771 -927
rect -687 -2903 -653 -927
rect -569 -2903 -535 -927
rect -451 -2903 -417 -927
rect -333 -2903 -299 -927
rect -215 -2903 -181 -927
rect -97 -2903 -63 -927
rect 21 -2903 55 -927
rect 139 -2903 173 -927
rect 257 -2903 291 -927
rect 375 -2903 409 -927
rect 493 -2903 527 -927
rect 611 -2903 645 -927
rect 729 -2903 763 -927
rect 847 -2903 881 -927
rect 965 -2903 999 -927
rect 1083 -2903 1117 -927
rect 1201 -2903 1235 -927
rect 1319 -2903 1353 -927
rect 1437 -2903 1471 -927
rect 1555 -2903 1589 -927
rect 1673 -2903 1707 -927
<< psubdiff >>
rect -2454 -3284 -2358 -3250
rect -1580 -3284 -1484 -3250
rect -2454 -3346 -2420 -3284
rect -1518 -3346 -1484 -3284
rect -2454 -5564 -2420 -5502
rect 1087 -3284 1183 -3250
rect 1961 -3284 2057 -3250
rect 1087 -3346 1121 -3284
rect -1289 -3460 -1193 -3426
rect 797 -3460 893 -3426
rect -1289 -3522 -1255 -3460
rect 859 -3522 893 -3460
rect -1289 -4240 -1255 -4178
rect 859 -4240 893 -4178
rect -1289 -4274 -1193 -4240
rect 797 -4274 893 -4240
rect -1518 -5564 -1484 -5502
rect -2454 -5598 -2358 -5564
rect -1580 -5598 -1484 -5564
rect -1245 -4400 -1149 -4366
rect 753 -4400 849 -4366
rect -1245 -4462 -1211 -4400
rect -3724 -5818 -3628 -5784
rect -2972 -5818 -2876 -5784
rect -3724 -5880 -3690 -5818
rect -2910 -5880 -2876 -5818
rect -3724 -6812 -3690 -6730
rect 815 -4462 849 -4400
rect -1245 -6680 -1211 -6618
rect 2023 -3346 2057 -3284
rect 1087 -5564 1121 -5502
rect 2128 -3652 2224 -3618
rect 2664 -3652 2760 -3618
rect 2128 -3714 2162 -3652
rect 2726 -3714 2760 -3652
rect 2128 -4880 2162 -4818
rect 2726 -4880 2760 -4818
rect 2128 -4914 2224 -4880
rect 2664 -4914 2760 -4880
rect 2023 -5564 2057 -5502
rect 1087 -5598 1183 -5564
rect 1961 -5598 2057 -5564
rect 815 -6680 849 -6618
rect -1245 -6714 -1149 -6680
rect 753 -6714 849 -6680
rect -2910 -6812 -2876 -6730
rect -3724 -6846 -3628 -6812
rect -2972 -6846 -2876 -6812
<< nsubdiff >>
rect -2217 -766 -2121 -732
rect 1725 -766 1821 -732
rect -2217 -828 -2183 -766
rect 1787 -828 1821 -766
rect -2217 -3064 -2183 -3002
rect 1787 -3064 1821 -3002
rect -2217 -3098 -2121 -3064
rect 1725 -3098 1821 -3064
<< psubdiffcont >>
rect -2358 -3284 -1580 -3250
rect -2454 -5502 -2420 -3346
rect -1518 -5502 -1484 -3346
rect 1183 -3284 1961 -3250
rect -1193 -3460 797 -3426
rect -1289 -4178 -1255 -3522
rect 859 -4178 893 -3522
rect -1193 -4274 797 -4240
rect -2358 -5598 -1580 -5564
rect -1149 -4400 753 -4366
rect -3628 -5818 -2972 -5784
rect -3724 -6730 -3690 -5880
rect -2910 -6730 -2876 -5880
rect -1245 -6618 -1211 -4462
rect 815 -6618 849 -4462
rect 1087 -5502 1121 -3346
rect 2023 -5502 2057 -3346
rect 2224 -3652 2664 -3618
rect 2128 -4818 2162 -3714
rect 2726 -4818 2760 -3714
rect 2224 -4914 2664 -4880
rect 1183 -5598 1961 -5564
rect -1149 -6714 753 -6680
rect -3628 -6846 -2972 -6812
<< nsubdiffcont >>
rect -2121 -766 1725 -732
rect -2217 -3002 -2183 -828
rect 1787 -3002 1821 -828
rect -2121 -3098 1725 -3064
<< poly >>
rect -2060 -834 -1994 -818
rect -2060 -868 -2044 -834
rect -2010 -868 -1994 -834
rect -2060 -884 -1994 -868
rect -1942 -834 -1876 -818
rect -1942 -868 -1926 -834
rect -1892 -868 -1876 -834
rect -1942 -884 -1876 -868
rect -1824 -834 -1758 -818
rect -1824 -868 -1808 -834
rect -1774 -868 -1758 -834
rect -1824 -884 -1758 -868
rect -1706 -834 -1640 -818
rect -1706 -868 -1690 -834
rect -1656 -868 -1640 -834
rect -1706 -884 -1640 -868
rect -1588 -834 -1522 -818
rect -1588 -868 -1572 -834
rect -1538 -868 -1522 -834
rect -1588 -884 -1522 -868
rect -1470 -834 -1404 -818
rect -1470 -868 -1454 -834
rect -1420 -868 -1404 -834
rect -1470 -884 -1404 -868
rect -1352 -834 -1286 -818
rect -1352 -868 -1336 -834
rect -1302 -868 -1286 -834
rect -1352 -884 -1286 -868
rect -1234 -834 -1168 -818
rect -1234 -868 -1218 -834
rect -1184 -868 -1168 -834
rect -1234 -884 -1168 -868
rect -1116 -834 -1050 -818
rect -1116 -868 -1100 -834
rect -1066 -868 -1050 -834
rect -1116 -884 -1050 -868
rect -998 -834 -932 -818
rect -998 -868 -982 -834
rect -948 -868 -932 -834
rect -998 -884 -932 -868
rect -880 -834 -814 -818
rect -880 -868 -864 -834
rect -830 -868 -814 -834
rect -880 -884 -814 -868
rect -762 -834 -696 -818
rect -762 -868 -746 -834
rect -712 -868 -696 -834
rect -762 -884 -696 -868
rect -644 -884 -578 -818
rect -526 -884 -460 -818
rect -408 -884 -342 -818
rect -290 -884 -224 -818
rect -172 -884 -106 -818
rect -54 -884 12 -818
rect 64 -884 130 -818
rect 182 -884 248 -818
rect 300 -834 366 -818
rect 300 -868 316 -834
rect 350 -868 366 -834
rect 300 -884 366 -868
rect 418 -834 484 -818
rect 418 -868 434 -834
rect 468 -868 484 -834
rect 418 -884 484 -868
rect 536 -834 602 -818
rect 536 -868 552 -834
rect 586 -868 602 -834
rect 536 -884 602 -868
rect 654 -834 720 -818
rect 654 -868 670 -834
rect 704 -868 720 -834
rect 654 -884 720 -868
rect 772 -834 838 -818
rect 772 -868 788 -834
rect 822 -868 838 -834
rect 772 -884 838 -868
rect 890 -834 956 -818
rect 890 -868 906 -834
rect 940 -868 956 -834
rect 890 -884 956 -868
rect 1008 -834 1074 -818
rect 1008 -868 1024 -834
rect 1058 -868 1074 -834
rect 1008 -884 1074 -868
rect 1126 -834 1192 -818
rect 1126 -868 1142 -834
rect 1176 -868 1192 -834
rect 1126 -884 1192 -868
rect 1244 -834 1310 -818
rect 1244 -868 1260 -834
rect 1294 -868 1310 -834
rect 1244 -884 1310 -868
rect 1362 -834 1428 -818
rect 1362 -868 1378 -834
rect 1412 -868 1428 -834
rect 1362 -884 1428 -868
rect 1480 -834 1546 -818
rect 1480 -868 1496 -834
rect 1530 -868 1546 -834
rect 1480 -884 1546 -868
rect 1598 -834 1664 -818
rect 1598 -868 1614 -834
rect 1648 -868 1664 -834
rect 1598 -884 1664 -868
rect -2057 -915 -1997 -884
rect -1939 -915 -1879 -884
rect -1821 -915 -1761 -884
rect -1703 -915 -1643 -884
rect -1585 -915 -1525 -884
rect -1467 -915 -1407 -884
rect -1349 -915 -1289 -884
rect -1231 -915 -1171 -884
rect -1113 -915 -1053 -884
rect -995 -915 -935 -884
rect -877 -915 -817 -884
rect -759 -915 -699 -884
rect -641 -915 -581 -884
rect -523 -915 -463 -884
rect -405 -915 -345 -884
rect -287 -915 -227 -884
rect -169 -915 -109 -884
rect -51 -915 9 -884
rect 67 -915 127 -884
rect 185 -915 245 -884
rect 303 -915 363 -884
rect 421 -915 481 -884
rect 539 -915 599 -884
rect 657 -915 717 -884
rect 775 -915 835 -884
rect 893 -915 953 -884
rect 1011 -915 1071 -884
rect 1129 -915 1189 -884
rect 1247 -915 1307 -884
rect 1365 -915 1425 -884
rect 1483 -915 1543 -884
rect 1601 -915 1661 -884
rect -2057 -2946 -1997 -2915
rect -1939 -2946 -1879 -2915
rect -1821 -2946 -1761 -2915
rect -1703 -2946 -1643 -2915
rect -1585 -2946 -1525 -2915
rect -1467 -2946 -1407 -2915
rect -1349 -2946 -1289 -2915
rect -1231 -2946 -1171 -2915
rect -1113 -2946 -1053 -2915
rect -995 -2946 -935 -2915
rect -877 -2946 -817 -2915
rect -759 -2946 -699 -2915
rect -641 -2946 -581 -2915
rect -523 -2946 -463 -2915
rect -405 -2946 -345 -2915
rect -287 -2946 -227 -2915
rect -169 -2946 -109 -2915
rect -51 -2946 9 -2915
rect 67 -2946 127 -2915
rect 185 -2946 245 -2915
rect 303 -2946 363 -2915
rect 421 -2946 481 -2915
rect 539 -2946 599 -2915
rect 657 -2946 717 -2915
rect 775 -2946 835 -2915
rect 893 -2946 953 -2915
rect 1011 -2946 1071 -2915
rect 1129 -2946 1189 -2915
rect 1247 -2946 1307 -2915
rect 1365 -2946 1425 -2915
rect 1483 -2946 1543 -2915
rect 1601 -2946 1661 -2915
rect -2060 -2962 -1994 -2946
rect -2060 -2996 -2044 -2962
rect -2010 -2996 -1994 -2962
rect -2060 -3012 -1994 -2996
rect -1942 -2962 -1876 -2946
rect -1942 -2996 -1926 -2962
rect -1892 -2996 -1876 -2962
rect -1942 -3012 -1876 -2996
rect -1824 -2962 -1758 -2946
rect -1824 -2996 -1808 -2962
rect -1774 -2996 -1758 -2962
rect -1824 -3012 -1758 -2996
rect -1706 -2962 -1640 -2946
rect -1706 -2996 -1690 -2962
rect -1656 -2996 -1640 -2962
rect -1706 -3012 -1640 -2996
rect -1588 -2962 -1522 -2946
rect -1588 -2996 -1572 -2962
rect -1538 -2996 -1522 -2962
rect -1588 -3012 -1522 -2996
rect -1470 -2962 -1404 -2946
rect -1470 -2996 -1454 -2962
rect -1420 -2996 -1404 -2962
rect -1470 -3012 -1404 -2996
rect -1352 -2962 -1286 -2946
rect -1352 -2996 -1336 -2962
rect -1302 -2996 -1286 -2962
rect -1352 -3012 -1286 -2996
rect -1234 -2962 -1168 -2946
rect -1234 -2996 -1218 -2962
rect -1184 -2996 -1168 -2962
rect -1234 -3012 -1168 -2996
rect -1116 -2962 -1050 -2946
rect -1116 -2996 -1100 -2962
rect -1066 -2996 -1050 -2962
rect -1116 -3012 -1050 -2996
rect -998 -2962 -932 -2946
rect -998 -2996 -982 -2962
rect -948 -2996 -932 -2962
rect -998 -3012 -932 -2996
rect -880 -2962 -814 -2946
rect -880 -2996 -864 -2962
rect -830 -2996 -814 -2962
rect -880 -3012 -814 -2996
rect -762 -2962 -696 -2946
rect -762 -2996 -746 -2962
rect -712 -2996 -696 -2962
rect -762 -3012 -696 -2996
rect -644 -2962 -578 -2946
rect -644 -2996 -628 -2962
rect -594 -2996 -578 -2962
rect -644 -3012 -578 -2996
rect -526 -2962 -460 -2946
rect -526 -2996 -510 -2962
rect -476 -2996 -460 -2962
rect -526 -3012 -460 -2996
rect -408 -2962 -342 -2946
rect -408 -2996 -392 -2962
rect -358 -2996 -342 -2962
rect -408 -3012 -342 -2996
rect -290 -2962 -224 -2946
rect -290 -2996 -274 -2962
rect -240 -2996 -224 -2962
rect -290 -3012 -224 -2996
rect -172 -2962 -106 -2946
rect -172 -2996 -156 -2962
rect -122 -2996 -106 -2962
rect -172 -3012 -106 -2996
rect -54 -2962 12 -2946
rect -54 -2996 -38 -2962
rect -4 -2996 12 -2962
rect -54 -3012 12 -2996
rect 64 -2962 130 -2946
rect 64 -2996 80 -2962
rect 114 -2996 130 -2962
rect 64 -3012 130 -2996
rect 182 -2962 248 -2946
rect 182 -2996 198 -2962
rect 232 -2996 248 -2962
rect 182 -3012 248 -2996
rect 300 -2962 366 -2946
rect 300 -2996 316 -2962
rect 350 -2996 366 -2962
rect 300 -3012 366 -2996
rect 418 -2962 484 -2946
rect 418 -2996 434 -2962
rect 468 -2996 484 -2962
rect 418 -3012 484 -2996
rect 536 -2962 602 -2946
rect 536 -2996 552 -2962
rect 586 -2996 602 -2962
rect 536 -3012 602 -2996
rect 654 -2962 720 -2946
rect 654 -2996 670 -2962
rect 704 -2996 720 -2962
rect 654 -3012 720 -2996
rect 772 -2962 838 -2946
rect 772 -2996 788 -2962
rect 822 -2996 838 -2962
rect 772 -3012 838 -2996
rect 890 -2962 956 -2946
rect 890 -2996 906 -2962
rect 940 -2996 956 -2962
rect 890 -3012 956 -2996
rect 1008 -2962 1074 -2946
rect 1008 -2996 1024 -2962
rect 1058 -2996 1074 -2962
rect 1008 -3012 1074 -2996
rect 1126 -2962 1192 -2946
rect 1126 -2996 1142 -2962
rect 1176 -2996 1192 -2962
rect 1126 -3012 1192 -2996
rect 1244 -2962 1310 -2946
rect 1244 -2996 1260 -2962
rect 1294 -2996 1310 -2962
rect 1244 -3012 1310 -2996
rect 1362 -2962 1428 -2946
rect 1362 -2996 1378 -2962
rect 1412 -2996 1428 -2962
rect 1362 -3012 1428 -2996
rect 1480 -2962 1546 -2946
rect 1480 -2996 1496 -2962
rect 1530 -2996 1546 -2962
rect 1480 -3012 1546 -2996
rect 1598 -2962 1664 -2946
rect 1598 -2996 1614 -2962
rect 1648 -2996 1664 -2962
rect 1598 -3012 1664 -2996
rect -2297 -3352 -2231 -3336
rect -2297 -3386 -2281 -3352
rect -2247 -3386 -2231 -3352
rect -2297 -3402 -2231 -3386
rect -2179 -3352 -2113 -3336
rect -2179 -3386 -2163 -3352
rect -2129 -3386 -2113 -3352
rect -2179 -3402 -2113 -3386
rect -2061 -3352 -1995 -3336
rect -2061 -3386 -2045 -3352
rect -2011 -3386 -1995 -3352
rect -2061 -3402 -1995 -3386
rect -1943 -3352 -1877 -3336
rect -1943 -3386 -1927 -3352
rect -1893 -3386 -1877 -3352
rect -1943 -3402 -1877 -3386
rect -1825 -3352 -1759 -3336
rect -1825 -3386 -1809 -3352
rect -1775 -3386 -1759 -3352
rect -1825 -3402 -1759 -3386
rect -1707 -3352 -1641 -3336
rect -1707 -3386 -1691 -3352
rect -1657 -3386 -1641 -3352
rect -1707 -3402 -1641 -3386
rect -2294 -3424 -2234 -3402
rect -2176 -3424 -2116 -3402
rect -2058 -3424 -1998 -3402
rect -1940 -3424 -1880 -3402
rect -1822 -3424 -1762 -3402
rect -1704 -3424 -1644 -3402
rect -2294 -5446 -2234 -5424
rect -2176 -5446 -2116 -5424
rect -2058 -5446 -1998 -5424
rect -1940 -5446 -1880 -5424
rect -1822 -5446 -1762 -5424
rect -1704 -5446 -1644 -5424
rect -2297 -5462 -2231 -5446
rect -2297 -5496 -2281 -5462
rect -2247 -5496 -2231 -5462
rect -2297 -5512 -2231 -5496
rect -2179 -5462 -2113 -5446
rect -2179 -5496 -2163 -5462
rect -2129 -5496 -2113 -5462
rect -2179 -5512 -2113 -5496
rect -2061 -5462 -1995 -5446
rect -2061 -5496 -2045 -5462
rect -2011 -5496 -1995 -5462
rect -2061 -5512 -1995 -5496
rect -1943 -5462 -1877 -5446
rect -1943 -5496 -1927 -5462
rect -1893 -5496 -1877 -5462
rect -1943 -5512 -1877 -5496
rect -1825 -5462 -1759 -5446
rect -1825 -5496 -1809 -5462
rect -1775 -5496 -1759 -5462
rect -1825 -5512 -1759 -5496
rect -1707 -5462 -1641 -5446
rect -1707 -5496 -1691 -5462
rect -1657 -5496 -1641 -5462
rect -1707 -5512 -1641 -5496
rect -1125 -3524 -999 -3496
rect -1125 -3558 -1079 -3524
rect -1045 -3558 -999 -3524
rect -1125 -3574 -999 -3558
rect 603 -3524 729 -3496
rect 603 -3558 649 -3524
rect 683 -3558 729 -3524
rect 603 -3574 729 -3558
rect -1125 -3600 -1095 -3574
rect -1029 -3600 -999 -3574
rect -933 -3600 -903 -3574
rect -837 -3600 -807 -3574
rect -741 -3600 -711 -3574
rect -645 -3600 -615 -3574
rect -549 -3600 -519 -3574
rect -453 -3600 -423 -3574
rect -357 -3600 -327 -3574
rect -261 -3600 -231 -3574
rect -165 -3600 -135 -3574
rect -69 -3600 -39 -3574
rect 27 -3600 57 -3574
rect 123 -3600 153 -3574
rect 219 -3600 249 -3574
rect 315 -3600 345 -3574
rect 411 -3600 441 -3574
rect 507 -3600 537 -3574
rect 603 -3600 633 -3574
rect 699 -3600 729 -3574
rect -1125 -4126 -1095 -4100
rect -1029 -4126 -999 -4100
rect -933 -4122 -903 -4100
rect -837 -4122 -807 -4100
rect -933 -4150 -807 -4122
rect -933 -4184 -887 -4150
rect -853 -4184 -807 -4150
rect -933 -4200 -807 -4184
rect -741 -4122 -711 -4100
rect -645 -4122 -615 -4100
rect -741 -4150 -615 -4122
rect -741 -4184 -695 -4150
rect -661 -4184 -615 -4150
rect -741 -4200 -615 -4184
rect -549 -4122 -519 -4100
rect -453 -4122 -423 -4100
rect -549 -4150 -423 -4122
rect -549 -4184 -503 -4150
rect -469 -4184 -423 -4150
rect -549 -4200 -423 -4184
rect -357 -4122 -327 -4100
rect -261 -4122 -231 -4100
rect -357 -4150 -231 -4122
rect -357 -4184 -311 -4150
rect -277 -4184 -231 -4150
rect -357 -4200 -231 -4184
rect -165 -4122 -135 -4100
rect -69 -4122 -39 -4100
rect -165 -4150 -39 -4122
rect -165 -4184 -119 -4150
rect -85 -4184 -39 -4150
rect -165 -4200 -39 -4184
rect 27 -4122 57 -4100
rect 123 -4122 153 -4100
rect 27 -4150 153 -4122
rect 27 -4184 73 -4150
rect 107 -4184 153 -4150
rect 27 -4200 153 -4184
rect 219 -4122 249 -4100
rect 315 -4122 345 -4100
rect 219 -4150 345 -4122
rect 219 -4184 265 -4150
rect 299 -4184 345 -4150
rect 219 -4200 345 -4184
rect 411 -4122 441 -4100
rect 507 -4122 537 -4100
rect 411 -4150 537 -4122
rect 603 -4126 633 -4100
rect 699 -4126 729 -4100
rect 411 -4184 457 -4150
rect 491 -4184 537 -4150
rect 411 -4200 537 -4184
rect -3638 -5964 -3550 -5948
rect -3638 -5998 -3622 -5964
rect -3588 -5978 -3550 -5964
rect -3050 -5978 -3024 -5948
rect -3588 -5998 -3572 -5978
rect -3638 -6044 -3572 -5998
rect -3638 -6074 -3550 -6044
rect -3050 -6074 -3024 -6044
rect -3638 -6156 -3550 -6140
rect -3638 -6190 -3622 -6156
rect -3588 -6170 -3550 -6156
rect -3050 -6170 -3024 -6140
rect -3588 -6190 -3572 -6170
rect -3638 -6236 -3572 -6190
rect -3638 -6266 -3550 -6236
rect -3050 -6266 -3024 -6236
rect -1085 -4468 -685 -4452
rect -1085 -4502 -1069 -4468
rect -701 -4502 -685 -4468
rect -1085 -4540 -685 -4502
rect -627 -4468 -227 -4452
rect -627 -4502 -611 -4468
rect -243 -4502 -227 -4468
rect -627 -4540 -227 -4502
rect -169 -4468 231 -4452
rect -169 -4502 -153 -4468
rect 215 -4502 231 -4468
rect -169 -4540 231 -4502
rect 289 -4468 689 -4452
rect 289 -4502 305 -4468
rect 673 -4502 689 -4468
rect 289 -4540 689 -4502
rect -1085 -6578 -685 -6540
rect -1085 -6612 -1069 -6578
rect -701 -6612 -685 -6578
rect -1085 -6628 -685 -6612
rect -627 -6578 -227 -6540
rect -627 -6612 -611 -6578
rect -243 -6612 -227 -6578
rect -627 -6628 -227 -6612
rect -169 -6578 231 -6540
rect -169 -6612 -153 -6578
rect 215 -6612 231 -6578
rect -169 -6628 231 -6612
rect 289 -6578 689 -6540
rect 289 -6612 305 -6578
rect 673 -6612 689 -6578
rect 289 -6628 689 -6612
rect 1244 -3352 1310 -3336
rect 1244 -3386 1260 -3352
rect 1294 -3386 1310 -3352
rect 1244 -3402 1310 -3386
rect 1362 -3352 1428 -3336
rect 1362 -3386 1378 -3352
rect 1412 -3386 1428 -3352
rect 1362 -3402 1428 -3386
rect 1480 -3352 1546 -3336
rect 1480 -3386 1496 -3352
rect 1530 -3386 1546 -3352
rect 1480 -3402 1546 -3386
rect 1598 -3352 1664 -3336
rect 1598 -3386 1614 -3352
rect 1648 -3386 1664 -3352
rect 1598 -3402 1664 -3386
rect 1716 -3352 1782 -3336
rect 1716 -3386 1732 -3352
rect 1766 -3386 1782 -3352
rect 1716 -3402 1782 -3386
rect 1834 -3352 1900 -3336
rect 1834 -3386 1850 -3352
rect 1884 -3386 1900 -3352
rect 1834 -3402 1900 -3386
rect 1247 -3424 1307 -3402
rect 1365 -3424 1425 -3402
rect 1483 -3424 1543 -3402
rect 1601 -3424 1661 -3402
rect 1719 -3424 1779 -3402
rect 1837 -3424 1897 -3402
rect 1247 -5446 1307 -5424
rect 1365 -5446 1425 -5424
rect 1483 -5446 1543 -5424
rect 1601 -5446 1661 -5424
rect 1719 -5446 1779 -5424
rect 1837 -5446 1897 -5424
rect 1244 -5462 1310 -5446
rect 1244 -5496 1260 -5462
rect 1294 -5496 1310 -5462
rect 1244 -5512 1310 -5496
rect 1362 -5462 1428 -5446
rect 1362 -5496 1378 -5462
rect 1412 -5496 1428 -5462
rect 1362 -5512 1428 -5496
rect 1480 -5462 1546 -5446
rect 1480 -5496 1496 -5462
rect 1530 -5496 1546 -5462
rect 1480 -5512 1546 -5496
rect 1598 -5462 1664 -5446
rect 1598 -5496 1614 -5462
rect 1648 -5496 1664 -5462
rect 1598 -5512 1664 -5496
rect 1716 -5462 1782 -5446
rect 1716 -5496 1732 -5462
rect 1766 -5496 1782 -5462
rect 1716 -5512 1782 -5496
rect 1834 -5462 1900 -5446
rect 1834 -5496 1850 -5462
rect 1884 -5496 1900 -5462
rect 1834 -5512 1900 -5496
<< polycont >>
rect -2044 -868 -2010 -834
rect -1926 -868 -1892 -834
rect -1808 -868 -1774 -834
rect -1690 -868 -1656 -834
rect -1572 -868 -1538 -834
rect -1454 -868 -1420 -834
rect -1336 -868 -1302 -834
rect -1218 -868 -1184 -834
rect -1100 -868 -1066 -834
rect -982 -868 -948 -834
rect -864 -868 -830 -834
rect -746 -868 -712 -834
rect 316 -868 350 -834
rect 434 -868 468 -834
rect 552 -868 586 -834
rect 670 -868 704 -834
rect 788 -868 822 -834
rect 906 -868 940 -834
rect 1024 -868 1058 -834
rect 1142 -868 1176 -834
rect 1260 -868 1294 -834
rect 1378 -868 1412 -834
rect 1496 -868 1530 -834
rect 1614 -868 1648 -834
rect -2044 -2996 -2010 -2962
rect -1926 -2996 -1892 -2962
rect -1808 -2996 -1774 -2962
rect -1690 -2996 -1656 -2962
rect -1572 -2996 -1538 -2962
rect -1454 -2996 -1420 -2962
rect -1336 -2996 -1302 -2962
rect -1218 -2996 -1184 -2962
rect -1100 -2996 -1066 -2962
rect -982 -2996 -948 -2962
rect -864 -2996 -830 -2962
rect -746 -2996 -712 -2962
rect -628 -2996 -594 -2962
rect -510 -2996 -476 -2962
rect -392 -2996 -358 -2962
rect -274 -2996 -240 -2962
rect -156 -2996 -122 -2962
rect -38 -2996 -4 -2962
rect 80 -2996 114 -2962
rect 198 -2996 232 -2962
rect 316 -2996 350 -2962
rect 434 -2996 468 -2962
rect 552 -2996 586 -2962
rect 670 -2996 704 -2962
rect 788 -2996 822 -2962
rect 906 -2996 940 -2962
rect 1024 -2996 1058 -2962
rect 1142 -2996 1176 -2962
rect 1260 -2996 1294 -2962
rect 1378 -2996 1412 -2962
rect 1496 -2996 1530 -2962
rect 1614 -2996 1648 -2962
rect -2281 -3386 -2247 -3352
rect -2163 -3386 -2129 -3352
rect -2045 -3386 -2011 -3352
rect -1927 -3386 -1893 -3352
rect -1809 -3386 -1775 -3352
rect -1691 -3386 -1657 -3352
rect -2281 -5496 -2247 -5462
rect -2163 -5496 -2129 -5462
rect -2045 -5496 -2011 -5462
rect -1927 -5496 -1893 -5462
rect -1809 -5496 -1775 -5462
rect -1691 -5496 -1657 -5462
rect -1079 -3558 -1045 -3524
rect 649 -3558 683 -3524
rect -887 -4184 -853 -4150
rect -695 -4184 -661 -4150
rect -503 -4184 -469 -4150
rect -311 -4184 -277 -4150
rect -119 -4184 -85 -4150
rect 73 -4184 107 -4150
rect 265 -4184 299 -4150
rect 457 -4184 491 -4150
rect -3622 -5998 -3588 -5964
rect -3622 -6190 -3588 -6156
rect -1069 -4502 -701 -4468
rect -611 -4502 -243 -4468
rect -153 -4502 215 -4468
rect 305 -4502 673 -4468
rect -1069 -6612 -701 -6578
rect -611 -6612 -243 -6578
rect -153 -6612 215 -6578
rect 305 -6612 673 -6578
rect 1260 -3386 1294 -3352
rect 1378 -3386 1412 -3352
rect 1496 -3386 1530 -3352
rect 1614 -3386 1648 -3352
rect 1732 -3386 1766 -3352
rect 1850 -3386 1884 -3352
rect 1260 -5496 1294 -5462
rect 1378 -5496 1412 -5462
rect 1496 -5496 1530 -5462
rect 1614 -5496 1648 -5462
rect 1732 -5496 1766 -5462
rect 1850 -5496 1884 -5462
<< xpolycontact >>
rect -3594 -6504 -3162 -6434
rect -3594 -6670 -3162 -6600
rect 2258 -4180 2396 -3748
rect 2492 -4180 2630 -3748
<< ppolyres >>
rect 2258 -4646 2396 -4180
rect 2492 -4646 2630 -4180
rect 2258 -4784 2630 -4646
<< xpolyres >>
rect -3162 -6504 -3026 -6434
rect -3096 -6600 -3026 -6504
rect -3162 -6670 -3026 -6600
<< locali >>
rect -2217 -766 -2121 -732
rect 1725 -766 1821 -732
rect -2217 -828 -2183 -766
rect 1787 -828 1821 -766
rect -2060 -868 -2044 -834
rect -2010 -868 -1994 -834
rect -1942 -868 -1926 -834
rect -1892 -868 -1876 -834
rect -1824 -868 -1808 -834
rect -1774 -868 -1758 -834
rect -1706 -868 -1690 -834
rect -1656 -868 -1640 -834
rect -1588 -868 -1572 -834
rect -1538 -868 -1522 -834
rect -1470 -868 -1454 -834
rect -1420 -868 -1404 -834
rect -1352 -868 -1336 -834
rect -1302 -868 -1286 -834
rect -1234 -868 -1218 -834
rect -1184 -868 -1168 -834
rect -1116 -868 -1100 -834
rect -1066 -868 -1050 -834
rect -998 -868 -982 -834
rect -948 -868 -932 -834
rect -880 -868 -864 -834
rect -830 -868 -814 -834
rect -762 -868 -746 -834
rect -712 -868 -696 -834
rect 300 -868 316 -834
rect 350 -868 366 -834
rect 418 -868 434 -834
rect 468 -868 484 -834
rect 536 -868 552 -834
rect 586 -868 602 -834
rect 654 -868 670 -834
rect 704 -868 720 -834
rect 772 -868 788 -834
rect 822 -868 838 -834
rect 890 -868 906 -834
rect 940 -868 956 -834
rect 1008 -868 1024 -834
rect 1058 -868 1074 -834
rect 1126 -868 1142 -834
rect 1176 -868 1192 -834
rect 1244 -868 1260 -834
rect 1294 -868 1310 -834
rect 1362 -868 1378 -834
rect 1412 -868 1428 -834
rect 1480 -868 1496 -834
rect 1530 -868 1546 -834
rect 1598 -868 1614 -834
rect 1648 -868 1664 -834
rect -2103 -927 -2069 -911
rect -2103 -2919 -2069 -2903
rect -1985 -927 -1951 -911
rect -1985 -2919 -1951 -2903
rect -1867 -927 -1833 -911
rect -1867 -2919 -1833 -2903
rect -1749 -927 -1715 -911
rect -1749 -2919 -1715 -2903
rect -1631 -927 -1597 -911
rect -1631 -2919 -1597 -2903
rect -1513 -927 -1479 -911
rect -1513 -2919 -1479 -2903
rect -1395 -927 -1361 -911
rect -1395 -2919 -1361 -2903
rect -1277 -927 -1243 -911
rect -1277 -2919 -1243 -2903
rect -1159 -927 -1125 -911
rect -1159 -2919 -1125 -2903
rect -1041 -927 -1007 -911
rect -1041 -2919 -1007 -2903
rect -923 -927 -889 -911
rect -923 -2919 -889 -2903
rect -805 -927 -771 -911
rect -805 -2919 -771 -2903
rect -687 -927 -653 -911
rect -687 -2919 -653 -2903
rect -569 -927 -535 -911
rect -569 -2919 -535 -2903
rect -451 -927 -417 -911
rect -451 -2919 -417 -2903
rect -333 -927 -299 -911
rect -333 -2919 -299 -2903
rect -215 -927 -181 -911
rect -215 -2919 -181 -2903
rect -97 -927 -63 -911
rect -97 -2919 -63 -2903
rect 21 -927 55 -911
rect 21 -2919 55 -2903
rect 139 -927 173 -911
rect 139 -2919 173 -2903
rect 257 -927 291 -911
rect 257 -2919 291 -2903
rect 375 -927 409 -911
rect 375 -2919 409 -2903
rect 493 -927 527 -911
rect 493 -2919 527 -2903
rect 611 -927 645 -911
rect 611 -2919 645 -2903
rect 729 -927 763 -911
rect 729 -2919 763 -2903
rect 847 -927 881 -911
rect 847 -2919 881 -2903
rect 965 -927 999 -911
rect 965 -2919 999 -2903
rect 1083 -927 1117 -911
rect 1083 -2919 1117 -2903
rect 1201 -927 1235 -911
rect 1201 -2919 1235 -2903
rect 1319 -927 1353 -911
rect 1319 -2919 1353 -2903
rect 1437 -927 1471 -911
rect 1437 -2919 1471 -2903
rect 1555 -927 1589 -911
rect 1555 -2919 1589 -2903
rect 1673 -927 1707 -911
rect 1673 -2919 1707 -2903
rect -2060 -2996 -2044 -2962
rect -2010 -2996 -1994 -2962
rect -1942 -2996 -1926 -2962
rect -1892 -2996 -1876 -2962
rect -1824 -2996 -1808 -2962
rect -1774 -2996 -1758 -2962
rect -1706 -2996 -1690 -2962
rect -1656 -2996 -1640 -2962
rect -1588 -2996 -1572 -2962
rect -1538 -2996 -1522 -2962
rect -1470 -2996 -1454 -2962
rect -1420 -2996 -1404 -2962
rect -1352 -2996 -1336 -2962
rect -1302 -2996 -1286 -2962
rect -1234 -2996 -1218 -2962
rect -1184 -2996 -1168 -2962
rect -1116 -2996 -1100 -2962
rect -1066 -2996 -1050 -2962
rect -998 -2996 -982 -2962
rect -948 -2996 -932 -2962
rect -880 -2996 -864 -2962
rect -830 -2996 -814 -2962
rect -762 -2996 -746 -2962
rect -712 -2996 -696 -2962
rect -644 -2996 -628 -2962
rect -594 -2996 -578 -2962
rect -526 -2996 -510 -2962
rect -476 -2996 -460 -2962
rect -408 -2996 -392 -2962
rect -358 -2996 -342 -2962
rect -290 -2996 -274 -2962
rect -240 -2996 -224 -2962
rect -172 -2996 -156 -2962
rect -122 -2996 -106 -2962
rect -54 -2996 -38 -2962
rect -4 -2996 12 -2962
rect 64 -2996 80 -2962
rect 114 -2996 130 -2962
rect 182 -2996 198 -2962
rect 232 -2996 248 -2962
rect 300 -2996 316 -2962
rect 350 -2996 366 -2962
rect 418 -2996 434 -2962
rect 468 -2996 484 -2962
rect 536 -2996 552 -2962
rect 586 -2996 602 -2962
rect 654 -2996 670 -2962
rect 704 -2996 720 -2962
rect 772 -2996 788 -2962
rect 822 -2996 838 -2962
rect 890 -2996 906 -2962
rect 940 -2996 956 -2962
rect 1008 -2996 1024 -2962
rect 1058 -2996 1074 -2962
rect 1126 -2996 1142 -2962
rect 1176 -2996 1192 -2962
rect 1244 -2996 1260 -2962
rect 1294 -2996 1310 -2962
rect 1362 -2996 1378 -2962
rect 1412 -2996 1428 -2962
rect 1480 -2996 1496 -2962
rect 1530 -2996 1546 -2962
rect 1598 -2996 1614 -2962
rect 1648 -2996 1664 -2962
rect -2217 -3064 -2183 -3002
rect 1787 -3064 1821 -3002
rect -2217 -3098 -2121 -3064
rect 1725 -3098 1821 -3064
rect -2454 -3284 -2358 -3250
rect -1580 -3284 -1484 -3250
rect -2454 -3346 -2420 -3284
rect -1518 -3346 -1484 -3284
rect -2297 -3386 -2281 -3352
rect -2247 -3386 -2231 -3352
rect -2179 -3386 -2163 -3352
rect -2129 -3386 -2113 -3352
rect -2061 -3386 -2045 -3352
rect -2011 -3386 -1995 -3352
rect -1943 -3386 -1927 -3352
rect -1893 -3386 -1877 -3352
rect -1825 -3386 -1809 -3352
rect -1775 -3386 -1759 -3352
rect -1707 -3386 -1691 -3352
rect -1657 -3386 -1641 -3352
rect -2340 -3436 -2306 -3420
rect -2340 -5428 -2306 -5412
rect -2222 -3436 -2188 -3420
rect -2222 -5428 -2188 -5412
rect -2104 -3436 -2070 -3420
rect -2104 -5428 -2070 -5412
rect -1986 -3436 -1952 -3420
rect -1986 -5428 -1952 -5412
rect -1868 -3436 -1834 -3420
rect -1868 -5428 -1834 -5412
rect -1750 -3436 -1716 -3420
rect -1750 -5428 -1716 -5412
rect -1632 -3436 -1598 -3420
rect -1632 -5428 -1598 -5412
rect 1087 -3284 1183 -3250
rect 1961 -3284 2057 -3250
rect 1087 -3346 1121 -3284
rect 2023 -3346 2057 -3284
rect 1244 -3386 1260 -3352
rect 1294 -3386 1310 -3352
rect 1362 -3386 1378 -3352
rect 1412 -3386 1428 -3352
rect 1480 -3386 1496 -3352
rect 1530 -3386 1546 -3352
rect 1598 -3386 1614 -3352
rect 1648 -3386 1664 -3352
rect 1716 -3386 1732 -3352
rect 1766 -3386 1782 -3352
rect 1834 -3386 1850 -3352
rect 1884 -3386 1900 -3352
rect -1289 -3460 -1193 -3426
rect 797 -3460 893 -3426
rect -1289 -3522 -1255 -3460
rect 859 -3522 893 -3460
rect -1095 -3558 -1079 -3524
rect -1045 -3558 -1029 -3524
rect 633 -3558 649 -3524
rect 683 -3558 699 -3524
rect -1175 -3612 -1141 -3596
rect -1175 -4104 -1141 -4088
rect -1079 -3612 -1045 -3596
rect -1079 -4104 -1045 -4088
rect -983 -3612 -949 -3596
rect -983 -4104 -949 -4088
rect -887 -3612 -853 -3596
rect -887 -4104 -853 -4088
rect -791 -3612 -757 -3596
rect -791 -4104 -757 -4088
rect -695 -3612 -661 -3596
rect -695 -4104 -661 -4088
rect -599 -3612 -565 -3596
rect -599 -4104 -565 -4088
rect -503 -3612 -469 -3596
rect -503 -4104 -469 -4088
rect -407 -3612 -373 -3596
rect -407 -4104 -373 -4088
rect -311 -3612 -277 -3596
rect -311 -4104 -277 -4088
rect -215 -3612 -181 -3596
rect -215 -4104 -181 -4088
rect -119 -3612 -85 -3596
rect -119 -4104 -85 -4088
rect -23 -3612 11 -3596
rect -23 -4104 11 -4088
rect 73 -3612 107 -3596
rect 73 -4104 107 -4088
rect 169 -3612 203 -3596
rect 169 -4104 203 -4088
rect 265 -3612 299 -3596
rect 265 -4104 299 -4088
rect 361 -3612 395 -3596
rect 361 -4104 395 -4088
rect 457 -3612 491 -3596
rect 457 -4104 491 -4088
rect 553 -3612 587 -3596
rect 553 -4104 587 -4088
rect 649 -3612 683 -3596
rect 649 -4104 683 -4088
rect 745 -3612 779 -3596
rect 745 -4104 779 -4088
rect -1289 -4240 -1255 -4178
rect -903 -4184 -887 -4150
rect -853 -4184 -837 -4150
rect -711 -4184 -695 -4150
rect -661 -4184 -645 -4150
rect -519 -4184 -503 -4150
rect -469 -4184 -453 -4150
rect -327 -4184 -311 -4150
rect -277 -4184 -261 -4150
rect -135 -4184 -119 -4150
rect -85 -4184 -69 -4150
rect 57 -4184 73 -4150
rect 107 -4184 123 -4150
rect 249 -4184 265 -4150
rect 299 -4184 315 -4150
rect 441 -4184 457 -4150
rect 491 -4184 507 -4150
rect 859 -4240 893 -4178
rect -1289 -4274 -1193 -4240
rect 797 -4274 893 -4240
rect -2297 -5496 -2281 -5462
rect -2247 -5496 -2231 -5462
rect -2179 -5496 -2163 -5462
rect -2129 -5496 -2113 -5462
rect -2061 -5496 -2045 -5462
rect -2011 -5496 -1995 -5462
rect -1943 -5496 -1927 -5462
rect -1893 -5496 -1877 -5462
rect -1825 -5496 -1809 -5462
rect -1775 -5496 -1759 -5462
rect -1707 -5496 -1691 -5462
rect -1657 -5496 -1641 -5462
rect -2454 -5564 -2420 -5502
rect -1518 -5564 -1484 -5502
rect -2454 -5598 -2358 -5564
rect -1580 -5598 -1484 -5564
rect -1245 -4400 -1149 -4366
rect 753 -4400 849 -4366
rect -1245 -4462 -1211 -4400
rect 815 -4462 849 -4400
rect -1085 -4502 -1069 -4468
rect -701 -4502 -685 -4468
rect -627 -4502 -611 -4468
rect -243 -4502 -227 -4468
rect -169 -4502 -153 -4468
rect 215 -4502 231 -4468
rect 289 -4502 305 -4468
rect 673 -4502 689 -4468
rect -3758 -5784 -2842 -5750
rect -3758 -5818 -3628 -5784
rect -2972 -5818 -2842 -5784
rect -3758 -5880 -3690 -5818
rect -3758 -6730 -3724 -5880
rect -2910 -5880 -2842 -5818
rect -3554 -5932 -3538 -5898
rect -3062 -5932 -3046 -5898
rect -3622 -5964 -3588 -5948
rect -3622 -6014 -3588 -5998
rect -3554 -6028 -3538 -5994
rect -3062 -6028 -3046 -5994
rect -3554 -6124 -3538 -6090
rect -3062 -6124 -3046 -6090
rect -3622 -6156 -3588 -6140
rect -3622 -6206 -3588 -6190
rect -3554 -6220 -3538 -6186
rect -3062 -6220 -2910 -6186
rect -3633 -6316 -3538 -6282
rect -3062 -6316 -3046 -6282
rect -3633 -6434 -3582 -6316
rect -3633 -6504 -3594 -6434
rect -3633 -6608 -3594 -6600
rect -3633 -6661 -3610 -6608
rect -3633 -6670 -3594 -6661
rect -3758 -6812 -3690 -6730
rect -2876 -5920 -2842 -5880
rect -2876 -5940 -2720 -5920
rect -2876 -6730 -2800 -5940
rect -2910 -6812 -2800 -6730
rect -3758 -6846 -3628 -6812
rect -2972 -6846 -2800 -6812
rect -3758 -6860 -2800 -6846
rect -2740 -6860 -2720 -5940
rect -1131 -4552 -1097 -4536
rect -1131 -6544 -1097 -6528
rect -673 -4552 -639 -4536
rect -673 -6544 -639 -6528
rect -215 -4552 -181 -4536
rect -215 -6544 -181 -6528
rect 243 -4552 277 -4536
rect 243 -6544 277 -6528
rect 701 -4552 735 -4536
rect 701 -6544 735 -6528
rect 1201 -3436 1235 -3420
rect 1201 -5428 1235 -5412
rect 1319 -3436 1353 -3420
rect 1319 -5428 1353 -5412
rect 1437 -3436 1471 -3420
rect 1437 -5428 1471 -5412
rect 1555 -3436 1589 -3420
rect 1555 -5428 1589 -5412
rect 1673 -3436 1707 -3420
rect 1673 -5428 1707 -5412
rect 1791 -3436 1825 -3420
rect 1791 -5428 1825 -5412
rect 1909 -3436 1943 -3420
rect 1909 -5428 1943 -5412
rect 2128 -3640 2224 -3618
rect 2057 -3652 2224 -3640
rect 2664 -3652 2760 -3618
rect 2057 -3714 2162 -3652
rect 2057 -4818 2128 -3714
rect 2726 -3714 2760 -3652
rect 2057 -4880 2162 -4818
rect 2726 -4880 2760 -4818
rect 2128 -4914 2224 -4880
rect 2664 -4914 2760 -4880
rect 1244 -5496 1260 -5462
rect 1294 -5496 1310 -5462
rect 1362 -5496 1378 -5462
rect 1412 -5496 1428 -5462
rect 1480 -5496 1496 -5462
rect 1530 -5496 1546 -5462
rect 1598 -5496 1614 -5462
rect 1648 -5496 1664 -5462
rect 1716 -5496 1732 -5462
rect 1766 -5496 1782 -5462
rect 1834 -5496 1850 -5462
rect 1884 -5496 1900 -5462
rect 1087 -5564 1121 -5502
rect 2023 -5564 2057 -5502
rect 1087 -5598 1183 -5564
rect 1961 -5598 2057 -5564
rect -1085 -6612 -1069 -6578
rect -701 -6612 -685 -6578
rect -627 -6612 -611 -6578
rect -243 -6612 -227 -6578
rect -169 -6612 -153 -6578
rect 215 -6612 231 -6578
rect 289 -6612 305 -6578
rect 673 -6612 689 -6578
rect -1245 -6680 -1211 -6618
rect 815 -6680 849 -6618
rect -1245 -6714 -1149 -6680
rect 753 -6714 849 -6680
rect -3758 -6880 -2720 -6860
<< viali >>
rect -2044 -868 -2010 -834
rect -1926 -868 -1892 -834
rect -1808 -868 -1774 -834
rect -1690 -868 -1656 -834
rect -1572 -868 -1538 -834
rect -1454 -868 -1420 -834
rect -1336 -868 -1302 -834
rect -1218 -868 -1184 -834
rect -1100 -868 -1066 -834
rect -982 -868 -948 -834
rect -864 -868 -830 -834
rect -746 -868 -712 -834
rect 316 -868 350 -834
rect 434 -868 468 -834
rect 552 -868 586 -834
rect 670 -868 704 -834
rect 788 -868 822 -834
rect 906 -868 940 -834
rect 1024 -868 1058 -834
rect 1142 -868 1176 -834
rect 1260 -868 1294 -834
rect 1378 -868 1412 -834
rect 1496 -868 1530 -834
rect 1614 -868 1648 -834
rect -2217 -1315 -2183 -915
rect -2217 -2915 -2183 -2515
rect -2103 -2903 -2069 -927
rect -1985 -2903 -1951 -927
rect -1867 -2903 -1833 -927
rect -1749 -2903 -1715 -927
rect -1631 -2903 -1597 -927
rect -1513 -2903 -1479 -927
rect -1395 -2903 -1361 -927
rect -1277 -2903 -1243 -927
rect -1159 -2903 -1125 -927
rect -1041 -2903 -1007 -927
rect -923 -2903 -889 -927
rect -805 -2903 -771 -927
rect -687 -2903 -653 -927
rect -569 -2903 -535 -927
rect -451 -2903 -417 -927
rect -333 -2903 -299 -927
rect -215 -2903 -181 -927
rect -97 -2903 -63 -927
rect 21 -2903 55 -927
rect 139 -2903 173 -927
rect 257 -2903 291 -927
rect 375 -2903 409 -927
rect 493 -2903 527 -927
rect 611 -2903 645 -927
rect 729 -2903 763 -927
rect 847 -2903 881 -927
rect 965 -2903 999 -927
rect 1083 -2903 1117 -927
rect 1201 -2903 1235 -927
rect 1319 -2903 1353 -927
rect 1437 -2903 1471 -927
rect 1555 -2903 1589 -927
rect 1673 -2903 1707 -927
rect 1787 -1315 1821 -915
rect 1787 -2915 1821 -2515
rect -2044 -2996 -2010 -2962
rect -1926 -2996 -1892 -2962
rect -1808 -2996 -1774 -2962
rect -1690 -2996 -1656 -2962
rect -1572 -2996 -1538 -2962
rect -1454 -2996 -1420 -2962
rect -1336 -2996 -1302 -2962
rect -1218 -2996 -1184 -2962
rect -1100 -2996 -1066 -2962
rect -982 -2996 -948 -2962
rect -864 -2996 -830 -2962
rect -746 -2996 -712 -2962
rect -628 -2996 -594 -2962
rect -510 -2996 -476 -2962
rect -392 -2996 -358 -2962
rect -274 -2996 -240 -2962
rect -156 -2996 -122 -2962
rect -38 -2996 -4 -2962
rect 80 -2996 114 -2962
rect 198 -2996 232 -2962
rect 316 -2996 350 -2962
rect 434 -2996 468 -2962
rect 552 -2996 586 -2962
rect 670 -2996 704 -2962
rect 788 -2996 822 -2962
rect 906 -2996 940 -2962
rect 1024 -2996 1058 -2962
rect 1142 -2996 1176 -2962
rect 1260 -2996 1294 -2962
rect 1378 -2996 1412 -2962
rect 1496 -2996 1530 -2962
rect 1614 -2996 1648 -2962
rect -2281 -3386 -2247 -3352
rect -2163 -3386 -2129 -3352
rect -2045 -3386 -2011 -3352
rect -1927 -3386 -1893 -3352
rect -1809 -3386 -1775 -3352
rect -1691 -3386 -1657 -3352
rect -2454 -3824 -2420 -3424
rect -2454 -5424 -2420 -5024
rect -2340 -5412 -2306 -3436
rect -2222 -5412 -2188 -3436
rect -2104 -5412 -2070 -3436
rect -1986 -5412 -1952 -3436
rect -1868 -5412 -1834 -3436
rect -1750 -5412 -1716 -3436
rect -1632 -5412 -1598 -3436
rect -1518 -3824 -1484 -3424
rect 1260 -3386 1294 -3352
rect 1378 -3386 1412 -3352
rect 1496 -3386 1530 -3352
rect 1614 -3386 1648 -3352
rect 1732 -3386 1766 -3352
rect 1850 -3386 1884 -3352
rect -1079 -3558 -1045 -3524
rect 649 -3558 683 -3524
rect -1289 -4100 -1255 -3600
rect -1175 -4088 -1141 -3612
rect -1079 -4088 -1045 -3612
rect -983 -4088 -949 -3612
rect -887 -4088 -853 -3612
rect -791 -4088 -757 -3612
rect -695 -4088 -661 -3612
rect -599 -4088 -565 -3612
rect -503 -4088 -469 -3612
rect -407 -4088 -373 -3612
rect -311 -4088 -277 -3612
rect -215 -4088 -181 -3612
rect -119 -4088 -85 -3612
rect -23 -4088 11 -3612
rect 73 -4088 107 -3612
rect 169 -4088 203 -3612
rect 265 -4088 299 -3612
rect 361 -4088 395 -3612
rect 457 -4088 491 -3612
rect 553 -4088 587 -3612
rect 649 -4088 683 -3612
rect 745 -4088 779 -3612
rect 859 -4100 893 -3600
rect -887 -4184 -853 -4150
rect -695 -4184 -661 -4150
rect -503 -4184 -469 -4150
rect -311 -4184 -277 -4150
rect -119 -4184 -85 -4150
rect 73 -4184 107 -4150
rect 265 -4184 299 -4150
rect 457 -4184 491 -4150
rect 1087 -3824 1121 -3424
rect -1518 -5424 -1484 -5024
rect -2281 -5496 -2247 -5462
rect -2163 -5496 -2129 -5462
rect -2045 -5496 -2011 -5462
rect -1927 -5496 -1893 -5462
rect -1809 -5496 -1775 -5462
rect -1691 -5496 -1657 -5462
rect -1069 -4502 -701 -4468
rect -611 -4502 -243 -4468
rect -153 -4502 215 -4468
rect 305 -4502 673 -4468
rect -1245 -4940 -1211 -4540
rect -3538 -5932 -3062 -5898
rect -3622 -5998 -3588 -5964
rect -3538 -6028 -3062 -5994
rect -3538 -6124 -3062 -6090
rect -3622 -6190 -3588 -6156
rect -3538 -6220 -3062 -6186
rect -3538 -6316 -3062 -6282
rect -3610 -6661 -3594 -6608
rect -3594 -6661 -3178 -6608
rect -2800 -6860 -2740 -5940
rect -1245 -6540 -1211 -6140
rect -1131 -6528 -1097 -4552
rect -673 -6528 -639 -4552
rect -215 -6528 -181 -4552
rect 243 -6528 277 -4552
rect 701 -6528 735 -4552
rect 815 -4940 849 -4540
rect 1087 -5424 1121 -5024
rect 1201 -5412 1235 -3436
rect 1319 -5412 1353 -3436
rect 1437 -5412 1471 -3436
rect 1555 -5412 1589 -3436
rect 1673 -5412 1707 -3436
rect 1791 -5412 1825 -3436
rect 1909 -5412 1943 -3436
rect 2023 -3824 2057 -3424
rect 2272 -4160 2382 -3770
rect 2502 -4160 2612 -3770
rect 2023 -5424 2057 -5024
rect 1260 -5496 1294 -5462
rect 1378 -5496 1412 -5462
rect 1496 -5496 1530 -5462
rect 1614 -5496 1648 -5462
rect 1732 -5496 1766 -5462
rect 1850 -5496 1884 -5462
rect 815 -6540 849 -6140
rect -1069 -6612 -701 -6578
rect -611 -6612 -243 -6578
rect -153 -6612 215 -6578
rect 305 -6612 673 -6578
<< metal1 >>
rect -2112 -834 -1994 -828
rect -2112 -868 -2044 -834
rect -2010 -868 -1994 -834
rect -2112 -874 -1994 -868
rect -1942 -834 -696 -828
rect -1942 -868 -1926 -834
rect -1892 -868 -1808 -834
rect -1774 -868 -1690 -834
rect -1656 -868 -1572 -834
rect -1538 -868 -1454 -834
rect -1420 -868 -1336 -834
rect -1302 -868 -1218 -834
rect -1184 -868 -1100 -834
rect -1066 -868 -982 -834
rect -948 -868 -864 -834
rect -830 -868 -746 -834
rect -712 -868 -696 -834
rect -1942 -874 -696 -868
rect 300 -834 1546 -828
rect 300 -868 316 -834
rect 350 -868 434 -834
rect 468 -868 552 -834
rect 586 -868 670 -834
rect 704 -868 788 -834
rect 822 -868 906 -834
rect 940 -868 1024 -834
rect 1058 -868 1142 -834
rect 1176 -868 1260 -834
rect 1294 -868 1378 -834
rect 1412 -868 1496 -834
rect 1530 -868 1546 -834
rect 300 -874 1546 -868
rect 1598 -834 1716 -828
rect 1598 -868 1614 -834
rect 1648 -868 1716 -834
rect 1598 -874 1716 -868
rect -2223 -915 -2177 -903
rect -2112 -915 -2060 -874
rect -2223 -1315 -2217 -915
rect -2183 -927 -2060 -915
rect -2183 -1315 -2112 -927
rect -2223 -1327 -2177 -1315
rect -2223 -2515 -2177 -2503
rect -2223 -2915 -2217 -2515
rect -2183 -2903 -2112 -2515
rect -2183 -2915 -2060 -2903
rect -2223 -2927 -2177 -2915
rect -2112 -2956 -2060 -2915
rect -1994 -927 -1942 -915
rect -1994 -2916 -1942 -2903
rect -1876 -927 -1824 -915
rect -1876 -2915 -1824 -2903
rect -1758 -927 -1706 -915
rect -1758 -2915 -1706 -2903
rect -1640 -927 -1588 -915
rect -1640 -2915 -1588 -2903
rect -1522 -927 -1470 -915
rect -1522 -2915 -1470 -2903
rect -1404 -927 -1352 -915
rect -1404 -2915 -1352 -2903
rect -1286 -927 -1234 -915
rect -1286 -2915 -1234 -2903
rect -1168 -927 -1116 -915
rect -1168 -2915 -1116 -2903
rect -1050 -927 -998 -915
rect -1050 -2915 -998 -2903
rect -932 -927 -880 -915
rect -932 -2915 -880 -2903
rect -814 -927 -762 -874
rect -814 -2956 -762 -2903
rect -696 -927 -644 -915
rect -696 -2915 -644 -2903
rect -578 -927 -526 -914
rect -578 -2915 -526 -2903
rect -460 -927 -408 -915
rect -460 -2915 -408 -2903
rect -342 -927 -290 -915
rect -342 -2915 -290 -2903
rect -224 -927 -172 -915
rect -224 -2915 -172 -2903
rect -106 -927 -54 -915
rect -106 -2915 -54 -2903
rect 12 -927 64 -915
rect 12 -2915 64 -2903
rect 130 -927 182 -914
rect 130 -2915 182 -2903
rect 248 -927 300 -915
rect 248 -2915 300 -2903
rect 366 -927 418 -874
rect 1664 -915 1716 -874
rect 1781 -915 1827 -903
rect -290 -2956 -224 -2950
rect 366 -2956 418 -2903
rect 484 -927 536 -915
rect 484 -2915 536 -2903
rect 602 -927 654 -915
rect 602 -2915 654 -2903
rect 720 -927 772 -915
rect 720 -2915 772 -2903
rect 838 -927 890 -915
rect 838 -2915 890 -2903
rect 956 -927 1008 -915
rect 956 -2915 1008 -2903
rect 1074 -927 1126 -915
rect 1074 -2915 1126 -2903
rect 1192 -927 1244 -915
rect 1192 -2915 1244 -2903
rect 1310 -927 1362 -915
rect 1310 -2915 1362 -2903
rect 1428 -927 1480 -915
rect 1428 -2915 1480 -2903
rect 1546 -927 1598 -915
rect 1546 -2915 1598 -2903
rect 1664 -927 1787 -915
rect 1716 -1315 1787 -927
rect 1821 -1315 1827 -915
rect 1781 -1327 1827 -1315
rect 1781 -2515 1827 -2503
rect 1716 -2903 1787 -2515
rect 1664 -2915 1787 -2903
rect 1821 -2915 1827 -2515
rect 1664 -2956 1716 -2915
rect 1781 -2927 1827 -2915
rect -2112 -2962 -1994 -2956
rect -2112 -2996 -2044 -2962
rect -2010 -2996 -1994 -2962
rect -2112 -3002 -1994 -2996
rect -1942 -2962 -696 -2956
rect -1942 -2996 -1926 -2962
rect -1892 -2996 -1808 -2962
rect -1774 -2996 -1690 -2962
rect -1656 -2996 -1572 -2962
rect -1538 -2996 -1454 -2962
rect -1420 -2996 -1336 -2962
rect -1302 -2996 -1218 -2962
rect -1184 -2996 -1100 -2962
rect -1066 -2996 -982 -2962
rect -948 -2996 -864 -2962
rect -830 -2996 -746 -2962
rect -712 -2996 -696 -2962
rect -1942 -3002 -696 -2996
rect -644 -2962 -282 -2956
rect -644 -2996 -628 -2962
rect -594 -2996 -510 -2962
rect -476 -2996 -392 -2962
rect -358 -2996 -282 -2962
rect -644 -3002 -282 -2996
rect -290 -3008 -282 -3002
rect -230 -3008 -224 -2956
rect -168 -2962 248 -2956
rect -168 -2996 -156 -2962
rect -122 -2996 -38 -2962
rect -4 -2996 80 -2962
rect 114 -2996 198 -2962
rect 232 -2996 248 -2962
rect -168 -3000 248 -2996
rect -290 -3019 -224 -3008
rect -173 -3052 -167 -3000
rect -115 -3002 248 -3000
rect 300 -2962 1546 -2956
rect 300 -2996 316 -2962
rect 350 -2996 434 -2962
rect 468 -2996 552 -2962
rect 586 -2996 670 -2962
rect 704 -2996 788 -2962
rect 822 -2996 906 -2962
rect 940 -2996 1024 -2962
rect 1058 -2996 1142 -2962
rect 1176 -2996 1260 -2962
rect 1294 -2996 1378 -2962
rect 1412 -2996 1496 -2962
rect 1530 -2996 1546 -2962
rect 300 -3002 1546 -2996
rect 1598 -2962 1716 -2956
rect 1598 -2996 1614 -2962
rect 1648 -2996 1716 -2962
rect 1598 -3002 1716 -2996
rect -115 -3052 -109 -3002
rect -1995 -3242 -1943 -3236
rect -1995 -3346 -1943 -3294
rect 1546 -3242 1598 -3236
rect 1546 -3346 1598 -3294
rect -2349 -3352 -2231 -3346
rect -2349 -3386 -2281 -3352
rect -2247 -3386 -2231 -3352
rect -2349 -3392 -2231 -3386
rect -2179 -3352 -1763 -3346
rect -2179 -3386 -2163 -3352
rect -2129 -3386 -2045 -3352
rect -2011 -3386 -1927 -3352
rect -1893 -3386 -1809 -3352
rect -1775 -3386 -1763 -3352
rect -2179 -3392 -1763 -3386
rect -1703 -3352 -1589 -3346
rect -1703 -3386 -1691 -3352
rect -1657 -3386 -1589 -3352
rect -1703 -3392 -1589 -3386
rect -2460 -3424 -2414 -3412
rect -2349 -3424 -2297 -3392
rect -1641 -3424 -1589 -3392
rect 1192 -3352 1306 -3346
rect 1192 -3386 1260 -3352
rect 1294 -3386 1306 -3352
rect 1192 -3392 1306 -3386
rect 1366 -3352 1782 -3346
rect 1366 -3386 1378 -3352
rect 1412 -3386 1496 -3352
rect 1530 -3386 1614 -3352
rect 1648 -3386 1732 -3352
rect 1766 -3386 1782 -3352
rect 1366 -3392 1782 -3386
rect 1838 -3352 1952 -3346
rect 1838 -3386 1850 -3352
rect 1884 -3386 1952 -3352
rect 1838 -3392 1952 -3386
rect -1498 -3412 -1398 -3400
rect -1524 -3424 -1398 -3412
rect -2460 -3824 -2454 -3424
rect -2420 -3436 -2297 -3424
rect -2420 -3824 -2349 -3436
rect -2460 -3836 -2414 -3824
rect -2460 -5024 -2414 -5012
rect -2460 -5424 -2454 -5024
rect -2420 -5412 -2349 -5024
rect -2420 -5424 -2297 -5412
rect -2231 -3436 -2179 -3424
rect -2231 -5424 -2179 -5412
rect -2113 -3436 -2061 -3424
rect -2113 -5424 -2061 -5412
rect -1995 -3436 -1943 -3424
rect -1995 -5424 -1943 -5412
rect -1877 -3436 -1825 -3424
rect -1877 -5424 -1825 -5412
rect -1759 -3436 -1707 -3424
rect -1759 -5424 -1707 -5412
rect -1641 -3436 -1518 -3424
rect -1589 -3824 -1518 -3436
rect -1484 -3500 -1398 -3424
rect 1002 -3412 1102 -3400
rect 1002 -3424 1127 -3412
rect 1192 -3424 1244 -3392
rect 1900 -3424 1952 -3392
rect 2017 -3424 2063 -3412
rect 1002 -3500 1087 -3424
rect -1484 -3600 -1238 -3500
rect -1181 -3524 -1029 -3518
rect -1181 -3558 -1079 -3524
rect -1045 -3558 -1029 -3524
rect -1181 -3564 -1029 -3558
rect 633 -3524 785 -3518
rect 633 -3558 649 -3524
rect 683 -3558 785 -3524
rect 633 -3564 785 -3558
rect -1181 -3600 -1135 -3564
rect -1085 -3600 -1039 -3564
rect 643 -3600 689 -3564
rect 739 -3600 785 -3564
rect 842 -3600 1087 -3500
rect -1484 -3824 -1289 -3600
rect -1524 -3836 -1289 -3824
rect -1498 -4000 -1289 -3836
rect -1398 -4100 -1289 -4000
rect -1255 -4100 -1185 -3600
rect -1131 -4100 -1125 -3600
rect -1095 -4100 -1089 -3600
rect -1035 -4100 -1029 -3600
rect -999 -4100 -993 -3600
rect -939 -4100 -933 -3600
rect -903 -4100 -897 -3600
rect -843 -4100 -837 -3600
rect -807 -4100 -801 -3600
rect -747 -4100 -741 -3600
rect -711 -4100 -705 -3600
rect -651 -4100 -645 -3600
rect -615 -4100 -609 -3600
rect -555 -4100 -549 -3600
rect -519 -4100 -513 -3600
rect -459 -4100 -453 -3600
rect -423 -4100 -417 -3600
rect -363 -4100 -357 -3600
rect -327 -4100 -321 -3600
rect -267 -4100 -261 -3600
rect -231 -4100 -225 -3600
rect -171 -4100 -165 -3600
rect -135 -4100 -129 -3600
rect -75 -4100 -69 -3600
rect -39 -4100 -33 -3600
rect 21 -4100 27 -3600
rect 57 -4100 63 -3600
rect 117 -4100 123 -3600
rect 153 -4100 159 -3600
rect 213 -4100 219 -3600
rect 249 -4100 255 -3600
rect 309 -4100 315 -3600
rect 345 -4100 351 -3600
rect 405 -4100 411 -3600
rect 441 -4100 447 -3600
rect 501 -4100 507 -3600
rect 537 -4100 543 -3600
rect 597 -4100 603 -3600
rect 633 -4100 639 -3600
rect 693 -4100 699 -3600
rect 729 -4100 735 -3600
rect 789 -4100 859 -3600
rect 893 -3824 1087 -3600
rect 1121 -3436 1244 -3424
rect 1121 -3824 1192 -3436
rect 893 -3836 1127 -3824
rect 893 -4000 1102 -3836
rect 893 -4100 1002 -4000
rect -1398 -4400 -1238 -4100
rect -909 -4200 -903 -4144
rect -837 -4200 -831 -4144
rect -717 -4200 -711 -4144
rect -645 -4200 -639 -4144
rect -525 -4200 -519 -4144
rect -453 -4200 -447 -4144
rect -333 -4200 -327 -4144
rect -261 -4200 -255 -4144
rect -141 -4200 -135 -4144
rect -69 -4200 -63 -4144
rect 51 -4200 57 -4144
rect 123 -4200 129 -4144
rect 243 -4200 249 -4144
rect 315 -4200 321 -4144
rect 435 -4200 441 -4144
rect 507 -4200 513 -4144
rect -1398 -4540 -1198 -4400
rect -1142 -4438 -1078 -4430
rect -1078 -4468 685 -4462
rect -1078 -4502 -1069 -4468
rect -701 -4502 -611 -4468
rect -243 -4502 -153 -4468
rect 215 -4502 305 -4468
rect 673 -4502 685 -4468
rect -1142 -4508 685 -4502
rect -1142 -4510 -1078 -4508
rect 842 -4528 1002 -4100
rect 809 -4540 1002 -4528
rect -1398 -4900 -1245 -4540
rect -1498 -4940 -1245 -4900
rect -1211 -4552 -1088 -4540
rect -1211 -4940 -1140 -4552
rect -1498 -5000 -1198 -4940
rect -1498 -5012 -1238 -5000
rect -1524 -5024 -1238 -5012
rect -1589 -5412 -1518 -5024
rect -1641 -5424 -1518 -5412
rect -1484 -5424 -1238 -5024
rect -2460 -5436 -2414 -5424
rect -2349 -5456 -2297 -5424
rect -1641 -5456 -1589 -5424
rect -1524 -5436 -1238 -5424
rect -2349 -5462 -2231 -5456
rect -2349 -5496 -2281 -5462
rect -2247 -5496 -2231 -5462
rect -2349 -5502 -2231 -5496
rect -2179 -5462 -1763 -5456
rect -2179 -5496 -2163 -5462
rect -2129 -5496 -2045 -5462
rect -2011 -5496 -1927 -5462
rect -1893 -5496 -1809 -5462
rect -1775 -5496 -1763 -5462
rect -2179 -5502 -1763 -5496
rect -1703 -5462 -1589 -5456
rect -1703 -5496 -1691 -5462
rect -1657 -5496 -1589 -5462
rect -1703 -5502 -1589 -5496
rect -1498 -5500 -1238 -5436
rect -1398 -5560 -1238 -5500
rect -3550 -5898 -2942 -5892
rect -3550 -5932 -3538 -5898
rect -3062 -5932 -2942 -5898
rect -3550 -5938 -2942 -5932
rect -3628 -5964 -3582 -5948
rect -3628 -5994 -3622 -5964
rect -3763 -5998 -3622 -5994
rect -3588 -5998 -3582 -5964
rect -3763 -6028 -3582 -5998
rect -3551 -5994 -3534 -5985
rect -3065 -5994 -3050 -5985
rect -3551 -6028 -3538 -5994
rect -3062 -6028 -3050 -5994
rect -3763 -6884 -3729 -6028
rect -3551 -6037 -3534 -6028
rect -3065 -6037 -3050 -6028
rect -2982 -6084 -2942 -5938
rect -3550 -6090 -2942 -6084
rect -3550 -6124 -3538 -6090
rect -3062 -6124 -2942 -6090
rect -3550 -6130 -2942 -6124
rect -3628 -6156 -3582 -6140
rect -3628 -6186 -3622 -6156
rect -3769 -7084 -3729 -6884
rect -3701 -6190 -3622 -6186
rect -3588 -6190 -3582 -6156
rect -3701 -6220 -3582 -6190
rect -3550 -6186 -3050 -6180
rect -3550 -6220 -3538 -6186
rect -3062 -6220 -3050 -6186
rect -3701 -6884 -3667 -6220
rect -3550 -6226 -3050 -6220
rect -2982 -6276 -2942 -6130
rect -3550 -6282 -2942 -6276
rect -3550 -6316 -3538 -6282
rect -3062 -6316 -2942 -6282
rect -3550 -6322 -2942 -6316
rect -2820 -5940 -2580 -5920
rect -3633 -6670 -3610 -6600
rect -3181 -6608 -3162 -6600
rect -3178 -6661 -3162 -6608
rect -3181 -6670 -3162 -6661
rect -2820 -6860 -2800 -5940
rect -2600 -6860 -2580 -5940
rect -1398 -6780 -1378 -5560
rect -1318 -6128 -1238 -5560
rect -1318 -6140 -1205 -6128
rect -1318 -6540 -1245 -6140
rect -1211 -6528 -1140 -6140
rect -1211 -6540 -1088 -6528
rect -682 -4552 -630 -4540
rect -682 -6540 -630 -6528
rect -224 -4552 -172 -4540
rect -224 -6540 -172 -6528
rect 234 -4552 286 -4540
rect 234 -6540 286 -6528
rect 692 -4552 815 -4540
rect 744 -4940 815 -4552
rect 849 -4900 1002 -4540
rect 849 -4940 1102 -4900
rect 809 -4952 1102 -4940
rect 842 -5012 1102 -4952
rect 842 -5024 1127 -5012
rect 842 -5424 1087 -5024
rect 1121 -5412 1192 -5024
rect 1121 -5424 1244 -5412
rect 1310 -3436 1362 -3424
rect 1310 -5424 1362 -5412
rect 1428 -3436 1480 -3424
rect 1428 -5424 1480 -5412
rect 1546 -3436 1598 -3424
rect 1546 -5424 1598 -5412
rect 1664 -3436 1716 -3424
rect 1664 -5424 1716 -5412
rect 1782 -3436 1834 -3424
rect 1782 -5424 1834 -5412
rect 1900 -3436 2023 -3424
rect 1952 -3824 2023 -3436
rect 2057 -3824 2063 -3424
rect 2017 -3836 2063 -3824
rect 2252 -3770 2402 -3750
rect 2252 -4160 2272 -3770
rect 2382 -4160 2402 -3770
rect 2252 -4180 2402 -4160
rect 2482 -3770 2632 -3750
rect 2482 -4160 2502 -3770
rect 2612 -4160 2632 -3770
rect 2482 -4180 2632 -4160
rect 2017 -5024 2063 -5012
rect 1952 -5412 2023 -5024
rect 1900 -5424 2023 -5412
rect 2057 -5424 2063 -5024
rect 842 -5436 1127 -5424
rect 842 -5500 1102 -5436
rect 1192 -5456 1244 -5424
rect 1900 -5456 1952 -5424
rect 2017 -5436 2063 -5424
rect 1192 -5462 1306 -5456
rect 1192 -5496 1260 -5462
rect 1294 -5496 1306 -5462
rect 842 -5560 1002 -5500
rect 1192 -5502 1306 -5496
rect 1366 -5462 1782 -5456
rect 1366 -5496 1378 -5462
rect 1412 -5496 1496 -5462
rect 1530 -5496 1614 -5462
rect 1648 -5496 1732 -5462
rect 1766 -5496 1782 -5462
rect 1366 -5502 1782 -5496
rect 1838 -5462 1952 -5456
rect 1838 -5496 1850 -5462
rect 1884 -5496 1952 -5462
rect 1838 -5502 1952 -5496
rect 842 -6128 922 -5560
rect 809 -6140 922 -6128
rect 744 -6528 815 -6140
rect 692 -6540 815 -6528
rect 849 -6540 922 -6140
rect -1318 -6552 -1205 -6540
rect 809 -6552 922 -6540
rect -1318 -6780 -1238 -6552
rect -1081 -6578 685 -6572
rect -1081 -6612 -1069 -6578
rect -701 -6612 -611 -6578
rect -243 -6612 -153 -6578
rect 215 -6612 305 -6578
rect 673 -6612 685 -6578
rect -1081 -6618 685 -6612
rect -1398 -6800 -1238 -6780
rect 842 -6780 922 -6552
rect 982 -6780 1002 -5560
rect 842 -6800 1002 -6780
rect -2820 -6880 -2580 -6860
rect -3701 -7084 -3661 -6884
<< via1 >>
rect -2112 -2903 -2103 -927
rect -2103 -2903 -2069 -927
rect -2069 -2903 -2060 -927
rect -1994 -2903 -1985 -927
rect -1985 -2903 -1951 -927
rect -1951 -2903 -1942 -927
rect -1876 -2903 -1867 -927
rect -1867 -2903 -1833 -927
rect -1833 -2903 -1824 -927
rect -1758 -2903 -1749 -927
rect -1749 -2903 -1715 -927
rect -1715 -2903 -1706 -927
rect -1640 -2903 -1631 -927
rect -1631 -2903 -1597 -927
rect -1597 -2903 -1588 -927
rect -1522 -2903 -1513 -927
rect -1513 -2903 -1479 -927
rect -1479 -2903 -1470 -927
rect -1404 -2903 -1395 -927
rect -1395 -2903 -1361 -927
rect -1361 -2903 -1352 -927
rect -1286 -2903 -1277 -927
rect -1277 -2903 -1243 -927
rect -1243 -2903 -1234 -927
rect -1168 -2903 -1159 -927
rect -1159 -2903 -1125 -927
rect -1125 -2903 -1116 -927
rect -1050 -2903 -1041 -927
rect -1041 -2903 -1007 -927
rect -1007 -2903 -998 -927
rect -932 -2903 -923 -927
rect -923 -2903 -889 -927
rect -889 -2903 -880 -927
rect -814 -2903 -805 -927
rect -805 -2903 -771 -927
rect -771 -2903 -762 -927
rect -696 -2903 -687 -927
rect -687 -2903 -653 -927
rect -653 -2903 -644 -927
rect -578 -2903 -569 -927
rect -569 -2903 -535 -927
rect -535 -2903 -526 -927
rect -460 -2903 -451 -927
rect -451 -2903 -417 -927
rect -417 -2903 -408 -927
rect -342 -2903 -333 -927
rect -333 -2903 -299 -927
rect -299 -2903 -290 -927
rect -224 -2903 -215 -927
rect -215 -2903 -181 -927
rect -181 -2903 -172 -927
rect -106 -2903 -97 -927
rect -97 -2903 -63 -927
rect -63 -2903 -54 -927
rect 12 -2903 21 -927
rect 21 -2903 55 -927
rect 55 -2903 64 -927
rect 130 -2903 139 -927
rect 139 -2903 173 -927
rect 173 -2903 182 -927
rect 248 -2903 257 -927
rect 257 -2903 291 -927
rect 291 -2903 300 -927
rect 366 -2903 375 -927
rect 375 -2903 409 -927
rect 409 -2903 418 -927
rect 484 -2903 493 -927
rect 493 -2903 527 -927
rect 527 -2903 536 -927
rect 602 -2903 611 -927
rect 611 -2903 645 -927
rect 645 -2903 654 -927
rect 720 -2903 729 -927
rect 729 -2903 763 -927
rect 763 -2903 772 -927
rect 838 -2903 847 -927
rect 847 -2903 881 -927
rect 881 -2903 890 -927
rect 956 -2903 965 -927
rect 965 -2903 999 -927
rect 999 -2903 1008 -927
rect 1074 -2903 1083 -927
rect 1083 -2903 1117 -927
rect 1117 -2903 1126 -927
rect 1192 -2903 1201 -927
rect 1201 -2903 1235 -927
rect 1235 -2903 1244 -927
rect 1310 -2903 1319 -927
rect 1319 -2903 1353 -927
rect 1353 -2903 1362 -927
rect 1428 -2903 1437 -927
rect 1437 -2903 1471 -927
rect 1471 -2903 1480 -927
rect 1546 -2903 1555 -927
rect 1555 -2903 1589 -927
rect 1589 -2903 1598 -927
rect 1664 -2903 1673 -927
rect 1673 -2903 1707 -927
rect 1707 -2903 1716 -927
rect -282 -2962 -230 -2956
rect -282 -2996 -274 -2962
rect -274 -2996 -240 -2962
rect -240 -2996 -230 -2962
rect -282 -3008 -230 -2996
rect -167 -3052 -115 -3000
rect -1995 -3294 -1943 -3242
rect 1546 -3294 1598 -3242
rect -2349 -5412 -2340 -3436
rect -2340 -5412 -2306 -3436
rect -2306 -5412 -2297 -3436
rect -2231 -5412 -2222 -3436
rect -2222 -5412 -2188 -3436
rect -2188 -5412 -2179 -3436
rect -2113 -5412 -2104 -3436
rect -2104 -5412 -2070 -3436
rect -2070 -5412 -2061 -3436
rect -1995 -5412 -1986 -3436
rect -1986 -5412 -1952 -3436
rect -1952 -5412 -1943 -3436
rect -1877 -5412 -1868 -3436
rect -1868 -5412 -1834 -3436
rect -1834 -5412 -1825 -3436
rect -1759 -5412 -1750 -3436
rect -1750 -5412 -1716 -3436
rect -1716 -5412 -1707 -3436
rect -1641 -5412 -1632 -3436
rect -1632 -5412 -1598 -3436
rect -1598 -5412 -1589 -3436
rect -1185 -3612 -1131 -3600
rect -1185 -4088 -1175 -3612
rect -1175 -4088 -1141 -3612
rect -1141 -4088 -1131 -3612
rect -1185 -4100 -1131 -4088
rect -1089 -3612 -1035 -3600
rect -1089 -4088 -1079 -3612
rect -1079 -4088 -1045 -3612
rect -1045 -4088 -1035 -3612
rect -1089 -4100 -1035 -4088
rect -993 -3612 -939 -3600
rect -993 -4088 -983 -3612
rect -983 -4088 -949 -3612
rect -949 -4088 -939 -3612
rect -993 -4100 -939 -4088
rect -897 -3612 -843 -3600
rect -897 -4088 -887 -3612
rect -887 -4088 -853 -3612
rect -853 -4088 -843 -3612
rect -897 -4100 -843 -4088
rect -801 -3612 -747 -3600
rect -801 -4088 -791 -3612
rect -791 -4088 -757 -3612
rect -757 -4088 -747 -3612
rect -801 -4100 -747 -4088
rect -705 -3612 -651 -3600
rect -705 -4088 -695 -3612
rect -695 -4088 -661 -3612
rect -661 -4088 -651 -3612
rect -705 -4100 -651 -4088
rect -609 -3612 -555 -3600
rect -609 -4088 -599 -3612
rect -599 -4088 -565 -3612
rect -565 -4088 -555 -3612
rect -609 -4100 -555 -4088
rect -513 -3612 -459 -3600
rect -513 -4088 -503 -3612
rect -503 -4088 -469 -3612
rect -469 -4088 -459 -3612
rect -513 -4100 -459 -4088
rect -417 -3612 -363 -3600
rect -417 -4088 -407 -3612
rect -407 -4088 -373 -3612
rect -373 -4088 -363 -3612
rect -417 -4100 -363 -4088
rect -321 -3612 -267 -3600
rect -321 -4088 -311 -3612
rect -311 -4088 -277 -3612
rect -277 -4088 -267 -3612
rect -321 -4100 -267 -4088
rect -225 -3612 -171 -3600
rect -225 -4088 -215 -3612
rect -215 -4088 -181 -3612
rect -181 -4088 -171 -3612
rect -225 -4100 -171 -4088
rect -129 -3612 -75 -3600
rect -129 -4088 -119 -3612
rect -119 -4088 -85 -3612
rect -85 -4088 -75 -3612
rect -129 -4100 -75 -4088
rect -33 -3612 21 -3600
rect -33 -4088 -23 -3612
rect -23 -4088 11 -3612
rect 11 -4088 21 -3612
rect -33 -4100 21 -4088
rect 63 -3612 117 -3600
rect 63 -4088 73 -3612
rect 73 -4088 107 -3612
rect 107 -4088 117 -3612
rect 63 -4100 117 -4088
rect 159 -3612 213 -3600
rect 159 -4088 169 -3612
rect 169 -4088 203 -3612
rect 203 -4088 213 -3612
rect 159 -4100 213 -4088
rect 255 -3612 309 -3600
rect 255 -4088 265 -3612
rect 265 -4088 299 -3612
rect 299 -4088 309 -3612
rect 255 -4100 309 -4088
rect 351 -3612 405 -3600
rect 351 -4088 361 -3612
rect 361 -4088 395 -3612
rect 395 -4088 405 -3612
rect 351 -4100 405 -4088
rect 447 -3612 501 -3600
rect 447 -4088 457 -3612
rect 457 -4088 491 -3612
rect 491 -4088 501 -3612
rect 447 -4100 501 -4088
rect 543 -3612 597 -3600
rect 543 -4088 553 -3612
rect 553 -4088 587 -3612
rect 587 -4088 597 -3612
rect 543 -4100 597 -4088
rect 639 -3612 693 -3600
rect 639 -4088 649 -3612
rect 649 -4088 683 -3612
rect 683 -4088 693 -3612
rect 639 -4100 693 -4088
rect 735 -3612 789 -3600
rect 735 -4088 745 -3612
rect 745 -4088 779 -3612
rect 779 -4088 789 -3612
rect 735 -4100 789 -4088
rect -903 -4150 -837 -4144
rect -903 -4184 -887 -4150
rect -887 -4184 -853 -4150
rect -853 -4184 -837 -4150
rect -903 -4200 -837 -4184
rect -711 -4150 -645 -4144
rect -711 -4184 -695 -4150
rect -695 -4184 -661 -4150
rect -661 -4184 -645 -4150
rect -711 -4200 -645 -4184
rect -519 -4150 -453 -4144
rect -519 -4184 -503 -4150
rect -503 -4184 -469 -4150
rect -469 -4184 -453 -4150
rect -519 -4200 -453 -4184
rect -327 -4150 -261 -4144
rect -327 -4184 -311 -4150
rect -311 -4184 -277 -4150
rect -277 -4184 -261 -4150
rect -327 -4200 -261 -4184
rect -135 -4150 -69 -4144
rect -135 -4184 -119 -4150
rect -119 -4184 -85 -4150
rect -85 -4184 -69 -4150
rect -135 -4200 -69 -4184
rect 57 -4150 123 -4144
rect 57 -4184 73 -4150
rect 73 -4184 107 -4150
rect 107 -4184 123 -4150
rect 57 -4200 123 -4184
rect 249 -4150 315 -4144
rect 249 -4184 265 -4150
rect 265 -4184 299 -4150
rect 299 -4184 315 -4150
rect 249 -4200 315 -4184
rect 441 -4150 507 -4144
rect 441 -4184 457 -4150
rect 457 -4184 491 -4150
rect 491 -4184 507 -4150
rect 441 -4200 507 -4184
rect -1142 -4502 -1078 -4438
rect -3534 -5994 -3065 -5985
rect -3534 -6028 -3065 -5994
rect -3534 -6037 -3065 -6028
rect -3610 -6608 -3181 -6600
rect -3610 -6661 -3181 -6608
rect -3610 -6670 -3181 -6661
rect -2800 -6860 -2740 -5940
rect -2740 -6860 -2600 -5940
rect -1378 -6780 -1318 -5560
rect -1140 -6528 -1131 -4552
rect -1131 -6528 -1097 -4552
rect -1097 -6528 -1088 -4552
rect -682 -6528 -673 -4552
rect -673 -6528 -639 -4552
rect -639 -6528 -630 -4552
rect -224 -6528 -215 -4552
rect -215 -6528 -181 -4552
rect -181 -6528 -172 -4552
rect 234 -6528 243 -4552
rect 243 -6528 277 -4552
rect 277 -6528 286 -4552
rect 692 -6528 701 -4552
rect 701 -6528 735 -4552
rect 735 -6528 744 -4552
rect 1192 -5412 1201 -3436
rect 1201 -5412 1235 -3436
rect 1235 -5412 1244 -3436
rect 1310 -5412 1319 -3436
rect 1319 -5412 1353 -3436
rect 1353 -5412 1362 -3436
rect 1428 -5412 1437 -3436
rect 1437 -5412 1471 -3436
rect 1471 -5412 1480 -3436
rect 1546 -5412 1555 -3436
rect 1555 -5412 1589 -3436
rect 1589 -5412 1598 -3436
rect 1664 -5412 1673 -3436
rect 1673 -5412 1707 -3436
rect 1707 -5412 1716 -3436
rect 1782 -5412 1791 -3436
rect 1791 -5412 1825 -3436
rect 1825 -5412 1834 -3436
rect 1900 -5412 1909 -3436
rect 1909 -5412 1943 -3436
rect 1943 -5412 1952 -3436
rect 2272 -4160 2382 -3770
rect 2502 -4160 2612 -3770
rect 922 -6780 982 -5560
<< metal2 >>
rect -2000 0 1400 100
rect -2000 -400 -1900 0
rect -2090 -500 -1900 -400
rect 1300 -400 1400 0
rect 1300 -500 1694 -400
rect -2090 -600 1694 -500
rect -2090 -664 -1990 -600
rect -1598 -664 -1498 -600
rect -1198 -664 -1098 -600
rect -798 -664 -698 -600
rect -398 -664 -298 -600
rect -98 -664 2 -600
rect 302 -664 402 -600
rect 702 -664 802 -600
rect 1102 -664 1202 -600
rect 1594 -664 1694 -600
rect -2112 -766 1716 -664
rect -2112 -927 -2060 -766
rect -2112 -2915 -2060 -2903
rect -1994 -927 -1942 -915
rect -1994 -3012 -1942 -2903
rect -1876 -927 -1824 -766
rect -1876 -2915 -1824 -2903
rect -1758 -927 -1706 -915
rect -1758 -3012 -1706 -2903
rect -1640 -927 -1588 -766
rect -1640 -2915 -1588 -2903
rect -1522 -927 -1470 -915
rect -1522 -3012 -1470 -2903
rect -1404 -927 -1352 -766
rect -1404 -2915 -1352 -2903
rect -1286 -927 -1234 -915
rect -1286 -3012 -1234 -2903
rect -1168 -927 -1116 -766
rect -1168 -2915 -1116 -2903
rect -1050 -927 -998 -915
rect -1994 -3064 -1234 -3012
rect -1050 -3012 -998 -2903
rect -932 -927 -880 -766
rect -932 -2915 -880 -2903
rect -814 -927 -762 -915
rect -814 -3012 -762 -2903
rect -696 -927 -644 -766
rect -696 -2915 -644 -2903
rect -578 -927 -526 -915
rect -578 -2915 -526 -2903
rect -460 -927 -408 -766
rect -460 -2915 -408 -2903
rect -342 -927 -290 -915
rect -342 -2922 -290 -2903
rect -224 -927 -172 -766
rect -224 -2916 -172 -2903
rect -106 -927 -54 -915
rect -342 -3012 -310 -2922
rect -106 -2944 -54 -2903
rect 12 -927 64 -766
rect 12 -2915 64 -2903
rect 130 -927 182 -915
rect 130 -2915 182 -2903
rect 248 -927 300 -766
rect 248 -2915 300 -2903
rect 366 -927 418 -915
rect -258 -2950 -52 -2944
rect -1050 -3042 -310 -3012
rect -282 -2956 -52 -2950
rect -230 -2972 -52 -2956
rect -282 -3014 -230 -3008
rect -173 -3042 -167 -3000
rect -1050 -3052 -167 -3042
rect -115 -3052 -109 -3000
rect -1050 -3064 -109 -3052
rect -81 -3012 -52 -2972
rect 366 -3010 418 -2903
rect 484 -927 536 -766
rect 602 -927 654 -915
rect 484 -2915 536 -2903
rect 601 -2903 602 -2835
rect 601 -2915 654 -2903
rect 720 -927 772 -766
rect 838 -927 890 -915
rect 720 -2915 772 -2903
rect 837 -2903 838 -2835
rect 837 -2915 890 -2903
rect 956 -927 1008 -766
rect 1074 -927 1126 -915
rect 956 -2915 1008 -2903
rect 1073 -2903 1074 -2835
rect 1073 -2915 1126 -2903
rect 1192 -927 1244 -766
rect 1310 -927 1362 -915
rect 1192 -2915 1244 -2903
rect 1309 -2903 1310 -2835
rect 1309 -2915 1362 -2903
rect 1428 -927 1480 -766
rect 1546 -927 1598 -915
rect 1428 -2915 1480 -2903
rect 1545 -2903 1546 -2835
rect 182 -3011 418 -3010
rect 601 -3011 653 -2915
rect 182 -3012 653 -3011
rect -81 -3062 653 -3012
rect -81 -3064 182 -3062
rect 366 -3063 653 -3062
rect 837 -3012 889 -2915
rect 1073 -3012 1125 -2915
rect 1309 -3012 1361 -2915
rect 1545 -3012 1598 -2903
rect 1664 -927 1716 -766
rect 1664 -2915 1716 -2903
rect -1758 -3134 -1706 -3064
rect -2113 -3186 -1706 -3134
rect -2113 -3231 -2061 -3186
rect -1877 -3231 -1825 -3186
rect -2113 -3240 -1825 -3231
rect -2113 -3296 -1997 -3240
rect -1941 -3296 -1825 -3240
rect -2113 -3305 -1825 -3296
rect -2349 -3436 -2297 -3424
rect -2349 -5564 -2297 -5412
rect -2231 -3436 -2179 -3424
rect -2231 -5564 -2179 -5412
rect -2113 -3436 -2061 -3305
rect -2113 -5424 -2061 -5412
rect -1995 -3436 -1943 -3424
rect -1995 -5564 -1943 -5412
rect -1877 -3436 -1825 -3305
rect -814 -3390 -762 -3064
rect -342 -3070 -109 -3064
rect 366 -3390 418 -3063
rect 837 -3064 1598 -3012
rect 1672 -3060 1802 -3050
rect 1309 -3134 1361 -3064
rect 1672 -3134 1682 -3060
rect 1309 -3150 1682 -3134
rect 1792 -3150 1802 -3060
rect 1309 -3186 1802 -3150
rect -1877 -5424 -1825 -5412
rect -1759 -3436 -1707 -3424
rect -1759 -5540 -1707 -5412
rect -1641 -3436 -1589 -3424
rect -903 -3530 -261 -3390
rect -903 -3600 -837 -3530
rect -711 -3600 -645 -3530
rect -519 -3600 -453 -3530
rect -327 -3600 -261 -3530
rect -135 -3530 507 -3390
rect -135 -3600 -69 -3530
rect 57 -3600 123 -3530
rect 249 -3600 315 -3530
rect 441 -3600 507 -3530
rect 1192 -3436 1244 -3424
rect -1191 -4100 -1185 -3600
rect -1131 -4100 -1125 -3600
rect -1095 -4100 -1089 -3600
rect -1035 -4100 -1029 -3600
rect -999 -4100 -993 -3600
rect -939 -4100 -933 -3600
rect -903 -4100 -897 -3600
rect -843 -4100 -837 -3600
rect -807 -4100 -801 -3600
rect -747 -4100 -741 -3600
rect -711 -4100 -705 -3600
rect -651 -4100 -645 -3600
rect -615 -4100 -609 -3600
rect -555 -4100 -549 -3600
rect -519 -4100 -513 -3600
rect -459 -4100 -453 -3600
rect -423 -4100 -417 -3600
rect -363 -4100 -357 -3600
rect -327 -4100 -321 -3600
rect -267 -4100 -261 -3600
rect -231 -4100 -225 -3600
rect -171 -4100 -165 -3600
rect -135 -4100 -129 -3600
rect -75 -4100 -69 -3600
rect -39 -4100 -33 -3600
rect 21 -4100 27 -3600
rect 57 -4100 63 -3600
rect 117 -4100 123 -3600
rect 153 -4100 159 -3600
rect 213 -4100 219 -3600
rect 249 -4100 255 -3600
rect 309 -4100 315 -3600
rect 345 -4100 351 -3600
rect 405 -4100 411 -3600
rect 441 -4100 447 -3600
rect 501 -4100 507 -3600
rect 537 -4100 543 -3600
rect 597 -4100 603 -3600
rect 633 -4100 639 -3600
rect 693 -4100 699 -3600
rect 729 -4100 735 -3600
rect 789 -4100 795 -3600
rect -993 -4260 -939 -4100
rect -903 -4144 -837 -4138
rect -903 -4220 -837 -4206
rect -801 -4260 -747 -4100
rect -711 -4144 -645 -4138
rect -711 -4220 -645 -4206
rect -609 -4260 -555 -4100
rect -519 -4144 -453 -4138
rect -519 -4220 -453 -4206
rect -417 -4260 -363 -4100
rect -327 -4144 -261 -4138
rect -327 -4220 -261 -4206
rect -225 -4260 -171 -4100
rect -135 -4144 -69 -4138
rect -135 -4220 -69 -4206
rect -33 -4260 21 -4100
rect 57 -4144 123 -4138
rect 57 -4220 123 -4206
rect 159 -4260 213 -4100
rect 249 -4144 315 -4138
rect 249 -4220 315 -4206
rect 351 -4260 405 -4100
rect 441 -4144 507 -4138
rect 441 -4220 507 -4206
rect 543 -4260 597 -4100
rect -993 -4330 597 -4260
rect -993 -4416 -939 -4330
rect -801 -4416 -747 -4330
rect -609 -4416 -555 -4330
rect -417 -4416 -363 -4330
rect -225 -4416 -171 -4330
rect -33 -4416 21 -4330
rect 159 -4416 213 -4330
rect 351 -4416 405 -4330
rect 543 -4416 597 -4330
rect -1400 -4438 -1078 -4430
rect -1400 -4440 -1142 -4438
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1142 -4440
rect -1400 -4502 -1142 -4500
rect -1400 -4510 -1078 -4502
rect -993 -4508 597 -4416
rect -1641 -5540 -1589 -5412
rect -1140 -4552 -1088 -4540
rect -1759 -5560 -1298 -5540
rect -1759 -5564 -1378 -5560
rect -2398 -5634 -1378 -5564
rect -3300 -5768 -3050 -5749
rect -3300 -5985 -3280 -5768
rect -3070 -5985 -3050 -5768
rect -2398 -5800 -2298 -5634
rect -2198 -5800 -2098 -5634
rect -1998 -5800 -1898 -5634
rect -1798 -5640 -1378 -5634
rect -1798 -5800 -1698 -5640
rect -1598 -5800 -1498 -5640
rect -1398 -5800 -1378 -5640
rect -3551 -6037 -3534 -5985
rect -3065 -6037 -3050 -5985
rect -2820 -5940 -2580 -5920
rect -3633 -6670 -3610 -6600
rect -3181 -6670 -3162 -6600
rect -3600 -6848 -3400 -6670
rect -3600 -7084 -3520 -6848
rect -2820 -6860 -2800 -5940
rect -2600 -6700 -2580 -5940
rect -2440 -6000 -1378 -5800
rect -2440 -6300 -1498 -6000
rect -1398 -6300 -1378 -6000
rect -2440 -6400 -1378 -6300
rect -2440 -6700 -1498 -6400
rect -1398 -6700 -1378 -6400
rect -2600 -6780 -1378 -6700
rect -1318 -6700 -1298 -5560
rect -1140 -6680 -1088 -6528
rect -682 -4552 -630 -4508
rect -682 -6540 -630 -6528
rect -224 -4552 -172 -4540
rect -224 -6680 -172 -6528
rect 234 -4552 286 -4508
rect 234 -6540 286 -6528
rect 692 -4552 744 -4540
rect 1192 -5540 1244 -5412
rect 1310 -3436 1362 -3424
rect 1310 -5540 1362 -5412
rect 1428 -3436 1480 -3186
rect 1541 -3240 1602 -3231
rect 1541 -3296 1544 -3240
rect 1600 -3296 1602 -3240
rect 1541 -3305 1602 -3296
rect 1428 -5424 1480 -5412
rect 1546 -3436 1598 -3424
rect 692 -6680 744 -6528
rect -1140 -6700 744 -6680
rect 902 -5560 1362 -5540
rect 902 -6700 922 -5560
rect -1318 -6780 922 -6700
rect 982 -5564 1362 -5560
rect 1546 -5564 1598 -5412
rect 1664 -3436 1716 -3186
rect 1664 -5424 1716 -5412
rect 1782 -3436 1834 -3424
rect 1782 -5564 1834 -5412
rect 1900 -3436 1952 -3424
rect 2252 -3770 2402 -3750
rect 2252 -4160 2272 -3770
rect 2382 -4160 2402 -3770
rect 2252 -4180 2402 -4160
rect 2482 -3770 2632 -3750
rect 2482 -4160 2502 -3770
rect 2612 -4160 2632 -3770
rect 2482 -4180 2632 -4160
rect 1900 -5564 1952 -5412
rect 982 -5634 1952 -5564
rect 982 -5640 1402 -5634
rect 982 -5900 1002 -5640
rect 1102 -5800 1202 -5640
rect 1302 -5800 1402 -5640
rect 1502 -5800 1602 -5634
rect 1702 -5800 1802 -5634
rect 1102 -5900 2000 -5800
rect 982 -6000 2000 -5900
rect 982 -6300 1002 -6000
rect 1102 -6300 2000 -6000
rect 982 -6400 2000 -6300
rect 982 -6700 1002 -6400
rect 1102 -6700 2000 -6400
rect 982 -6780 2000 -6700
rect -2600 -6860 2000 -6780
rect -2820 -7000 2000 -6860
rect -2600 -7100 -1200 -7000
rect -2600 -7700 -2500 -7100
rect -1300 -7700 -1200 -7100
rect -2600 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via2 >>
rect -1900 -500 1300 0
rect -1997 -3242 -1941 -3240
rect -1997 -3294 -1995 -3242
rect -1995 -3294 -1943 -3242
rect -1943 -3294 -1941 -3242
rect -1997 -3296 -1941 -3294
rect 1682 -3150 1792 -3060
rect -903 -4200 -837 -4150
rect -903 -4206 -837 -4200
rect -711 -4200 -645 -4150
rect -711 -4206 -645 -4200
rect -519 -4200 -453 -4150
rect -519 -4206 -453 -4200
rect -327 -4200 -261 -4150
rect -327 -4206 -261 -4200
rect -135 -4200 -69 -4150
rect -135 -4206 -69 -4200
rect 57 -4200 123 -4150
rect 57 -4206 123 -4200
rect 249 -4200 315 -4150
rect 249 -4206 315 -4200
rect 441 -4200 507 -4150
rect 441 -4206 507 -4200
rect -1390 -4500 -1230 -4440
rect -3280 -5985 -3070 -5768
rect -3280 -5988 -3070 -5985
rect -2800 -6860 -2600 -5940
rect 1544 -3242 1600 -3240
rect 1544 -3294 1546 -3242
rect 1546 -3294 1598 -3242
rect 1598 -3294 1600 -3242
rect 1544 -3296 1600 -3294
rect 2272 -4160 2382 -3770
rect 2502 -4160 2612 -3770
rect -2500 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< metal3 >>
rect -2000 0 1400 100
rect -7000 -7100 -4200 -200
rect -3800 -5500 -2500 -148
rect -2000 -500 -1900 0
rect 1300 -500 1400 0
rect -2000 -600 1400 -500
rect 1672 -3060 1802 -3050
rect 1672 -3150 1682 -3060
rect 1792 -3150 1802 -3060
rect 2002 -3100 2802 -400
rect 1672 -3160 1802 -3150
rect 2202 -3220 2802 -3100
rect -2005 -3240 2142 -3231
rect -2005 -3296 -1997 -3240
rect -1941 -3296 1544 -3240
rect 1600 -3296 2142 -3240
rect -2005 -3305 2142 -3296
rect -1938 -3336 1541 -3305
rect 2068 -3751 2142 -3305
rect 2202 -3380 2222 -3220
rect 2782 -3380 2802 -3220
rect 2202 -3460 2232 -3380
rect 2772 -3460 2802 -3380
rect 2202 -3490 2802 -3460
rect 2512 -3750 2582 -3490
rect 2252 -3751 2402 -3750
rect 2068 -3770 2402 -3751
rect 2068 -3825 2272 -3770
rect -909 -4150 -255 -4138
rect -909 -4206 -903 -4150
rect -837 -4206 -711 -4150
rect -645 -4206 -519 -4150
rect -453 -4206 -327 -4150
rect -261 -4206 -255 -4150
rect -909 -4220 -255 -4206
rect -141 -4150 513 -4138
rect -141 -4206 -135 -4150
rect -69 -4206 57 -4150
rect 123 -4206 249 -4150
rect 315 -4206 441 -4150
rect 507 -4206 513 -4150
rect 2252 -4160 2272 -3825
rect 2382 -4160 2402 -3770
rect 2252 -4180 2402 -4160
rect 2482 -3770 2632 -3750
rect 2482 -4160 2502 -3770
rect 2612 -4160 2632 -3770
rect 2482 -4180 2632 -4160
rect -141 -4220 513 -4206
rect -1400 -4440 -1220 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1220 -4440
rect -3800 -5700 -2100 -5500
rect -1400 -5700 -1220 -4500
rect -3800 -5748 -2500 -5700
rect -3800 -5768 -2900 -5748
rect -3800 -5988 -3280 -5768
rect -3070 -5988 -2900 -5768
rect -3800 -6248 -2900 -5988
rect -3800 -6648 -3700 -6248
rect -3000 -6648 -2900 -6248
rect -3800 -6748 -2900 -6648
rect -2820 -5940 -2500 -5920
rect -2820 -6860 -2800 -5940
rect -2520 -6860 -2500 -5940
rect -2400 -6000 -1220 -5700
rect -2820 -6880 -2500 -6860
rect -7000 -7700 -6900 -7100
rect -4300 -7700 -4200 -7100
rect -7000 -7800 -4200 -7700
rect -2600 -7100 -1200 -7000
rect -2600 -7700 -2500 -7100
rect -1300 -7700 -1200 -7100
rect -2600 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via3 >>
rect -1900 -500 1300 0
rect 1682 -3150 1792 -3060
rect 2222 -3380 2782 -3220
rect 2232 -3460 2772 -3380
rect -3700 -6648 -3000 -6248
rect -2720 -6860 -2600 -5940
rect -2600 -6860 -2520 -5940
rect -6900 -7700 -4300 -7100
rect -2500 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< mimcap >>
rect -3700 -288 -2600 -248
rect -6900 -340 -4300 -300
rect -6900 -6460 -6860 -340
rect -4340 -6460 -4300 -340
rect -3700 -5608 -3660 -288
rect -2640 -5608 -2600 -288
rect 2032 -450 2772 -430
rect 2032 -3050 2052 -450
rect 2752 -3050 2772 -450
rect 2032 -3070 2772 -3050
rect -3700 -5648 -2600 -5608
rect -6900 -6500 -4300 -6460
<< mimcapcontact >>
rect -6860 -6460 -4340 -340
rect -3660 -5608 -2640 -288
rect 2052 -3050 2752 -450
<< metal4 >>
rect -6800 100 1400 600
rect -6800 -200 -4400 100
rect -2000 0 1400 100
rect -7000 -340 -4200 -200
rect -7000 -6460 -6860 -340
rect -4340 -6460 -4200 -340
rect -3800 -288 -2500 -148
rect -3800 -5608 -3660 -288
rect -2640 -5608 -2500 -288
rect -2000 -500 -1900 0
rect 1300 -500 1400 0
rect -2000 -600 1400 -500
rect 2002 -450 2802 -400
rect 2002 -3040 2052 -450
rect 1672 -3050 2052 -3040
rect 2752 -3050 2802 -450
rect 1672 -3060 2802 -3050
rect 1672 -3150 1682 -3060
rect 1792 -3100 2802 -3060
rect 1792 -3150 1802 -3100
rect 1672 -3160 1802 -3150
rect 2202 -3220 2802 -3200
rect 2202 -3380 2222 -3220
rect 2202 -3460 2232 -3380
rect 2782 -3380 2802 -3220
rect 2772 -3460 2802 -3380
rect 2202 -3490 2802 -3460
rect -3800 -5748 -2500 -5608
rect -2740 -5940 -2500 -5748
rect -7000 -6600 -4200 -6460
rect -3800 -6248 -2900 -6148
rect -3800 -6648 -3700 -6248
rect -3000 -6648 -2900 -6248
rect -3800 -6748 -2900 -6648
rect -2740 -6860 -2720 -5940
rect -2520 -6860 -2500 -5940
rect -2740 -6880 -2500 -6860
rect -2740 -7000 -2501 -6880
rect -7000 -7100 -4200 -7000
rect -7000 -7700 -6900 -7100
rect -4300 -7300 -4200 -7100
rect -2740 -7100 2000 -7000
rect -2740 -7300 -2500 -7100
rect -4300 -7700 -2500 -7300
rect -1300 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect -7000 -7800 2000 -7700
<< via4 >>
rect 2232 -3460 2772 -3220
rect -3700 -6648 -3000 -6248
rect -6900 -7700 -4300 -7100
<< mimcap2 >>
rect -3700 -288 -2600 -248
rect -6900 -340 -4300 -300
rect -6900 -6460 -6860 -340
rect -4340 -6460 -4300 -340
rect -3700 -5608 -3660 -288
rect -2640 -5608 -2600 -288
rect 2032 -450 2772 -430
rect 2032 -3050 2052 -450
rect 2752 -3050 2772 -450
rect 2032 -3070 2772 -3050
rect -3700 -5648 -2600 -5608
rect -6900 -6500 -4300 -6460
<< mimcap2contact >>
rect -6860 -6460 -4340 -340
rect -3660 -5608 -2640 -288
rect 2052 -3050 2752 -450
<< metal5 >>
rect -7000 -340 -4200 -200
rect -7000 -6460 -6860 -340
rect -4340 -6460 -4200 -340
rect -7000 -7100 -4200 -6460
rect -3800 -288 -2500 -148
rect -3800 -5608 -3660 -288
rect -2640 -5608 -2500 -288
rect 2002 -450 2802 -400
rect 2002 -3050 2052 -450
rect 2752 -3050 2802 -450
rect 2002 -3100 2802 -3050
rect 2202 -3220 2802 -3100
rect 2202 -3460 2232 -3220
rect 2772 -3460 2802 -3220
rect 2202 -3490 2802 -3460
rect -3800 -5748 -2500 -5608
rect -3800 -6248 -2900 -5748
rect -3800 -6648 -3700 -6248
rect -3000 -6648 -2900 -6248
rect -3800 -6748 -2900 -6648
rect -7000 -7700 -6900 -7100
rect -4300 -7700 -4200 -7100
rect -7000 -7800 -4200 -7700
<< comment >>
rect -198 -5100 -195 -560
<< labels >>
rlabel metal3 -660 -4200 -620 -4180 1 VIN
rlabel metal3 120 -4200 160 -4180 1 VIP
rlabel metal4 -3820 320 -3440 600 1 VHI
rlabel metal4 -3440 -7800 -3260 -7300 1 VLO
rlabel metal1 -3701 -7084 -3661 -7044 1 SBAR
rlabel metal1 -3769 -7084 -3729 -7044 1 S
rlabel metal2 -3600 -7084 -3520 -7004 1 VREF
rlabel metal3 -2080 -5780 -2020 -5720 1 VREF_GATED
rlabel metal2 1682 -3186 1802 -3134 1 VOP
<< end >>
