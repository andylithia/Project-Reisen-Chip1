magic
tech sky130A
timestamp 1671154469
<< pwell >>
rect -4007 2516 -2880 2976
<< nmoslvt >>
rect -3907 2621 -3892 2871
rect -3859 2621 -3844 2871
rect -3811 2621 -3796 2871
rect -3763 2621 -3748 2871
rect -3715 2621 -3700 2871
rect -3667 2621 -3652 2871
rect -3619 2621 -3604 2871
rect -3571 2621 -3556 2871
rect -3523 2621 -3508 2871
rect -3475 2621 -3460 2871
rect -3427 2621 -3412 2871
rect -3379 2621 -3364 2871
rect -3331 2621 -3316 2871
rect -3283 2621 -3268 2871
rect -3235 2621 -3220 2871
rect -3187 2621 -3172 2871
rect -3139 2621 -3124 2871
rect -3091 2621 -3076 2871
rect -3043 2621 -3028 2871
rect -2995 2621 -2980 2871
<< ndiff >>
rect -3938 2865 -3907 2871
rect -3938 2627 -3932 2865
rect -3915 2627 -3907 2865
rect -3938 2621 -3907 2627
rect -3892 2865 -3859 2871
rect -3892 2627 -3884 2865
rect -3867 2627 -3859 2865
rect -3892 2621 -3859 2627
rect -3844 2865 -3811 2871
rect -3844 2627 -3836 2865
rect -3819 2627 -3811 2865
rect -3844 2621 -3811 2627
rect -3796 2865 -3763 2871
rect -3796 2627 -3788 2865
rect -3771 2627 -3763 2865
rect -3796 2621 -3763 2627
rect -3748 2865 -3715 2871
rect -3748 2627 -3740 2865
rect -3723 2627 -3715 2865
rect -3748 2621 -3715 2627
rect -3700 2865 -3667 2871
rect -3700 2627 -3692 2865
rect -3675 2627 -3667 2865
rect -3700 2621 -3667 2627
rect -3652 2865 -3619 2871
rect -3652 2627 -3644 2865
rect -3627 2627 -3619 2865
rect -3652 2621 -3619 2627
rect -3604 2865 -3571 2871
rect -3604 2627 -3596 2865
rect -3579 2627 -3571 2865
rect -3604 2621 -3571 2627
rect -3556 2865 -3523 2871
rect -3556 2627 -3548 2865
rect -3531 2627 -3523 2865
rect -3556 2621 -3523 2627
rect -3508 2865 -3475 2871
rect -3508 2627 -3500 2865
rect -3483 2627 -3475 2865
rect -3508 2621 -3475 2627
rect -3460 2865 -3427 2871
rect -3460 2627 -3452 2865
rect -3435 2627 -3427 2865
rect -3460 2621 -3427 2627
rect -3412 2865 -3379 2871
rect -3412 2627 -3404 2865
rect -3387 2627 -3379 2865
rect -3412 2621 -3379 2627
rect -3364 2865 -3331 2871
rect -3364 2627 -3356 2865
rect -3339 2627 -3331 2865
rect -3364 2621 -3331 2627
rect -3316 2865 -3283 2871
rect -3316 2627 -3308 2865
rect -3291 2627 -3283 2865
rect -3316 2621 -3283 2627
rect -3268 2865 -3235 2871
rect -3268 2627 -3260 2865
rect -3243 2627 -3235 2865
rect -3268 2621 -3235 2627
rect -3220 2865 -3187 2871
rect -3220 2627 -3212 2865
rect -3195 2627 -3187 2865
rect -3220 2621 -3187 2627
rect -3172 2865 -3139 2871
rect -3172 2627 -3164 2865
rect -3147 2627 -3139 2865
rect -3172 2621 -3139 2627
rect -3124 2865 -3091 2871
rect -3124 2627 -3116 2865
rect -3099 2627 -3091 2865
rect -3124 2621 -3091 2627
rect -3076 2865 -3043 2871
rect -3076 2627 -3068 2865
rect -3051 2627 -3043 2865
rect -3076 2621 -3043 2627
rect -3028 2865 -2995 2871
rect -3028 2627 -3020 2865
rect -3003 2627 -2995 2865
rect -3028 2621 -2995 2627
rect -2980 2865 -2949 2871
rect -2980 2627 -2972 2865
rect -2955 2627 -2949 2865
rect -2980 2621 -2949 2627
<< ndiffc >>
rect -3932 2627 -3915 2865
rect -3884 2627 -3867 2865
rect -3836 2627 -3819 2865
rect -3788 2627 -3771 2865
rect -3740 2627 -3723 2865
rect -3692 2627 -3675 2865
rect -3644 2627 -3627 2865
rect -3596 2627 -3579 2865
rect -3548 2627 -3531 2865
rect -3500 2627 -3483 2865
rect -3452 2627 -3435 2865
rect -3404 2627 -3387 2865
rect -3356 2627 -3339 2865
rect -3308 2627 -3291 2865
rect -3260 2627 -3243 2865
rect -3212 2627 -3195 2865
rect -3164 2627 -3147 2865
rect -3116 2627 -3099 2865
rect -3068 2627 -3051 2865
rect -3020 2627 -3003 2865
rect -2972 2627 -2955 2865
<< psubdiff >>
rect -3989 2941 -3941 2958
rect -2946 2941 -2898 2958
rect -3989 2910 -3972 2941
rect -2915 2910 -2898 2941
rect -3989 2551 -3972 2582
rect -2915 2551 -2898 2582
rect -3989 2534 -3941 2551
rect -2946 2534 -2898 2551
<< psubdiffcont >>
rect -3941 2941 -2946 2958
rect -3989 2582 -3972 2910
rect -2915 2582 -2898 2910
rect -3941 2534 -2946 2551
<< poly >>
rect -3811 2913 -3748 2921
rect -3811 2896 -3788 2913
rect -3771 2896 -3748 2913
rect -3907 2871 -3892 2884
rect -3859 2871 -3844 2884
rect -3811 2882 -3748 2896
rect -3811 2871 -3796 2882
rect -3763 2871 -3748 2882
rect -3715 2913 -3652 2921
rect -3715 2896 -3692 2913
rect -3675 2896 -3652 2913
rect -3715 2882 -3652 2896
rect -3715 2871 -3700 2882
rect -3667 2871 -3652 2882
rect -3619 2913 -3556 2921
rect -3619 2896 -3596 2913
rect -3579 2896 -3556 2913
rect -3619 2882 -3556 2896
rect -3619 2871 -3604 2882
rect -3571 2871 -3556 2882
rect -3523 2913 -3460 2921
rect -3523 2896 -3500 2913
rect -3483 2896 -3460 2913
rect -3523 2882 -3460 2896
rect -3523 2871 -3508 2882
rect -3475 2871 -3460 2882
rect -3427 2913 -3364 2921
rect -3427 2896 -3404 2913
rect -3387 2896 -3364 2913
rect -3427 2882 -3364 2896
rect -3427 2871 -3412 2882
rect -3379 2871 -3364 2882
rect -3331 2913 -3268 2921
rect -3331 2896 -3308 2913
rect -3291 2896 -3268 2913
rect -3331 2882 -3268 2896
rect -3331 2871 -3316 2882
rect -3283 2871 -3268 2882
rect -3235 2913 -3172 2921
rect -3235 2896 -3212 2913
rect -3195 2896 -3172 2913
rect -3235 2882 -3172 2896
rect -3235 2871 -3220 2882
rect -3187 2871 -3172 2882
rect -3139 2913 -3076 2921
rect -3139 2896 -3116 2913
rect -3099 2896 -3076 2913
rect -3139 2882 -3076 2896
rect -3139 2871 -3124 2882
rect -3091 2871 -3076 2882
rect -3043 2871 -3028 2884
rect -2995 2871 -2980 2884
rect -3907 2608 -3892 2621
rect -3859 2608 -3844 2621
rect -3811 2608 -3796 2621
rect -3763 2608 -3748 2621
rect -3715 2608 -3700 2621
rect -3667 2608 -3652 2621
rect -3619 2608 -3604 2621
rect -3571 2608 -3556 2621
rect -3523 2608 -3508 2621
rect -3475 2608 -3460 2621
rect -3427 2608 -3412 2621
rect -3379 2608 -3364 2621
rect -3331 2608 -3316 2621
rect -3283 2608 -3268 2621
rect -3235 2608 -3220 2621
rect -3187 2608 -3172 2621
rect -3139 2608 -3124 2621
rect -3091 2608 -3076 2621
rect -3043 2608 -3028 2621
rect -2995 2608 -2980 2621
rect -3907 2600 -3844 2608
rect -3907 2583 -3884 2600
rect -3867 2583 -3844 2600
rect -3907 2569 -3844 2583
rect -3043 2600 -2980 2608
rect -3043 2583 -3020 2600
rect -3003 2583 -2980 2600
rect -3043 2569 -2980 2583
<< polycont >>
rect -3788 2896 -3771 2913
rect -3692 2896 -3675 2913
rect -3596 2896 -3579 2913
rect -3500 2896 -3483 2913
rect -3404 2896 -3387 2913
rect -3308 2896 -3291 2913
rect -3212 2896 -3195 2913
rect -3116 2896 -3099 2913
rect -3884 2583 -3867 2600
rect -3020 2583 -3003 2600
<< locali >>
rect -3989 2941 -3941 2958
rect -2946 2941 -2898 2958
rect -3989 2910 -3972 2941
rect -3796 2896 -3788 2913
rect -3771 2896 -3763 2913
rect -3700 2896 -3692 2913
rect -3675 2896 -3667 2913
rect -3604 2896 -3596 2913
rect -3579 2896 -3571 2913
rect -3508 2896 -3500 2913
rect -3483 2896 -3475 2913
rect -3412 2896 -3404 2913
rect -3387 2896 -3379 2913
rect -3316 2896 -3308 2913
rect -3291 2896 -3283 2913
rect -3220 2896 -3212 2913
rect -3195 2896 -3187 2913
rect -3124 2896 -3116 2913
rect -3099 2896 -3091 2913
rect -2915 2910 -2898 2941
rect -3932 2865 -3915 2873
rect -3932 2619 -3915 2627
rect -3884 2865 -3867 2873
rect -3884 2619 -3867 2627
rect -3836 2865 -3819 2873
rect -3836 2619 -3819 2627
rect -3788 2865 -3771 2873
rect -3788 2619 -3771 2627
rect -3740 2865 -3723 2873
rect -3740 2619 -3723 2627
rect -3692 2865 -3675 2873
rect -3692 2619 -3675 2627
rect -3644 2865 -3627 2873
rect -3644 2619 -3627 2627
rect -3596 2865 -3579 2873
rect -3596 2619 -3579 2627
rect -3548 2865 -3531 2873
rect -3548 2619 -3531 2627
rect -3500 2865 -3483 2873
rect -3500 2619 -3483 2627
rect -3452 2865 -3435 2873
rect -3452 2619 -3435 2627
rect -3404 2865 -3387 2873
rect -3404 2619 -3387 2627
rect -3356 2865 -3339 2873
rect -3356 2619 -3339 2627
rect -3308 2865 -3291 2873
rect -3308 2619 -3291 2627
rect -3260 2865 -3243 2873
rect -3260 2619 -3243 2627
rect -3212 2865 -3195 2873
rect -3212 2619 -3195 2627
rect -3164 2865 -3147 2873
rect -3164 2619 -3147 2627
rect -3116 2865 -3099 2873
rect -3116 2619 -3099 2627
rect -3068 2865 -3051 2873
rect -3068 2619 -3051 2627
rect -3020 2865 -3003 2873
rect -3020 2619 -3003 2627
rect -2972 2865 -2955 2873
rect -2972 2619 -2955 2627
rect -3892 2583 -3884 2600
rect -3867 2583 -3859 2600
rect -3028 2583 -3020 2600
rect -3003 2583 -2995 2600
rect -3989 2551 -3972 2582
rect -2915 2551 -2898 2582
rect -3989 2534 -3941 2551
rect -2946 2534 -2898 2551
<< viali >>
rect -3788 2896 -3771 2913
rect -3692 2896 -3675 2913
rect -3596 2896 -3579 2913
rect -3500 2896 -3483 2913
rect -3404 2896 -3387 2913
rect -3308 2896 -3291 2913
rect -3212 2896 -3195 2913
rect -3116 2896 -3099 2913
rect -3989 2621 -3972 2871
rect -3932 2627 -3915 2865
rect -3884 2627 -3867 2865
rect -3836 2627 -3819 2865
rect -3788 2627 -3771 2865
rect -3740 2627 -3723 2865
rect -3692 2627 -3675 2865
rect -3644 2627 -3627 2865
rect -3596 2627 -3579 2865
rect -3548 2627 -3531 2865
rect -3500 2627 -3483 2865
rect -3452 2627 -3435 2865
rect -3404 2627 -3387 2865
rect -3356 2627 -3339 2865
rect -3308 2627 -3291 2865
rect -3260 2627 -3243 2865
rect -3212 2627 -3195 2865
rect -3164 2627 -3147 2865
rect -3116 2627 -3099 2865
rect -3068 2627 -3051 2865
rect -3020 2627 -3003 2865
rect -2972 2627 -2955 2865
rect -2915 2621 -2898 2871
rect -3884 2583 -3867 2600
rect -3020 2583 -3003 2600
<< metal1 >>
rect -3799 2893 -3796 2921
rect -3763 2893 -3760 2921
rect -3703 2893 -3700 2921
rect -3667 2893 -3664 2921
rect -3607 2893 -3604 2921
rect -3571 2893 -3568 2921
rect -3511 2893 -3508 2921
rect -3475 2893 -3472 2921
rect -3415 2893 -3412 2921
rect -3379 2893 -3376 2921
rect -3319 2893 -3316 2921
rect -3283 2893 -3280 2921
rect -3223 2893 -3220 2921
rect -3187 2893 -3184 2921
rect -3127 2893 -3124 2921
rect -3091 2893 -3088 2921
rect -3992 2871 -3969 2877
rect -2918 2871 -2895 2877
rect -3992 2621 -3989 2871
rect -3972 2621 -3937 2871
rect -3910 2621 -3907 2871
rect -3892 2621 -3889 2871
rect -3862 2621 -3859 2871
rect -3844 2621 -3841 2871
rect -3814 2621 -3811 2871
rect -3796 2621 -3793 2871
rect -3766 2621 -3763 2871
rect -3748 2621 -3745 2871
rect -3718 2621 -3715 2871
rect -3700 2621 -3697 2871
rect -3670 2621 -3667 2871
rect -3652 2621 -3649 2871
rect -3622 2621 -3619 2871
rect -3604 2621 -3601 2871
rect -3574 2621 -3571 2871
rect -3556 2621 -3553 2871
rect -3526 2621 -3523 2871
rect -3508 2621 -3505 2871
rect -3478 2621 -3475 2871
rect -3460 2621 -3457 2871
rect -3430 2621 -3427 2871
rect -3412 2621 -3409 2871
rect -3382 2621 -3379 2871
rect -3364 2621 -3361 2871
rect -3334 2621 -3331 2871
rect -3316 2621 -3313 2871
rect -3286 2621 -3283 2871
rect -3268 2621 -3265 2871
rect -3238 2621 -3235 2871
rect -3220 2621 -3217 2871
rect -3190 2621 -3187 2871
rect -3172 2621 -3169 2871
rect -3142 2621 -3139 2871
rect -3124 2621 -3121 2871
rect -3094 2621 -3091 2871
rect -3076 2621 -3073 2871
rect -3046 2621 -3043 2871
rect -3028 2621 -3025 2871
rect -2998 2621 -2995 2871
rect -2980 2621 -2977 2871
rect -2950 2621 -2915 2871
rect -2898 2621 -2895 2871
rect -3992 2615 -3969 2621
rect -3935 2603 -3912 2621
rect -3887 2603 -3864 2621
rect -3023 2603 -3000 2621
rect -2975 2603 -2952 2621
rect -2918 2615 -2895 2621
rect -3935 2600 -3859 2603
rect -3935 2583 -3884 2600
rect -3867 2583 -3859 2600
rect -3935 2580 -3859 2583
rect -3028 2600 -2952 2603
rect -3028 2583 -3020 2600
rect -3003 2583 -2952 2600
rect -3028 2580 -2952 2583
<< via1 >>
rect -3796 2913 -3763 2921
rect -3796 2896 -3788 2913
rect -3788 2896 -3771 2913
rect -3771 2896 -3763 2913
rect -3796 2893 -3763 2896
rect -3700 2913 -3667 2921
rect -3700 2896 -3692 2913
rect -3692 2896 -3675 2913
rect -3675 2896 -3667 2913
rect -3700 2893 -3667 2896
rect -3604 2913 -3571 2921
rect -3604 2896 -3596 2913
rect -3596 2896 -3579 2913
rect -3579 2896 -3571 2913
rect -3604 2893 -3571 2896
rect -3508 2913 -3475 2921
rect -3508 2896 -3500 2913
rect -3500 2896 -3483 2913
rect -3483 2896 -3475 2913
rect -3508 2893 -3475 2896
rect -3412 2913 -3379 2921
rect -3412 2896 -3404 2913
rect -3404 2896 -3387 2913
rect -3387 2896 -3379 2913
rect -3412 2893 -3379 2896
rect -3316 2913 -3283 2921
rect -3316 2896 -3308 2913
rect -3308 2896 -3291 2913
rect -3291 2896 -3283 2913
rect -3316 2893 -3283 2896
rect -3220 2913 -3187 2921
rect -3220 2896 -3212 2913
rect -3212 2896 -3195 2913
rect -3195 2896 -3187 2913
rect -3220 2893 -3187 2896
rect -3124 2913 -3091 2921
rect -3124 2896 -3116 2913
rect -3116 2896 -3099 2913
rect -3099 2896 -3091 2913
rect -3124 2893 -3091 2896
rect -3937 2865 -3910 2871
rect -3937 2627 -3932 2865
rect -3932 2627 -3915 2865
rect -3915 2627 -3910 2865
rect -3937 2621 -3910 2627
rect -3889 2865 -3862 2871
rect -3889 2627 -3884 2865
rect -3884 2627 -3867 2865
rect -3867 2627 -3862 2865
rect -3889 2621 -3862 2627
rect -3841 2865 -3814 2871
rect -3841 2627 -3836 2865
rect -3836 2627 -3819 2865
rect -3819 2627 -3814 2865
rect -3841 2621 -3814 2627
rect -3793 2865 -3766 2871
rect -3793 2627 -3788 2865
rect -3788 2627 -3771 2865
rect -3771 2627 -3766 2865
rect -3793 2621 -3766 2627
rect -3745 2865 -3718 2871
rect -3745 2627 -3740 2865
rect -3740 2627 -3723 2865
rect -3723 2627 -3718 2865
rect -3745 2621 -3718 2627
rect -3697 2865 -3670 2871
rect -3697 2627 -3692 2865
rect -3692 2627 -3675 2865
rect -3675 2627 -3670 2865
rect -3697 2621 -3670 2627
rect -3649 2865 -3622 2871
rect -3649 2627 -3644 2865
rect -3644 2627 -3627 2865
rect -3627 2627 -3622 2865
rect -3649 2621 -3622 2627
rect -3601 2865 -3574 2871
rect -3601 2627 -3596 2865
rect -3596 2627 -3579 2865
rect -3579 2627 -3574 2865
rect -3601 2621 -3574 2627
rect -3553 2865 -3526 2871
rect -3553 2627 -3548 2865
rect -3548 2627 -3531 2865
rect -3531 2627 -3526 2865
rect -3553 2621 -3526 2627
rect -3505 2865 -3478 2871
rect -3505 2627 -3500 2865
rect -3500 2627 -3483 2865
rect -3483 2627 -3478 2865
rect -3505 2621 -3478 2627
rect -3457 2865 -3430 2871
rect -3457 2627 -3452 2865
rect -3452 2627 -3435 2865
rect -3435 2627 -3430 2865
rect -3457 2621 -3430 2627
rect -3409 2865 -3382 2871
rect -3409 2627 -3404 2865
rect -3404 2627 -3387 2865
rect -3387 2627 -3382 2865
rect -3409 2621 -3382 2627
rect -3361 2865 -3334 2871
rect -3361 2627 -3356 2865
rect -3356 2627 -3339 2865
rect -3339 2627 -3334 2865
rect -3361 2621 -3334 2627
rect -3313 2865 -3286 2871
rect -3313 2627 -3308 2865
rect -3308 2627 -3291 2865
rect -3291 2627 -3286 2865
rect -3313 2621 -3286 2627
rect -3265 2865 -3238 2871
rect -3265 2627 -3260 2865
rect -3260 2627 -3243 2865
rect -3243 2627 -3238 2865
rect -3265 2621 -3238 2627
rect -3217 2865 -3190 2871
rect -3217 2627 -3212 2865
rect -3212 2627 -3195 2865
rect -3195 2627 -3190 2865
rect -3217 2621 -3190 2627
rect -3169 2865 -3142 2871
rect -3169 2627 -3164 2865
rect -3164 2627 -3147 2865
rect -3147 2627 -3142 2865
rect -3169 2621 -3142 2627
rect -3121 2865 -3094 2871
rect -3121 2627 -3116 2865
rect -3116 2627 -3099 2865
rect -3099 2627 -3094 2865
rect -3121 2621 -3094 2627
rect -3073 2865 -3046 2871
rect -3073 2627 -3068 2865
rect -3068 2627 -3051 2865
rect -3051 2627 -3046 2865
rect -3073 2621 -3046 2627
rect -3025 2865 -2998 2871
rect -3025 2627 -3020 2865
rect -3020 2627 -3003 2865
rect -3003 2627 -2998 2865
rect -3025 2621 -2998 2627
rect -2977 2865 -2950 2871
rect -2977 2627 -2972 2865
rect -2972 2627 -2955 2865
rect -2955 2627 -2950 2865
rect -2977 2621 -2950 2627
<< metal2 >>
rect -3841 2951 -3046 2986
rect -3841 2871 -3814 2951
rect -3796 2924 -3763 2931
rect -3796 2890 -3763 2893
rect -3745 2871 -3718 2951
rect -3700 2924 -3667 2931
rect -3700 2890 -3667 2893
rect -3649 2871 -3622 2951
rect -3604 2924 -3571 2931
rect -3604 2890 -3571 2893
rect -3553 2871 -3526 2951
rect -3508 2924 -3475 2931
rect -3508 2890 -3475 2893
rect -3457 2871 -3430 2951
rect -3412 2924 -3379 2931
rect -3412 2890 -3379 2893
rect -3361 2871 -3334 2951
rect -3316 2924 -3283 2931
rect -3316 2890 -3283 2893
rect -3265 2871 -3238 2951
rect -3220 2924 -3187 2931
rect -3220 2890 -3187 2893
rect -3169 2871 -3142 2951
rect -3124 2924 -3091 2931
rect -3124 2890 -3091 2893
rect -3073 2871 -3046 2951
rect -3940 2621 -3937 2871
rect -3910 2621 -3907 2871
rect -3892 2621 -3889 2871
rect -3862 2621 -3859 2871
rect -3844 2621 -3841 2871
rect -3814 2621 -3811 2871
rect -3796 2621 -3793 2871
rect -3766 2621 -3763 2871
rect -3748 2621 -3745 2871
rect -3718 2621 -3715 2871
rect -3700 2621 -3697 2871
rect -3670 2621 -3667 2871
rect -3652 2621 -3649 2871
rect -3622 2621 -3619 2871
rect -3604 2621 -3601 2871
rect -3574 2621 -3571 2871
rect -3556 2621 -3553 2871
rect -3526 2621 -3523 2871
rect -3508 2621 -3505 2871
rect -3478 2621 -3475 2871
rect -3460 2621 -3457 2871
rect -3430 2621 -3427 2871
rect -3412 2621 -3409 2871
rect -3382 2621 -3379 2871
rect -3364 2621 -3361 2871
rect -3334 2621 -3331 2871
rect -3316 2621 -3313 2871
rect -3286 2621 -3283 2871
rect -3268 2621 -3265 2871
rect -3238 2621 -3235 2871
rect -3220 2621 -3217 2871
rect -3190 2621 -3187 2871
rect -3172 2621 -3169 2871
rect -3142 2621 -3139 2871
rect -3124 2621 -3121 2871
rect -3094 2621 -3091 2871
rect -3076 2621 -3073 2871
rect -3046 2621 -3043 2871
rect -3028 2621 -3025 2871
rect -2998 2621 -2995 2871
rect -2980 2621 -2977 2871
rect -2950 2621 -2947 2871
rect -3796 2586 -3763 2621
rect -3700 2586 -3667 2621
rect -3604 2586 -3571 2621
rect -3508 2586 -3475 2621
rect -3796 2516 -3475 2586
rect -3412 2586 -3379 2621
rect -3316 2586 -3283 2621
rect -3220 2586 -3187 2621
rect -3124 2586 -3091 2621
rect -3412 2516 -3091 2586
<< via2 >>
rect -3796 2921 -3763 2924
rect -3796 2896 -3763 2921
rect -3700 2921 -3667 2924
rect -3700 2896 -3667 2921
rect -3604 2921 -3571 2924
rect -3604 2896 -3571 2921
rect -3508 2921 -3475 2924
rect -3508 2896 -3475 2921
rect -3412 2921 -3379 2924
rect -3412 2896 -3379 2921
rect -3316 2921 -3283 2924
rect -3316 2896 -3283 2921
rect -3220 2921 -3187 2924
rect -3220 2896 -3187 2921
rect -3124 2921 -3091 2924
rect -3124 2896 -3091 2921
<< metal3 >>
rect -3799 2924 -3472 2931
rect -3799 2896 -3796 2924
rect -3763 2896 -3700 2924
rect -3667 2896 -3604 2924
rect -3571 2896 -3508 2924
rect -3475 2896 -3472 2924
rect -3799 2890 -3472 2896
rect -3415 2924 -3088 2931
rect -3415 2896 -3412 2924
rect -3379 2896 -3316 2924
rect -3283 2896 -3220 2924
rect -3187 2896 -3124 2924
rect -3091 2896 -3088 2924
rect -3415 2890 -3088 2896
<< labels >>
rlabel metal2 -3841 2977 -3800 2986 1 CS
rlabel metal3 -3761 2923 -3747 2931 1 G1
rlabel metal3 -3331 2923 -3317 2931 1 G2
rlabel metal2 -3796 2516 -3782 2524 1 D1
rlabel metal2 -3412 2516 -3398 2524 1 D2
rlabel metal1 -3935 2580 -3912 2603 1 GND
<< end >>
