magic
tech sky130A
magscale 1 2
timestamp 1672341527
<< locali >>
rect 45140 16699 45260 16750
rect 45140 16665 45183 16699
rect 45217 16665 45260 16699
rect 45140 16627 45260 16665
rect 45140 16593 45183 16627
rect 45217 16593 45260 16627
rect 45140 16555 45260 16593
rect 45140 16521 45183 16555
rect 45217 16521 45260 16555
rect 45140 16483 45260 16521
rect 45140 16449 45183 16483
rect 45217 16449 45260 16483
rect 45140 16411 45260 16449
rect 45140 16377 45183 16411
rect 45217 16377 45260 16411
rect 45140 16339 45260 16377
rect 45140 16305 45183 16339
rect 45217 16305 45260 16339
rect 45140 16267 45260 16305
rect 45140 16233 45183 16267
rect 45217 16233 45260 16267
rect 45140 16195 45260 16233
rect 45140 16161 45183 16195
rect 45217 16161 45260 16195
rect 45140 16123 45260 16161
rect 45140 16089 45183 16123
rect 45217 16089 45260 16123
rect 45140 16051 45260 16089
rect 45140 16017 45183 16051
rect 45217 16017 45260 16051
rect 45140 15979 45260 16017
rect 45140 15945 45183 15979
rect 45217 15945 45260 15979
rect 45140 15907 45260 15945
rect 45140 15873 45183 15907
rect 45217 15873 45260 15907
rect 45140 15835 45260 15873
rect 45140 15801 45183 15835
rect 45217 15801 45260 15835
rect 45140 15750 45260 15801
<< viali >>
rect 45183 16665 45217 16699
rect 45183 16593 45217 16627
rect 45183 16521 45217 16555
rect 45183 16449 45217 16483
rect 45183 16377 45217 16411
rect 45183 16305 45217 16339
rect 45183 16233 45217 16267
rect 45183 16161 45217 16195
rect 45183 16089 45217 16123
rect 45183 16017 45217 16051
rect 45183 15945 45217 15979
rect 45183 15873 45217 15907
rect 45183 15801 45217 15835
<< metal1 >>
rect 45360 26406 45440 26440
rect 45360 26354 45374 26406
rect 45426 26354 45440 26406
rect 45360 26342 45440 26354
rect 45360 26290 45374 26342
rect 45426 26290 45440 26342
rect 45360 26278 45440 26290
rect 45360 26226 45374 26278
rect 45426 26226 45440 26278
rect 45360 26214 45440 26226
rect 45360 26162 45374 26214
rect 45426 26162 45440 26214
rect 45360 26150 45440 26162
rect 45360 26098 45374 26150
rect 45426 26098 45440 26150
rect 45360 26086 45440 26098
rect 45360 26034 45374 26086
rect 45426 26034 45440 26086
rect 45360 26000 45440 26034
rect 45140 16724 45260 16750
rect 45140 16672 45174 16724
rect 45226 16672 45260 16724
rect 45140 16665 45183 16672
rect 45217 16665 45260 16672
rect 45140 16660 45260 16665
rect 45140 16608 45174 16660
rect 45226 16608 45260 16660
rect 45140 16596 45183 16608
rect 45217 16596 45260 16608
rect 45140 16544 45174 16596
rect 45226 16544 45260 16596
rect 45140 16532 45183 16544
rect 45217 16532 45260 16544
rect 45140 16480 45174 16532
rect 45226 16480 45260 16532
rect 45140 16468 45183 16480
rect 45217 16468 45260 16480
rect 45140 16416 45174 16468
rect 45226 16416 45260 16468
rect 45140 16411 45260 16416
rect 45140 16404 45183 16411
rect 45217 16404 45260 16411
rect 45140 16352 45174 16404
rect 45226 16352 45260 16404
rect 45140 16340 45260 16352
rect 45140 16288 45174 16340
rect 45226 16288 45260 16340
rect 45140 16276 45260 16288
rect 45140 16224 45174 16276
rect 45226 16224 45260 16276
rect 45140 16212 45260 16224
rect 45140 16160 45174 16212
rect 45226 16160 45260 16212
rect 45140 16148 45260 16160
rect 45140 16096 45174 16148
rect 45226 16096 45260 16148
rect 45140 16089 45183 16096
rect 45217 16089 45260 16096
rect 45140 16084 45260 16089
rect 45140 16032 45174 16084
rect 45226 16032 45260 16084
rect 45140 16020 45183 16032
rect 45217 16020 45260 16032
rect 45140 15968 45174 16020
rect 45226 15968 45260 16020
rect 45140 15956 45183 15968
rect 45217 15956 45260 15968
rect 45140 15904 45174 15956
rect 45226 15904 45260 15956
rect 45140 15892 45183 15904
rect 45217 15892 45260 15904
rect 45140 15840 45174 15892
rect 45226 15840 45260 15892
rect 45140 15835 45260 15840
rect 45140 15828 45183 15835
rect 45217 15828 45260 15835
rect 45140 15776 45174 15828
rect 45226 15776 45260 15828
rect 45140 15750 45260 15776
rect 45360 5966 45440 6000
rect 45360 5914 45374 5966
rect 45426 5914 45440 5966
rect 45360 5902 45440 5914
rect 45360 5850 45374 5902
rect 45426 5850 45440 5902
rect 45360 5838 45440 5850
rect 45360 5786 45374 5838
rect 45426 5786 45440 5838
rect 45360 5774 45440 5786
rect 45360 5722 45374 5774
rect 45426 5722 45440 5774
rect 45360 5710 45440 5722
rect 45360 5658 45374 5710
rect 45426 5658 45440 5710
rect 45360 5646 45440 5658
rect 45360 5594 45374 5646
rect 45426 5594 45440 5646
rect 45360 5560 45440 5594
<< via1 >>
rect 45374 26354 45426 26406
rect 45374 26290 45426 26342
rect 45374 26226 45426 26278
rect 45374 26162 45426 26214
rect 45374 26098 45426 26150
rect 45374 26034 45426 26086
rect 45174 16699 45226 16724
rect 45174 16672 45183 16699
rect 45183 16672 45217 16699
rect 45217 16672 45226 16699
rect 45174 16627 45226 16660
rect 45174 16608 45183 16627
rect 45183 16608 45217 16627
rect 45217 16608 45226 16627
rect 45174 16593 45183 16596
rect 45183 16593 45217 16596
rect 45217 16593 45226 16596
rect 45174 16555 45226 16593
rect 45174 16544 45183 16555
rect 45183 16544 45217 16555
rect 45217 16544 45226 16555
rect 45174 16521 45183 16532
rect 45183 16521 45217 16532
rect 45217 16521 45226 16532
rect 45174 16483 45226 16521
rect 45174 16480 45183 16483
rect 45183 16480 45217 16483
rect 45217 16480 45226 16483
rect 45174 16449 45183 16468
rect 45183 16449 45217 16468
rect 45217 16449 45226 16468
rect 45174 16416 45226 16449
rect 45174 16377 45183 16404
rect 45183 16377 45217 16404
rect 45217 16377 45226 16404
rect 45174 16352 45226 16377
rect 45174 16339 45226 16340
rect 45174 16305 45183 16339
rect 45183 16305 45217 16339
rect 45217 16305 45226 16339
rect 45174 16288 45226 16305
rect 45174 16267 45226 16276
rect 45174 16233 45183 16267
rect 45183 16233 45217 16267
rect 45217 16233 45226 16267
rect 45174 16224 45226 16233
rect 45174 16195 45226 16212
rect 45174 16161 45183 16195
rect 45183 16161 45217 16195
rect 45217 16161 45226 16195
rect 45174 16160 45226 16161
rect 45174 16123 45226 16148
rect 45174 16096 45183 16123
rect 45183 16096 45217 16123
rect 45217 16096 45226 16123
rect 45174 16051 45226 16084
rect 45174 16032 45183 16051
rect 45183 16032 45217 16051
rect 45217 16032 45226 16051
rect 45174 16017 45183 16020
rect 45183 16017 45217 16020
rect 45217 16017 45226 16020
rect 45174 15979 45226 16017
rect 45174 15968 45183 15979
rect 45183 15968 45217 15979
rect 45217 15968 45226 15979
rect 45174 15945 45183 15956
rect 45183 15945 45217 15956
rect 45217 15945 45226 15956
rect 45174 15907 45226 15945
rect 45174 15904 45183 15907
rect 45183 15904 45217 15907
rect 45217 15904 45226 15907
rect 45174 15873 45183 15892
rect 45183 15873 45217 15892
rect 45217 15873 45226 15892
rect 45174 15840 45226 15873
rect 45174 15801 45183 15828
rect 45183 15801 45217 15828
rect 45217 15801 45226 15828
rect 45174 15776 45226 15801
rect 45374 5914 45426 5966
rect 45374 5850 45426 5902
rect 45374 5786 45426 5838
rect 45374 5722 45426 5774
rect 45374 5658 45426 5710
rect 45374 5594 45426 5646
<< metal2 >>
rect 45330 26408 45470 26440
rect 45330 26352 45372 26408
rect 45428 26352 45470 26408
rect 45330 26342 45470 26352
rect 45330 26328 45374 26342
rect 45426 26328 45470 26342
rect 45330 26272 45372 26328
rect 45428 26272 45470 26328
rect 45330 26248 45374 26272
rect 45426 26248 45470 26272
rect 45330 26192 45372 26248
rect 45428 26192 45470 26248
rect 45330 26168 45374 26192
rect 45426 26168 45470 26192
rect 45330 26112 45372 26168
rect 45428 26112 45470 26168
rect 45330 26098 45374 26112
rect 45426 26098 45470 26112
rect 45330 26088 45470 26098
rect 45330 26032 45372 26088
rect 45428 26032 45470 26088
rect 45330 26000 45470 26032
rect 45140 16724 45260 16750
rect 45140 16718 45174 16724
rect 45226 16718 45260 16724
rect 45140 16662 45172 16718
rect 45228 16662 45260 16718
rect 45140 16660 45260 16662
rect 45140 16638 45174 16660
rect 45226 16638 45260 16660
rect 45140 16582 45172 16638
rect 45228 16582 45260 16638
rect 45140 16558 45174 16582
rect 45226 16558 45260 16582
rect 45140 16502 45172 16558
rect 45228 16502 45260 16558
rect 45140 16480 45174 16502
rect 45226 16480 45260 16502
rect 45140 16478 45260 16480
rect 45140 16422 45172 16478
rect 45228 16422 45260 16478
rect 45140 16416 45174 16422
rect 45226 16416 45260 16422
rect 45140 16404 45260 16416
rect 45140 16398 45174 16404
rect 45226 16398 45260 16404
rect 45140 16342 45172 16398
rect 45228 16342 45260 16398
rect 45140 16340 45260 16342
rect 45140 16318 45174 16340
rect 45226 16318 45260 16340
rect 45140 16262 45172 16318
rect 45228 16262 45260 16318
rect 45140 16238 45174 16262
rect 45226 16238 45260 16262
rect 45140 16182 45172 16238
rect 45228 16182 45260 16238
rect 45140 16160 45174 16182
rect 45226 16160 45260 16182
rect 45140 16158 45260 16160
rect 45140 16102 45172 16158
rect 45228 16102 45260 16158
rect 45140 16096 45174 16102
rect 45226 16096 45260 16102
rect 45140 16084 45260 16096
rect 45140 16078 45174 16084
rect 45226 16078 45260 16084
rect 45140 16022 45172 16078
rect 45228 16022 45260 16078
rect 45140 16020 45260 16022
rect 45140 15998 45174 16020
rect 45226 15998 45260 16020
rect 45140 15942 45172 15998
rect 45228 15942 45260 15998
rect 45140 15918 45174 15942
rect 45226 15918 45260 15942
rect 45140 15862 45172 15918
rect 45228 15862 45260 15918
rect 45140 15840 45174 15862
rect 45226 15840 45260 15862
rect 45140 15838 45260 15840
rect 45140 15782 45172 15838
rect 45228 15782 45260 15838
rect 45140 15776 45174 15782
rect 45226 15776 45260 15782
rect 45140 15750 45260 15776
rect 45330 5968 45470 6000
rect 45330 5912 45372 5968
rect 45428 5912 45470 5968
rect 45330 5902 45470 5912
rect 45330 5888 45374 5902
rect 45426 5888 45470 5902
rect 45330 5832 45372 5888
rect 45428 5832 45470 5888
rect 45330 5808 45374 5832
rect 45426 5808 45470 5832
rect 45330 5752 45372 5808
rect 45428 5752 45470 5808
rect 45330 5728 45374 5752
rect 45426 5728 45470 5752
rect 45330 5672 45372 5728
rect 45428 5672 45470 5728
rect 45330 5658 45374 5672
rect 45426 5658 45470 5672
rect 45330 5648 45470 5658
rect 45330 5592 45372 5648
rect 45428 5592 45470 5648
rect 45330 5560 45470 5592
<< via2 >>
rect 45372 26406 45428 26408
rect 45372 26354 45374 26406
rect 45374 26354 45426 26406
rect 45426 26354 45428 26406
rect 45372 26352 45428 26354
rect 45372 26290 45374 26328
rect 45374 26290 45426 26328
rect 45426 26290 45428 26328
rect 45372 26278 45428 26290
rect 45372 26272 45374 26278
rect 45374 26272 45426 26278
rect 45426 26272 45428 26278
rect 45372 26226 45374 26248
rect 45374 26226 45426 26248
rect 45426 26226 45428 26248
rect 45372 26214 45428 26226
rect 45372 26192 45374 26214
rect 45374 26192 45426 26214
rect 45426 26192 45428 26214
rect 45372 26162 45374 26168
rect 45374 26162 45426 26168
rect 45426 26162 45428 26168
rect 45372 26150 45428 26162
rect 45372 26112 45374 26150
rect 45374 26112 45426 26150
rect 45426 26112 45428 26150
rect 45372 26086 45428 26088
rect 45372 26034 45374 26086
rect 45374 26034 45426 26086
rect 45426 26034 45428 26086
rect 45372 26032 45428 26034
rect 45172 16672 45174 16718
rect 45174 16672 45226 16718
rect 45226 16672 45228 16718
rect 45172 16662 45228 16672
rect 45172 16608 45174 16638
rect 45174 16608 45226 16638
rect 45226 16608 45228 16638
rect 45172 16596 45228 16608
rect 45172 16582 45174 16596
rect 45174 16582 45226 16596
rect 45226 16582 45228 16596
rect 45172 16544 45174 16558
rect 45174 16544 45226 16558
rect 45226 16544 45228 16558
rect 45172 16532 45228 16544
rect 45172 16502 45174 16532
rect 45174 16502 45226 16532
rect 45226 16502 45228 16532
rect 45172 16468 45228 16478
rect 45172 16422 45174 16468
rect 45174 16422 45226 16468
rect 45226 16422 45228 16468
rect 45172 16352 45174 16398
rect 45174 16352 45226 16398
rect 45226 16352 45228 16398
rect 45172 16342 45228 16352
rect 45172 16288 45174 16318
rect 45174 16288 45226 16318
rect 45226 16288 45228 16318
rect 45172 16276 45228 16288
rect 45172 16262 45174 16276
rect 45174 16262 45226 16276
rect 45226 16262 45228 16276
rect 45172 16224 45174 16238
rect 45174 16224 45226 16238
rect 45226 16224 45228 16238
rect 45172 16212 45228 16224
rect 45172 16182 45174 16212
rect 45174 16182 45226 16212
rect 45226 16182 45228 16212
rect 45172 16148 45228 16158
rect 45172 16102 45174 16148
rect 45174 16102 45226 16148
rect 45226 16102 45228 16148
rect 45172 16032 45174 16078
rect 45174 16032 45226 16078
rect 45226 16032 45228 16078
rect 45172 16022 45228 16032
rect 45172 15968 45174 15998
rect 45174 15968 45226 15998
rect 45226 15968 45228 15998
rect 45172 15956 45228 15968
rect 45172 15942 45174 15956
rect 45174 15942 45226 15956
rect 45226 15942 45228 15956
rect 45172 15904 45174 15918
rect 45174 15904 45226 15918
rect 45226 15904 45228 15918
rect 45172 15892 45228 15904
rect 45172 15862 45174 15892
rect 45174 15862 45226 15892
rect 45226 15862 45228 15892
rect 45172 15828 45228 15838
rect 45172 15782 45174 15828
rect 45174 15782 45226 15828
rect 45226 15782 45228 15828
rect 45372 5966 45428 5968
rect 45372 5914 45374 5966
rect 45374 5914 45426 5966
rect 45426 5914 45428 5966
rect 45372 5912 45428 5914
rect 45372 5850 45374 5888
rect 45374 5850 45426 5888
rect 45426 5850 45428 5888
rect 45372 5838 45428 5850
rect 45372 5832 45374 5838
rect 45374 5832 45426 5838
rect 45426 5832 45428 5838
rect 45372 5786 45374 5808
rect 45374 5786 45426 5808
rect 45426 5786 45428 5808
rect 45372 5774 45428 5786
rect 45372 5752 45374 5774
rect 45374 5752 45426 5774
rect 45426 5752 45428 5774
rect 45372 5722 45374 5728
rect 45374 5722 45426 5728
rect 45426 5722 45428 5728
rect 45372 5710 45428 5722
rect 45372 5672 45374 5710
rect 45374 5672 45426 5710
rect 45426 5672 45428 5710
rect 45372 5646 45428 5648
rect 45372 5594 45374 5646
rect 45374 5594 45426 5646
rect 45426 5594 45428 5646
rect 45372 5592 45428 5594
<< metal3 >>
rect 46000 46752 286000 46800
rect 46000 46448 47008 46752
rect 54992 46448 57008 46752
rect 64992 46448 67008 46752
rect 74992 46448 77008 46752
rect 84992 46448 87008 46752
rect 94992 46448 97008 46752
rect 104992 46448 107008 46752
rect 114992 46448 117008 46752
rect 124992 46448 127008 46752
rect 134992 46448 137008 46752
rect 144992 46448 147008 46752
rect 154992 46448 157008 46752
rect 164992 46448 167008 46752
rect 174992 46448 177008 46752
rect 184992 46448 187008 46752
rect 194992 46448 197008 46752
rect 204992 46448 207008 46752
rect 214992 46448 217008 46752
rect 224992 46448 227008 46752
rect 234992 46448 237008 46752
rect 244992 46448 247008 46752
rect 254992 46448 257008 46752
rect 264992 46448 267008 46752
rect 274992 46448 277008 46752
rect 284992 46448 286000 46752
rect 46000 46000 286000 46448
rect 45330 26412 45470 26440
rect 45330 26348 45368 26412
rect 45432 26348 45470 26412
rect 45330 26332 45470 26348
rect 45330 26268 45368 26332
rect 45432 26268 45470 26332
rect 45330 26252 45470 26268
rect 45330 26188 45368 26252
rect 45432 26188 45470 26252
rect 46000 26200 54400 46000
rect 56000 26200 64400 46000
rect 66000 26200 74400 46000
rect 76000 26200 84400 46000
rect 86000 26200 94400 46000
rect 96000 26200 104400 46000
rect 106000 26200 114400 46000
rect 116000 26200 124400 46000
rect 126000 26200 134400 46000
rect 136000 26200 144400 46000
rect 146000 26200 154400 46000
rect 156000 26200 164400 46000
rect 166000 26200 174400 46000
rect 176000 26200 184400 46000
rect 186000 26200 194400 46000
rect 196000 26200 204400 46000
rect 206000 26200 214400 46000
rect 216000 26200 224400 46000
rect 226000 26200 234400 46000
rect 236000 26200 244400 46000
rect 246000 26200 254400 46000
rect 256000 26200 264400 46000
rect 266000 26200 274400 46000
rect 276000 26200 284400 46000
rect 45330 26172 45470 26188
rect 45330 26108 45368 26172
rect 45432 26108 45470 26172
rect 45330 26092 45470 26108
rect 45330 26028 45368 26092
rect 45432 26028 45470 26092
rect 45330 26000 45470 26028
rect 47600 25800 54400 26200
rect 57600 25800 64400 26200
rect 67600 25800 74400 26200
rect 77600 25800 84400 26200
rect 87600 25800 94400 26200
rect 97600 25800 104400 26200
rect 107600 25800 114400 26200
rect 117600 25800 124400 26200
rect 127600 25800 134400 26200
rect 137600 25800 144400 26200
rect 147600 25800 154400 26200
rect 157600 25800 164400 26200
rect 167600 25800 174400 26200
rect 177600 25800 184400 26200
rect 187600 25800 194400 26200
rect 197600 25800 204400 26200
rect 207600 25800 214400 26200
rect 217600 25800 224400 26200
rect 227600 25800 234400 26200
rect 237600 25800 244400 26200
rect 247600 25800 254400 26200
rect 257600 25800 264400 26200
rect 267600 25800 274400 26200
rect 277600 25800 284400 26200
rect 45140 16722 45260 16750
rect 45140 16658 45168 16722
rect 45232 16658 45260 16722
rect 45140 16642 45260 16658
rect 45140 16578 45168 16642
rect 45232 16578 45260 16642
rect 45140 16562 45260 16578
rect 45140 16498 45168 16562
rect 45232 16498 45260 16562
rect 45140 16482 45260 16498
rect 45140 16418 45168 16482
rect 45232 16418 45260 16482
rect 45140 16402 45260 16418
rect 45140 16338 45168 16402
rect 45232 16338 45260 16402
rect 45140 16322 45260 16338
rect 45140 16258 45168 16322
rect 45232 16258 45260 16322
rect 45140 16242 45260 16258
rect 45140 16178 45168 16242
rect 45232 16178 45260 16242
rect 45140 16162 45260 16178
rect 45140 16098 45168 16162
rect 45232 16098 45260 16162
rect 45140 16082 45260 16098
rect 45140 16018 45168 16082
rect 45232 16018 45260 16082
rect 45140 16002 45260 16018
rect 45140 15938 45168 16002
rect 45232 15938 45260 16002
rect 45140 15922 45260 15938
rect 45140 15858 45168 15922
rect 45232 15858 45260 15922
rect 45140 15842 45260 15858
rect 45140 15778 45168 15842
rect 45232 15778 45260 15842
rect 45140 15750 45260 15778
rect 47600 6000 56000 25800
rect 57600 6000 66000 25800
rect 67600 6000 76000 25800
rect 77600 6000 86000 25800
rect 87600 6000 96000 25800
rect 97600 6000 106000 25800
rect 107600 6000 116000 25800
rect 117600 6000 126000 25800
rect 127600 6000 136000 25800
rect 137600 6000 146000 25800
rect 147600 6000 156000 25800
rect 157600 6000 166000 25800
rect 167600 6000 176000 25800
rect 177600 6000 186000 25800
rect 187600 6000 196000 25800
rect 197600 6000 206000 25800
rect 207600 6000 216000 25800
rect 217600 6000 226000 25800
rect 227600 6000 236000 25800
rect 237600 6000 246000 25800
rect 247600 6000 256000 25800
rect 257600 6000 266000 25800
rect 267600 6000 276000 25800
rect 277600 6000 286000 25800
rect 45330 5972 45470 6000
rect 45330 5908 45368 5972
rect 45432 5908 45470 5972
rect 45330 5892 45470 5908
rect 45330 5828 45368 5892
rect 45432 5828 45470 5892
rect 45330 5812 45470 5828
rect 45330 5748 45368 5812
rect 45432 5748 45470 5812
rect 45330 5732 45470 5748
rect 45330 5668 45368 5732
rect 45432 5668 45470 5732
rect 45330 5652 45470 5668
rect 45330 5588 45368 5652
rect 45432 5588 45470 5652
rect 45330 5560 45470 5588
rect 46000 5552 286000 6000
rect 46000 5248 47008 5552
rect 55952 5248 57008 5552
rect 65952 5248 67008 5552
rect 75952 5248 77008 5552
rect 85952 5248 87008 5552
rect 95952 5248 97008 5552
rect 105952 5248 107008 5552
rect 115952 5248 117008 5552
rect 125952 5248 127008 5552
rect 135952 5248 137008 5552
rect 145952 5248 147008 5552
rect 155952 5248 157008 5552
rect 165952 5248 167008 5552
rect 175952 5248 177008 5552
rect 185952 5248 187008 5552
rect 195952 5248 197008 5552
rect 205952 5248 207008 5552
rect 215952 5248 217008 5552
rect 225952 5248 227008 5552
rect 235952 5248 237008 5552
rect 245952 5248 247008 5552
rect 255952 5248 257008 5552
rect 265952 5248 267008 5552
rect 275952 5248 277008 5552
rect 285952 5248 286000 5552
rect 46000 5200 286000 5248
<< via3 >>
rect 47008 46448 54992 46752
rect 57008 46448 64992 46752
rect 67008 46448 74992 46752
rect 77008 46448 84992 46752
rect 87008 46448 94992 46752
rect 97008 46448 104992 46752
rect 107008 46448 114992 46752
rect 117008 46448 124992 46752
rect 127008 46448 134992 46752
rect 137008 46448 144992 46752
rect 147008 46448 154992 46752
rect 157008 46448 164992 46752
rect 167008 46448 174992 46752
rect 177008 46448 184992 46752
rect 187008 46448 194992 46752
rect 197008 46448 204992 46752
rect 207008 46448 214992 46752
rect 217008 46448 224992 46752
rect 227008 46448 234992 46752
rect 237008 46448 244992 46752
rect 247008 46448 254992 46752
rect 257008 46448 264992 46752
rect 267008 46448 274992 46752
rect 277008 46448 284992 46752
rect 45368 26408 45432 26412
rect 45368 26352 45372 26408
rect 45372 26352 45428 26408
rect 45428 26352 45432 26408
rect 45368 26348 45432 26352
rect 45368 26328 45432 26332
rect 45368 26272 45372 26328
rect 45372 26272 45428 26328
rect 45428 26272 45432 26328
rect 45368 26268 45432 26272
rect 45368 26248 45432 26252
rect 45368 26192 45372 26248
rect 45372 26192 45428 26248
rect 45428 26192 45432 26248
rect 45368 26188 45432 26192
rect 45368 26168 45432 26172
rect 45368 26112 45372 26168
rect 45372 26112 45428 26168
rect 45428 26112 45432 26168
rect 45368 26108 45432 26112
rect 45368 26088 45432 26092
rect 45368 26032 45372 26088
rect 45372 26032 45428 26088
rect 45428 26032 45432 26088
rect 45368 26028 45432 26032
rect 45168 16718 45232 16722
rect 45168 16662 45172 16718
rect 45172 16662 45228 16718
rect 45228 16662 45232 16718
rect 45168 16658 45232 16662
rect 45168 16638 45232 16642
rect 45168 16582 45172 16638
rect 45172 16582 45228 16638
rect 45228 16582 45232 16638
rect 45168 16578 45232 16582
rect 45168 16558 45232 16562
rect 45168 16502 45172 16558
rect 45172 16502 45228 16558
rect 45228 16502 45232 16558
rect 45168 16498 45232 16502
rect 45168 16478 45232 16482
rect 45168 16422 45172 16478
rect 45172 16422 45228 16478
rect 45228 16422 45232 16478
rect 45168 16418 45232 16422
rect 45168 16398 45232 16402
rect 45168 16342 45172 16398
rect 45172 16342 45228 16398
rect 45228 16342 45232 16398
rect 45168 16338 45232 16342
rect 45168 16318 45232 16322
rect 45168 16262 45172 16318
rect 45172 16262 45228 16318
rect 45228 16262 45232 16318
rect 45168 16258 45232 16262
rect 45168 16238 45232 16242
rect 45168 16182 45172 16238
rect 45172 16182 45228 16238
rect 45228 16182 45232 16238
rect 45168 16178 45232 16182
rect 45168 16158 45232 16162
rect 45168 16102 45172 16158
rect 45172 16102 45228 16158
rect 45228 16102 45232 16158
rect 45168 16098 45232 16102
rect 45168 16078 45232 16082
rect 45168 16022 45172 16078
rect 45172 16022 45228 16078
rect 45228 16022 45232 16078
rect 45168 16018 45232 16022
rect 45168 15998 45232 16002
rect 45168 15942 45172 15998
rect 45172 15942 45228 15998
rect 45228 15942 45232 15998
rect 45168 15938 45232 15942
rect 45168 15918 45232 15922
rect 45168 15862 45172 15918
rect 45172 15862 45228 15918
rect 45228 15862 45232 15918
rect 45168 15858 45232 15862
rect 45168 15838 45232 15842
rect 45168 15782 45172 15838
rect 45172 15782 45228 15838
rect 45228 15782 45232 15838
rect 45168 15778 45232 15782
rect 45368 5968 45432 5972
rect 45368 5912 45372 5968
rect 45372 5912 45428 5968
rect 45428 5912 45432 5968
rect 45368 5908 45432 5912
rect 45368 5888 45432 5892
rect 45368 5832 45372 5888
rect 45372 5832 45428 5888
rect 45428 5832 45432 5888
rect 45368 5828 45432 5832
rect 45368 5808 45432 5812
rect 45368 5752 45372 5808
rect 45372 5752 45428 5808
rect 45428 5752 45432 5808
rect 45368 5748 45432 5752
rect 45368 5728 45432 5732
rect 45368 5672 45372 5728
rect 45372 5672 45428 5728
rect 45428 5672 45432 5728
rect 45368 5668 45432 5672
rect 45368 5648 45432 5652
rect 45368 5592 45372 5648
rect 45372 5592 45428 5648
rect 45428 5592 45432 5648
rect 45368 5588 45432 5592
rect 47008 5248 55952 5552
rect 57008 5248 65952 5552
rect 67008 5248 75952 5552
rect 77008 5248 85952 5552
rect 87008 5248 95952 5552
rect 97008 5248 105952 5552
rect 107008 5248 115952 5552
rect 117008 5248 125952 5552
rect 127008 5248 135952 5552
rect 137008 5248 145952 5552
rect 147008 5248 155952 5552
rect 157008 5248 165952 5552
rect 167008 5248 175952 5552
rect 177008 5248 185952 5552
rect 187008 5248 195952 5552
rect 197008 5248 205952 5552
rect 207008 5248 215952 5552
rect 217008 5248 225952 5552
rect 227008 5248 235952 5552
rect 237008 5248 245952 5552
rect 247008 5248 255952 5552
rect 257008 5248 265952 5552
rect 267008 5248 275952 5552
rect 277008 5248 285952 5552
<< mimcap >>
rect 46040 45932 54360 45960
rect 46040 26268 46088 45932
rect 54312 26268 54360 45932
rect 46040 26240 54360 26268
rect 56040 45932 64360 45960
rect 56040 26268 56088 45932
rect 64312 26268 64360 45932
rect 56040 26240 64360 26268
rect 66040 45932 74360 45960
rect 66040 26268 66088 45932
rect 74312 26268 74360 45932
rect 66040 26240 74360 26268
rect 76040 45932 84360 45960
rect 76040 26268 76088 45932
rect 84312 26268 84360 45932
rect 76040 26240 84360 26268
rect 86040 45932 94360 45960
rect 86040 26268 86088 45932
rect 94312 26268 94360 45932
rect 86040 26240 94360 26268
rect 96040 45932 104360 45960
rect 96040 26268 96088 45932
rect 104312 26268 104360 45932
rect 96040 26240 104360 26268
rect 106040 45932 114360 45960
rect 106040 26268 106088 45932
rect 114312 26268 114360 45932
rect 106040 26240 114360 26268
rect 116040 45932 124360 45960
rect 116040 26268 116088 45932
rect 124312 26268 124360 45932
rect 116040 26240 124360 26268
rect 126040 45932 134360 45960
rect 126040 26268 126088 45932
rect 134312 26268 134360 45932
rect 126040 26240 134360 26268
rect 136040 45932 144360 45960
rect 136040 26268 136088 45932
rect 144312 26268 144360 45932
rect 136040 26240 144360 26268
rect 146040 45932 154360 45960
rect 146040 26268 146088 45932
rect 154312 26268 154360 45932
rect 146040 26240 154360 26268
rect 156040 45932 164360 45960
rect 156040 26268 156088 45932
rect 164312 26268 164360 45932
rect 156040 26240 164360 26268
rect 166040 45932 174360 45960
rect 166040 26268 166088 45932
rect 174312 26268 174360 45932
rect 166040 26240 174360 26268
rect 176040 45932 184360 45960
rect 176040 26268 176088 45932
rect 184312 26268 184360 45932
rect 176040 26240 184360 26268
rect 186040 45932 194360 45960
rect 186040 26268 186088 45932
rect 194312 26268 194360 45932
rect 186040 26240 194360 26268
rect 196040 45932 204360 45960
rect 196040 26268 196088 45932
rect 204312 26268 204360 45932
rect 196040 26240 204360 26268
rect 206040 45932 214360 45960
rect 206040 26268 206088 45932
rect 214312 26268 214360 45932
rect 206040 26240 214360 26268
rect 216040 45932 224360 45960
rect 216040 26268 216088 45932
rect 224312 26268 224360 45932
rect 216040 26240 224360 26268
rect 226040 45932 234360 45960
rect 226040 26268 226088 45932
rect 234312 26268 234360 45932
rect 226040 26240 234360 26268
rect 236040 45932 244360 45960
rect 236040 26268 236088 45932
rect 244312 26268 244360 45932
rect 236040 26240 244360 26268
rect 246040 45932 254360 45960
rect 246040 26268 246088 45932
rect 254312 26268 254360 45932
rect 246040 26240 254360 26268
rect 256040 45932 264360 45960
rect 256040 26268 256088 45932
rect 264312 26268 264360 45932
rect 256040 26240 264360 26268
rect 266040 45932 274360 45960
rect 266040 26268 266088 45932
rect 274312 26268 274360 45932
rect 266040 26240 274360 26268
rect 276040 45932 284360 45960
rect 276040 26268 276088 45932
rect 284312 26268 284360 45932
rect 276040 26240 284360 26268
rect 47640 25732 55960 25760
rect 47640 6068 47688 25732
rect 55912 6068 55960 25732
rect 47640 6040 55960 6068
rect 57640 25732 65960 25760
rect 57640 6068 57688 25732
rect 65912 6068 65960 25732
rect 57640 6040 65960 6068
rect 67640 25732 75960 25760
rect 67640 6068 67688 25732
rect 75912 6068 75960 25732
rect 67640 6040 75960 6068
rect 77640 25732 85960 25760
rect 77640 6068 77688 25732
rect 85912 6068 85960 25732
rect 77640 6040 85960 6068
rect 87640 25732 95960 25760
rect 87640 6068 87688 25732
rect 95912 6068 95960 25732
rect 87640 6040 95960 6068
rect 97640 25732 105960 25760
rect 97640 6068 97688 25732
rect 105912 6068 105960 25732
rect 97640 6040 105960 6068
rect 107640 25732 115960 25760
rect 107640 6068 107688 25732
rect 115912 6068 115960 25732
rect 107640 6040 115960 6068
rect 117640 25732 125960 25760
rect 117640 6068 117688 25732
rect 125912 6068 125960 25732
rect 117640 6040 125960 6068
rect 127640 25732 135960 25760
rect 127640 6068 127688 25732
rect 135912 6068 135960 25732
rect 127640 6040 135960 6068
rect 137640 25732 145960 25760
rect 137640 6068 137688 25732
rect 145912 6068 145960 25732
rect 137640 6040 145960 6068
rect 147640 25732 155960 25760
rect 147640 6068 147688 25732
rect 155912 6068 155960 25732
rect 147640 6040 155960 6068
rect 157640 25732 165960 25760
rect 157640 6068 157688 25732
rect 165912 6068 165960 25732
rect 157640 6040 165960 6068
rect 167640 25732 175960 25760
rect 167640 6068 167688 25732
rect 175912 6068 175960 25732
rect 167640 6040 175960 6068
rect 177640 25732 185960 25760
rect 177640 6068 177688 25732
rect 185912 6068 185960 25732
rect 177640 6040 185960 6068
rect 187640 25732 195960 25760
rect 187640 6068 187688 25732
rect 195912 6068 195960 25732
rect 187640 6040 195960 6068
rect 197640 25732 205960 25760
rect 197640 6068 197688 25732
rect 205912 6068 205960 25732
rect 197640 6040 205960 6068
rect 207640 25732 215960 25760
rect 207640 6068 207688 25732
rect 215912 6068 215960 25732
rect 207640 6040 215960 6068
rect 217640 25732 225960 25760
rect 217640 6068 217688 25732
rect 225912 6068 225960 25732
rect 217640 6040 225960 6068
rect 227640 25732 235960 25760
rect 227640 6068 227688 25732
rect 235912 6068 235960 25732
rect 227640 6040 235960 6068
rect 237640 25732 245960 25760
rect 237640 6068 237688 25732
rect 245912 6068 245960 25732
rect 237640 6040 245960 6068
rect 247640 25732 255960 25760
rect 247640 6068 247688 25732
rect 255912 6068 255960 25732
rect 247640 6040 255960 6068
rect 257640 25732 265960 25760
rect 257640 6068 257688 25732
rect 265912 6068 265960 25732
rect 257640 6040 265960 6068
rect 267640 25732 275960 25760
rect 267640 6068 267688 25732
rect 275912 6068 275960 25732
rect 267640 6040 275960 6068
rect 277640 25732 285960 25760
rect 277640 6068 277688 25732
rect 285912 6068 285960 25732
rect 277640 6040 285960 6068
<< mimcapcontact >>
rect 46088 26268 54312 45932
rect 56088 26268 64312 45932
rect 66088 26268 74312 45932
rect 76088 26268 84312 45932
rect 86088 26268 94312 45932
rect 96088 26268 104312 45932
rect 106088 26268 114312 45932
rect 116088 26268 124312 45932
rect 126088 26268 134312 45932
rect 136088 26268 144312 45932
rect 146088 26268 154312 45932
rect 156088 26268 164312 45932
rect 166088 26268 174312 45932
rect 176088 26268 184312 45932
rect 186088 26268 194312 45932
rect 196088 26268 204312 45932
rect 206088 26268 214312 45932
rect 216088 26268 224312 45932
rect 226088 26268 234312 45932
rect 236088 26268 244312 45932
rect 246088 26268 254312 45932
rect 256088 26268 264312 45932
rect 266088 26268 274312 45932
rect 276088 26268 284312 45932
rect 47688 6068 55912 25732
rect 57688 6068 65912 25732
rect 67688 6068 75912 25732
rect 77688 6068 85912 25732
rect 87688 6068 95912 25732
rect 97688 6068 105912 25732
rect 107688 6068 115912 25732
rect 117688 6068 125912 25732
rect 127688 6068 135912 25732
rect 137688 6068 145912 25732
rect 147688 6068 155912 25732
rect 157688 6068 165912 25732
rect 167688 6068 175912 25732
rect 177688 6068 185912 25732
rect 187688 6068 195912 25732
rect 197688 6068 205912 25732
rect 207688 6068 215912 25732
rect 217688 6068 225912 25732
rect 227688 6068 235912 25732
rect 237688 6068 245912 25732
rect 247688 6068 255912 25732
rect 257688 6068 265912 25732
rect 267688 6068 275912 25732
rect 277688 6068 285912 25732
<< metal4 >>
rect 46000 46752 286000 46800
rect 46000 46448 47008 46752
rect 54992 46448 57008 46752
rect 64992 46448 67008 46752
rect 74992 46448 77008 46752
rect 84992 46448 87008 46752
rect 94992 46448 97008 46752
rect 104992 46448 107008 46752
rect 114992 46448 117008 46752
rect 124992 46448 127008 46752
rect 134992 46448 137008 46752
rect 144992 46448 147008 46752
rect 154992 46448 157008 46752
rect 164992 46448 167008 46752
rect 174992 46448 177008 46752
rect 184992 46448 187008 46752
rect 194992 46448 197008 46752
rect 204992 46448 207008 46752
rect 214992 46448 217008 46752
rect 224992 46448 227008 46752
rect 234992 46448 237008 46752
rect 244992 46448 247008 46752
rect 254992 46448 257008 46752
rect 264992 46448 267008 46752
rect 274992 46448 277008 46752
rect 284992 46448 286000 46752
rect 46000 46400 286000 46448
rect 46000 45932 284400 46000
rect 43800 26412 45600 26600
rect 43800 26378 45368 26412
rect 43800 25822 44062 26378
rect 44938 26348 45368 26378
rect 45432 26400 45600 26412
rect 46000 26400 46088 45932
rect 45432 26348 46088 26400
rect 44938 26332 46088 26348
rect 44938 26268 45368 26332
rect 45432 26268 46088 26332
rect 54312 45600 56088 45932
rect 54312 26400 54400 45600
rect 56000 26400 56088 45600
rect 54312 26268 56088 26400
rect 64312 45600 66088 45932
rect 64312 26400 64400 45600
rect 66000 26400 66088 45600
rect 64312 26268 66088 26400
rect 74312 45600 76088 45932
rect 74312 26400 74400 45600
rect 76000 26400 76088 45600
rect 74312 26268 76088 26400
rect 84312 45600 86088 45932
rect 84312 26400 84400 45600
rect 86000 26400 86088 45600
rect 84312 26268 86088 26400
rect 94312 45600 96088 45932
rect 94312 26400 94400 45600
rect 96000 26400 96088 45600
rect 94312 26268 96088 26400
rect 104312 45600 106088 45932
rect 104312 26400 104400 45600
rect 106000 26400 106088 45600
rect 104312 26268 106088 26400
rect 114312 45600 116088 45932
rect 114312 26400 114400 45600
rect 116000 26400 116088 45600
rect 114312 26268 116088 26400
rect 124312 45600 126088 45932
rect 124312 26400 124400 45600
rect 126000 26400 126088 45600
rect 124312 26268 126088 26400
rect 134312 45600 136088 45932
rect 134312 26400 134400 45600
rect 136000 26400 136088 45600
rect 134312 26268 136088 26400
rect 144312 45600 146088 45932
rect 144312 26400 144400 45600
rect 146000 26400 146088 45600
rect 144312 26268 146088 26400
rect 154312 45600 156088 45932
rect 154312 26400 154400 45600
rect 156000 26400 156088 45600
rect 154312 26268 156088 26400
rect 164312 45600 166088 45932
rect 164312 26400 164400 45600
rect 166000 26400 166088 45600
rect 164312 26268 166088 26400
rect 174312 45600 176088 45932
rect 174312 26400 174400 45600
rect 176000 26400 176088 45600
rect 174312 26268 176088 26400
rect 184312 45600 186088 45932
rect 184312 26400 184400 45600
rect 186000 26400 186088 45600
rect 184312 26268 186088 26400
rect 194312 45600 196088 45932
rect 194312 26400 194400 45600
rect 196000 26400 196088 45600
rect 194312 26268 196088 26400
rect 204312 45600 206088 45932
rect 204312 26400 204400 45600
rect 206000 26400 206088 45600
rect 204312 26268 206088 26400
rect 214312 45600 216088 45932
rect 214312 26400 214400 45600
rect 216000 26400 216088 45600
rect 214312 26268 216088 26400
rect 224312 45600 226088 45932
rect 224312 26400 224400 45600
rect 226000 26400 226088 45600
rect 224312 26268 226088 26400
rect 234312 45600 236088 45932
rect 234312 26400 234400 45600
rect 236000 26400 236088 45600
rect 234312 26268 236088 26400
rect 244312 45600 246088 45932
rect 244312 26400 244400 45600
rect 246000 26400 246088 45600
rect 244312 26268 246088 26400
rect 254312 45600 256088 45932
rect 254312 26400 254400 45600
rect 256000 26400 256088 45600
rect 254312 26268 256088 26400
rect 264312 45600 266088 45932
rect 264312 26400 264400 45600
rect 266000 26400 266088 45600
rect 264312 26268 266088 26400
rect 274312 45600 276088 45932
rect 274312 26400 274400 45600
rect 276000 26400 276088 45600
rect 274312 26268 276088 26400
rect 284312 26268 284400 45932
rect 44938 26252 284400 26268
rect 44938 26188 45368 26252
rect 45432 26188 284400 26252
rect 44938 26172 284400 26188
rect 44938 26108 45368 26172
rect 45432 26108 284400 26172
rect 44938 26092 284400 26108
rect 44938 26028 45368 26092
rect 45432 26028 284400 26092
rect 44938 25822 284400 26028
rect 43800 25800 284400 25822
rect 43800 25732 286000 25800
rect 43800 25600 47688 25732
rect 45040 16722 45260 16750
rect 45040 16658 45168 16722
rect 45232 16658 45260 16722
rect 45040 16642 45260 16658
rect 45040 16578 45168 16642
rect 45232 16578 45260 16642
rect 45040 16562 45260 16578
rect 45040 16498 45168 16562
rect 45232 16498 45260 16562
rect 45040 16482 45260 16498
rect 45040 16418 45168 16482
rect 45232 16418 45260 16482
rect 45040 16402 45260 16418
rect 45040 16338 45168 16402
rect 45232 16338 45260 16402
rect 45040 16322 45260 16338
rect 45040 16258 45168 16322
rect 45232 16258 45260 16322
rect 45040 16242 45260 16258
rect 45040 16178 45168 16242
rect 45232 16178 45260 16242
rect 45040 16162 45260 16178
rect 45040 16098 45168 16162
rect 45232 16098 45260 16162
rect 45040 16082 45260 16098
rect 45040 16018 45168 16082
rect 45232 16018 45260 16082
rect 45040 16002 45260 16018
rect 45040 15938 45168 16002
rect 45232 15938 45260 16002
rect 45040 15922 45260 15938
rect 45040 15858 45168 15922
rect 45232 15858 45260 15922
rect 45040 15842 45260 15858
rect 45040 15778 45168 15842
rect 45232 15778 45260 15842
rect 45040 15750 45260 15778
rect 43800 6178 45600 6400
rect 43800 5622 44062 6178
rect 44938 5972 45600 6178
rect 47600 6068 47688 25600
rect 55912 25600 57688 25732
rect 55912 6400 56000 25600
rect 57600 6400 57688 25600
rect 55912 6068 57688 6400
rect 65912 25600 67688 25732
rect 65912 6400 66000 25600
rect 67600 6400 67688 25600
rect 65912 6068 67688 6400
rect 75912 25600 77688 25732
rect 75912 6400 76000 25600
rect 77600 6400 77688 25600
rect 75912 6068 77688 6400
rect 85912 25600 87688 25732
rect 85912 6400 86000 25600
rect 87600 6400 87688 25600
rect 85912 6068 87688 6400
rect 95912 25600 97688 25732
rect 95912 6400 96000 25600
rect 97600 6400 97688 25600
rect 95912 6068 97688 6400
rect 105912 25600 107688 25732
rect 105912 6400 106000 25600
rect 107600 6400 107688 25600
rect 105912 6068 107688 6400
rect 115912 25600 117688 25732
rect 115912 6400 116000 25600
rect 117600 6400 117688 25600
rect 115912 6068 117688 6400
rect 125912 25600 127688 25732
rect 125912 6400 126000 25600
rect 127600 6400 127688 25600
rect 125912 6068 127688 6400
rect 135912 25600 137688 25732
rect 135912 6400 136000 25600
rect 137600 6400 137688 25600
rect 135912 6068 137688 6400
rect 145912 25600 147688 25732
rect 145912 6400 146000 25600
rect 147600 6400 147688 25600
rect 145912 6068 147688 6400
rect 155912 25600 157688 25732
rect 155912 6400 156000 25600
rect 157600 6400 157688 25600
rect 155912 6068 157688 6400
rect 165912 25600 167688 25732
rect 165912 6400 166000 25600
rect 167600 6400 167688 25600
rect 165912 6068 167688 6400
rect 175912 25600 177688 25732
rect 175912 6400 176000 25600
rect 177600 6400 177688 25600
rect 175912 6068 177688 6400
rect 185912 25600 187688 25732
rect 185912 6400 186000 25600
rect 187600 6400 187688 25600
rect 185912 6068 187688 6400
rect 195912 25600 197688 25732
rect 195912 6400 196000 25600
rect 197600 6400 197688 25600
rect 195912 6068 197688 6400
rect 205912 25600 207688 25732
rect 205912 6400 206000 25600
rect 207600 6400 207688 25600
rect 205912 6068 207688 6400
rect 215912 25600 217688 25732
rect 215912 6400 216000 25600
rect 217600 6400 217688 25600
rect 215912 6068 217688 6400
rect 225912 25600 227688 25732
rect 225912 6400 226000 25600
rect 227600 6400 227688 25600
rect 225912 6068 227688 6400
rect 235912 25600 237688 25732
rect 235912 6400 236000 25600
rect 237600 6400 237688 25600
rect 235912 6068 237688 6400
rect 245912 25600 247688 25732
rect 245912 6400 246000 25600
rect 247600 6400 247688 25600
rect 245912 6068 247688 6400
rect 255912 25600 257688 25732
rect 255912 6400 256000 25600
rect 257600 6400 257688 25600
rect 255912 6068 257688 6400
rect 265912 25600 267688 25732
rect 265912 6400 266000 25600
rect 267600 6400 267688 25600
rect 265912 6068 267688 6400
rect 275912 25600 277688 25732
rect 275912 6400 276000 25600
rect 277600 6400 277688 25600
rect 275912 6068 277688 6400
rect 285912 6068 286000 25732
rect 47600 6000 286000 6068
rect 44938 5908 45368 5972
rect 45432 5908 45600 5972
rect 44938 5892 45600 5908
rect 44938 5828 45368 5892
rect 45432 5828 45600 5892
rect 44938 5812 45600 5828
rect 44938 5748 45368 5812
rect 45432 5800 45600 5812
rect 45432 5748 46000 5800
rect 44938 5732 46000 5748
rect 44938 5668 45368 5732
rect 45432 5668 46000 5732
rect 44938 5652 46000 5668
rect 44938 5622 45368 5652
rect 43800 5588 45368 5622
rect 45432 5600 46000 5652
rect 45432 5588 286000 5600
rect 43800 5552 286000 5588
rect 43800 5400 47008 5552
rect 46000 5248 47008 5400
rect 55952 5248 57008 5552
rect 65952 5248 67008 5552
rect 75952 5248 77008 5552
rect 85952 5248 87008 5552
rect 95952 5248 97008 5552
rect 105952 5248 107008 5552
rect 115952 5248 117008 5552
rect 125952 5248 127008 5552
rect 135952 5248 137008 5552
rect 145952 5248 147008 5552
rect 155952 5248 157008 5552
rect 165952 5248 167008 5552
rect 175952 5248 177008 5552
rect 185952 5248 187008 5552
rect 195952 5248 197008 5552
rect 205952 5248 207008 5552
rect 215952 5248 217008 5552
rect 225952 5248 227008 5552
rect 235952 5248 237008 5552
rect 245952 5248 247008 5552
rect 255952 5248 257008 5552
rect 265952 5248 267008 5552
rect 275952 5248 277008 5552
rect 285952 5248 286000 5552
rect 46000 5200 286000 5248
<< via4 >>
rect 47042 46482 47278 46718
rect 47362 46482 47598 46718
rect 47682 46482 47918 46718
rect 48002 46482 48238 46718
rect 48322 46482 48558 46718
rect 48642 46482 48878 46718
rect 48962 46482 49198 46718
rect 49282 46482 49518 46718
rect 49602 46482 49838 46718
rect 49922 46482 50158 46718
rect 50242 46482 50478 46718
rect 50562 46482 50798 46718
rect 50882 46482 51118 46718
rect 51202 46482 51438 46718
rect 51522 46482 51758 46718
rect 51842 46482 52078 46718
rect 52162 46482 52398 46718
rect 52482 46482 52718 46718
rect 52802 46482 53038 46718
rect 53122 46482 53358 46718
rect 53442 46482 53678 46718
rect 53762 46482 53998 46718
rect 54082 46482 54318 46718
rect 54402 46482 54638 46718
rect 54722 46482 54958 46718
rect 57042 46482 57278 46718
rect 57362 46482 57598 46718
rect 57682 46482 57918 46718
rect 58002 46482 58238 46718
rect 58322 46482 58558 46718
rect 58642 46482 58878 46718
rect 58962 46482 59198 46718
rect 59282 46482 59518 46718
rect 59602 46482 59838 46718
rect 59922 46482 60158 46718
rect 60242 46482 60478 46718
rect 60562 46482 60798 46718
rect 60882 46482 61118 46718
rect 61202 46482 61438 46718
rect 61522 46482 61758 46718
rect 61842 46482 62078 46718
rect 62162 46482 62398 46718
rect 62482 46482 62718 46718
rect 62802 46482 63038 46718
rect 63122 46482 63358 46718
rect 63442 46482 63678 46718
rect 63762 46482 63998 46718
rect 64082 46482 64318 46718
rect 64402 46482 64638 46718
rect 64722 46482 64958 46718
rect 67042 46482 67278 46718
rect 67362 46482 67598 46718
rect 67682 46482 67918 46718
rect 68002 46482 68238 46718
rect 68322 46482 68558 46718
rect 68642 46482 68878 46718
rect 68962 46482 69198 46718
rect 69282 46482 69518 46718
rect 69602 46482 69838 46718
rect 69922 46482 70158 46718
rect 70242 46482 70478 46718
rect 70562 46482 70798 46718
rect 70882 46482 71118 46718
rect 71202 46482 71438 46718
rect 71522 46482 71758 46718
rect 71842 46482 72078 46718
rect 72162 46482 72398 46718
rect 72482 46482 72718 46718
rect 72802 46482 73038 46718
rect 73122 46482 73358 46718
rect 73442 46482 73678 46718
rect 73762 46482 73998 46718
rect 74082 46482 74318 46718
rect 74402 46482 74638 46718
rect 74722 46482 74958 46718
rect 77042 46482 77278 46718
rect 77362 46482 77598 46718
rect 77682 46482 77918 46718
rect 78002 46482 78238 46718
rect 78322 46482 78558 46718
rect 78642 46482 78878 46718
rect 78962 46482 79198 46718
rect 79282 46482 79518 46718
rect 79602 46482 79838 46718
rect 79922 46482 80158 46718
rect 80242 46482 80478 46718
rect 80562 46482 80798 46718
rect 80882 46482 81118 46718
rect 81202 46482 81438 46718
rect 81522 46482 81758 46718
rect 81842 46482 82078 46718
rect 82162 46482 82398 46718
rect 82482 46482 82718 46718
rect 82802 46482 83038 46718
rect 83122 46482 83358 46718
rect 83442 46482 83678 46718
rect 83762 46482 83998 46718
rect 84082 46482 84318 46718
rect 84402 46482 84638 46718
rect 84722 46482 84958 46718
rect 87042 46482 87278 46718
rect 87362 46482 87598 46718
rect 87682 46482 87918 46718
rect 88002 46482 88238 46718
rect 88322 46482 88558 46718
rect 88642 46482 88878 46718
rect 88962 46482 89198 46718
rect 89282 46482 89518 46718
rect 89602 46482 89838 46718
rect 89922 46482 90158 46718
rect 90242 46482 90478 46718
rect 90562 46482 90798 46718
rect 90882 46482 91118 46718
rect 91202 46482 91438 46718
rect 91522 46482 91758 46718
rect 91842 46482 92078 46718
rect 92162 46482 92398 46718
rect 92482 46482 92718 46718
rect 92802 46482 93038 46718
rect 93122 46482 93358 46718
rect 93442 46482 93678 46718
rect 93762 46482 93998 46718
rect 94082 46482 94318 46718
rect 94402 46482 94638 46718
rect 94722 46482 94958 46718
rect 97042 46482 97278 46718
rect 97362 46482 97598 46718
rect 97682 46482 97918 46718
rect 98002 46482 98238 46718
rect 98322 46482 98558 46718
rect 98642 46482 98878 46718
rect 98962 46482 99198 46718
rect 99282 46482 99518 46718
rect 99602 46482 99838 46718
rect 99922 46482 100158 46718
rect 100242 46482 100478 46718
rect 100562 46482 100798 46718
rect 100882 46482 101118 46718
rect 101202 46482 101438 46718
rect 101522 46482 101758 46718
rect 101842 46482 102078 46718
rect 102162 46482 102398 46718
rect 102482 46482 102718 46718
rect 102802 46482 103038 46718
rect 103122 46482 103358 46718
rect 103442 46482 103678 46718
rect 103762 46482 103998 46718
rect 104082 46482 104318 46718
rect 104402 46482 104638 46718
rect 104722 46482 104958 46718
rect 107042 46482 107278 46718
rect 107362 46482 107598 46718
rect 107682 46482 107918 46718
rect 108002 46482 108238 46718
rect 108322 46482 108558 46718
rect 108642 46482 108878 46718
rect 108962 46482 109198 46718
rect 109282 46482 109518 46718
rect 109602 46482 109838 46718
rect 109922 46482 110158 46718
rect 110242 46482 110478 46718
rect 110562 46482 110798 46718
rect 110882 46482 111118 46718
rect 111202 46482 111438 46718
rect 111522 46482 111758 46718
rect 111842 46482 112078 46718
rect 112162 46482 112398 46718
rect 112482 46482 112718 46718
rect 112802 46482 113038 46718
rect 113122 46482 113358 46718
rect 113442 46482 113678 46718
rect 113762 46482 113998 46718
rect 114082 46482 114318 46718
rect 114402 46482 114638 46718
rect 114722 46482 114958 46718
rect 117042 46482 117278 46718
rect 117362 46482 117598 46718
rect 117682 46482 117918 46718
rect 118002 46482 118238 46718
rect 118322 46482 118558 46718
rect 118642 46482 118878 46718
rect 118962 46482 119198 46718
rect 119282 46482 119518 46718
rect 119602 46482 119838 46718
rect 119922 46482 120158 46718
rect 120242 46482 120478 46718
rect 120562 46482 120798 46718
rect 120882 46482 121118 46718
rect 121202 46482 121438 46718
rect 121522 46482 121758 46718
rect 121842 46482 122078 46718
rect 122162 46482 122398 46718
rect 122482 46482 122718 46718
rect 122802 46482 123038 46718
rect 123122 46482 123358 46718
rect 123442 46482 123678 46718
rect 123762 46482 123998 46718
rect 124082 46482 124318 46718
rect 124402 46482 124638 46718
rect 124722 46482 124958 46718
rect 127042 46482 127278 46718
rect 127362 46482 127598 46718
rect 127682 46482 127918 46718
rect 128002 46482 128238 46718
rect 128322 46482 128558 46718
rect 128642 46482 128878 46718
rect 128962 46482 129198 46718
rect 129282 46482 129518 46718
rect 129602 46482 129838 46718
rect 129922 46482 130158 46718
rect 130242 46482 130478 46718
rect 130562 46482 130798 46718
rect 130882 46482 131118 46718
rect 131202 46482 131438 46718
rect 131522 46482 131758 46718
rect 131842 46482 132078 46718
rect 132162 46482 132398 46718
rect 132482 46482 132718 46718
rect 132802 46482 133038 46718
rect 133122 46482 133358 46718
rect 133442 46482 133678 46718
rect 133762 46482 133998 46718
rect 134082 46482 134318 46718
rect 134402 46482 134638 46718
rect 134722 46482 134958 46718
rect 137042 46482 137278 46718
rect 137362 46482 137598 46718
rect 137682 46482 137918 46718
rect 138002 46482 138238 46718
rect 138322 46482 138558 46718
rect 138642 46482 138878 46718
rect 138962 46482 139198 46718
rect 139282 46482 139518 46718
rect 139602 46482 139838 46718
rect 139922 46482 140158 46718
rect 140242 46482 140478 46718
rect 140562 46482 140798 46718
rect 140882 46482 141118 46718
rect 141202 46482 141438 46718
rect 141522 46482 141758 46718
rect 141842 46482 142078 46718
rect 142162 46482 142398 46718
rect 142482 46482 142718 46718
rect 142802 46482 143038 46718
rect 143122 46482 143358 46718
rect 143442 46482 143678 46718
rect 143762 46482 143998 46718
rect 144082 46482 144318 46718
rect 144402 46482 144638 46718
rect 144722 46482 144958 46718
rect 147042 46482 147278 46718
rect 147362 46482 147598 46718
rect 147682 46482 147918 46718
rect 148002 46482 148238 46718
rect 148322 46482 148558 46718
rect 148642 46482 148878 46718
rect 148962 46482 149198 46718
rect 149282 46482 149518 46718
rect 149602 46482 149838 46718
rect 149922 46482 150158 46718
rect 150242 46482 150478 46718
rect 150562 46482 150798 46718
rect 150882 46482 151118 46718
rect 151202 46482 151438 46718
rect 151522 46482 151758 46718
rect 151842 46482 152078 46718
rect 152162 46482 152398 46718
rect 152482 46482 152718 46718
rect 152802 46482 153038 46718
rect 153122 46482 153358 46718
rect 153442 46482 153678 46718
rect 153762 46482 153998 46718
rect 154082 46482 154318 46718
rect 154402 46482 154638 46718
rect 154722 46482 154958 46718
rect 157042 46482 157278 46718
rect 157362 46482 157598 46718
rect 157682 46482 157918 46718
rect 158002 46482 158238 46718
rect 158322 46482 158558 46718
rect 158642 46482 158878 46718
rect 158962 46482 159198 46718
rect 159282 46482 159518 46718
rect 159602 46482 159838 46718
rect 159922 46482 160158 46718
rect 160242 46482 160478 46718
rect 160562 46482 160798 46718
rect 160882 46482 161118 46718
rect 161202 46482 161438 46718
rect 161522 46482 161758 46718
rect 161842 46482 162078 46718
rect 162162 46482 162398 46718
rect 162482 46482 162718 46718
rect 162802 46482 163038 46718
rect 163122 46482 163358 46718
rect 163442 46482 163678 46718
rect 163762 46482 163998 46718
rect 164082 46482 164318 46718
rect 164402 46482 164638 46718
rect 164722 46482 164958 46718
rect 167042 46482 167278 46718
rect 167362 46482 167598 46718
rect 167682 46482 167918 46718
rect 168002 46482 168238 46718
rect 168322 46482 168558 46718
rect 168642 46482 168878 46718
rect 168962 46482 169198 46718
rect 169282 46482 169518 46718
rect 169602 46482 169838 46718
rect 169922 46482 170158 46718
rect 170242 46482 170478 46718
rect 170562 46482 170798 46718
rect 170882 46482 171118 46718
rect 171202 46482 171438 46718
rect 171522 46482 171758 46718
rect 171842 46482 172078 46718
rect 172162 46482 172398 46718
rect 172482 46482 172718 46718
rect 172802 46482 173038 46718
rect 173122 46482 173358 46718
rect 173442 46482 173678 46718
rect 173762 46482 173998 46718
rect 174082 46482 174318 46718
rect 174402 46482 174638 46718
rect 174722 46482 174958 46718
rect 177042 46482 177278 46718
rect 177362 46482 177598 46718
rect 177682 46482 177918 46718
rect 178002 46482 178238 46718
rect 178322 46482 178558 46718
rect 178642 46482 178878 46718
rect 178962 46482 179198 46718
rect 179282 46482 179518 46718
rect 179602 46482 179838 46718
rect 179922 46482 180158 46718
rect 180242 46482 180478 46718
rect 180562 46482 180798 46718
rect 180882 46482 181118 46718
rect 181202 46482 181438 46718
rect 181522 46482 181758 46718
rect 181842 46482 182078 46718
rect 182162 46482 182398 46718
rect 182482 46482 182718 46718
rect 182802 46482 183038 46718
rect 183122 46482 183358 46718
rect 183442 46482 183678 46718
rect 183762 46482 183998 46718
rect 184082 46482 184318 46718
rect 184402 46482 184638 46718
rect 184722 46482 184958 46718
rect 187042 46482 187278 46718
rect 187362 46482 187598 46718
rect 187682 46482 187918 46718
rect 188002 46482 188238 46718
rect 188322 46482 188558 46718
rect 188642 46482 188878 46718
rect 188962 46482 189198 46718
rect 189282 46482 189518 46718
rect 189602 46482 189838 46718
rect 189922 46482 190158 46718
rect 190242 46482 190478 46718
rect 190562 46482 190798 46718
rect 190882 46482 191118 46718
rect 191202 46482 191438 46718
rect 191522 46482 191758 46718
rect 191842 46482 192078 46718
rect 192162 46482 192398 46718
rect 192482 46482 192718 46718
rect 192802 46482 193038 46718
rect 193122 46482 193358 46718
rect 193442 46482 193678 46718
rect 193762 46482 193998 46718
rect 194082 46482 194318 46718
rect 194402 46482 194638 46718
rect 194722 46482 194958 46718
rect 197042 46482 197278 46718
rect 197362 46482 197598 46718
rect 197682 46482 197918 46718
rect 198002 46482 198238 46718
rect 198322 46482 198558 46718
rect 198642 46482 198878 46718
rect 198962 46482 199198 46718
rect 199282 46482 199518 46718
rect 199602 46482 199838 46718
rect 199922 46482 200158 46718
rect 200242 46482 200478 46718
rect 200562 46482 200798 46718
rect 200882 46482 201118 46718
rect 201202 46482 201438 46718
rect 201522 46482 201758 46718
rect 201842 46482 202078 46718
rect 202162 46482 202398 46718
rect 202482 46482 202718 46718
rect 202802 46482 203038 46718
rect 203122 46482 203358 46718
rect 203442 46482 203678 46718
rect 203762 46482 203998 46718
rect 204082 46482 204318 46718
rect 204402 46482 204638 46718
rect 204722 46482 204958 46718
rect 207042 46482 207278 46718
rect 207362 46482 207598 46718
rect 207682 46482 207918 46718
rect 208002 46482 208238 46718
rect 208322 46482 208558 46718
rect 208642 46482 208878 46718
rect 208962 46482 209198 46718
rect 209282 46482 209518 46718
rect 209602 46482 209838 46718
rect 209922 46482 210158 46718
rect 210242 46482 210478 46718
rect 210562 46482 210798 46718
rect 210882 46482 211118 46718
rect 211202 46482 211438 46718
rect 211522 46482 211758 46718
rect 211842 46482 212078 46718
rect 212162 46482 212398 46718
rect 212482 46482 212718 46718
rect 212802 46482 213038 46718
rect 213122 46482 213358 46718
rect 213442 46482 213678 46718
rect 213762 46482 213998 46718
rect 214082 46482 214318 46718
rect 214402 46482 214638 46718
rect 214722 46482 214958 46718
rect 217042 46482 217278 46718
rect 217362 46482 217598 46718
rect 217682 46482 217918 46718
rect 218002 46482 218238 46718
rect 218322 46482 218558 46718
rect 218642 46482 218878 46718
rect 218962 46482 219198 46718
rect 219282 46482 219518 46718
rect 219602 46482 219838 46718
rect 219922 46482 220158 46718
rect 220242 46482 220478 46718
rect 220562 46482 220798 46718
rect 220882 46482 221118 46718
rect 221202 46482 221438 46718
rect 221522 46482 221758 46718
rect 221842 46482 222078 46718
rect 222162 46482 222398 46718
rect 222482 46482 222718 46718
rect 222802 46482 223038 46718
rect 223122 46482 223358 46718
rect 223442 46482 223678 46718
rect 223762 46482 223998 46718
rect 224082 46482 224318 46718
rect 224402 46482 224638 46718
rect 224722 46482 224958 46718
rect 227042 46482 227278 46718
rect 227362 46482 227598 46718
rect 227682 46482 227918 46718
rect 228002 46482 228238 46718
rect 228322 46482 228558 46718
rect 228642 46482 228878 46718
rect 228962 46482 229198 46718
rect 229282 46482 229518 46718
rect 229602 46482 229838 46718
rect 229922 46482 230158 46718
rect 230242 46482 230478 46718
rect 230562 46482 230798 46718
rect 230882 46482 231118 46718
rect 231202 46482 231438 46718
rect 231522 46482 231758 46718
rect 231842 46482 232078 46718
rect 232162 46482 232398 46718
rect 232482 46482 232718 46718
rect 232802 46482 233038 46718
rect 233122 46482 233358 46718
rect 233442 46482 233678 46718
rect 233762 46482 233998 46718
rect 234082 46482 234318 46718
rect 234402 46482 234638 46718
rect 234722 46482 234958 46718
rect 237042 46482 237278 46718
rect 237362 46482 237598 46718
rect 237682 46482 237918 46718
rect 238002 46482 238238 46718
rect 238322 46482 238558 46718
rect 238642 46482 238878 46718
rect 238962 46482 239198 46718
rect 239282 46482 239518 46718
rect 239602 46482 239838 46718
rect 239922 46482 240158 46718
rect 240242 46482 240478 46718
rect 240562 46482 240798 46718
rect 240882 46482 241118 46718
rect 241202 46482 241438 46718
rect 241522 46482 241758 46718
rect 241842 46482 242078 46718
rect 242162 46482 242398 46718
rect 242482 46482 242718 46718
rect 242802 46482 243038 46718
rect 243122 46482 243358 46718
rect 243442 46482 243678 46718
rect 243762 46482 243998 46718
rect 244082 46482 244318 46718
rect 244402 46482 244638 46718
rect 244722 46482 244958 46718
rect 247042 46482 247278 46718
rect 247362 46482 247598 46718
rect 247682 46482 247918 46718
rect 248002 46482 248238 46718
rect 248322 46482 248558 46718
rect 248642 46482 248878 46718
rect 248962 46482 249198 46718
rect 249282 46482 249518 46718
rect 249602 46482 249838 46718
rect 249922 46482 250158 46718
rect 250242 46482 250478 46718
rect 250562 46482 250798 46718
rect 250882 46482 251118 46718
rect 251202 46482 251438 46718
rect 251522 46482 251758 46718
rect 251842 46482 252078 46718
rect 252162 46482 252398 46718
rect 252482 46482 252718 46718
rect 252802 46482 253038 46718
rect 253122 46482 253358 46718
rect 253442 46482 253678 46718
rect 253762 46482 253998 46718
rect 254082 46482 254318 46718
rect 254402 46482 254638 46718
rect 254722 46482 254958 46718
rect 257042 46482 257278 46718
rect 257362 46482 257598 46718
rect 257682 46482 257918 46718
rect 258002 46482 258238 46718
rect 258322 46482 258558 46718
rect 258642 46482 258878 46718
rect 258962 46482 259198 46718
rect 259282 46482 259518 46718
rect 259602 46482 259838 46718
rect 259922 46482 260158 46718
rect 260242 46482 260478 46718
rect 260562 46482 260798 46718
rect 260882 46482 261118 46718
rect 261202 46482 261438 46718
rect 261522 46482 261758 46718
rect 261842 46482 262078 46718
rect 262162 46482 262398 46718
rect 262482 46482 262718 46718
rect 262802 46482 263038 46718
rect 263122 46482 263358 46718
rect 263442 46482 263678 46718
rect 263762 46482 263998 46718
rect 264082 46482 264318 46718
rect 264402 46482 264638 46718
rect 264722 46482 264958 46718
rect 267042 46482 267278 46718
rect 267362 46482 267598 46718
rect 267682 46482 267918 46718
rect 268002 46482 268238 46718
rect 268322 46482 268558 46718
rect 268642 46482 268878 46718
rect 268962 46482 269198 46718
rect 269282 46482 269518 46718
rect 269602 46482 269838 46718
rect 269922 46482 270158 46718
rect 270242 46482 270478 46718
rect 270562 46482 270798 46718
rect 270882 46482 271118 46718
rect 271202 46482 271438 46718
rect 271522 46482 271758 46718
rect 271842 46482 272078 46718
rect 272162 46482 272398 46718
rect 272482 46482 272718 46718
rect 272802 46482 273038 46718
rect 273122 46482 273358 46718
rect 273442 46482 273678 46718
rect 273762 46482 273998 46718
rect 274082 46482 274318 46718
rect 274402 46482 274638 46718
rect 274722 46482 274958 46718
rect 277042 46482 277278 46718
rect 277362 46482 277598 46718
rect 277682 46482 277918 46718
rect 278002 46482 278238 46718
rect 278322 46482 278558 46718
rect 278642 46482 278878 46718
rect 278962 46482 279198 46718
rect 279282 46482 279518 46718
rect 279602 46482 279838 46718
rect 279922 46482 280158 46718
rect 280242 46482 280478 46718
rect 280562 46482 280798 46718
rect 280882 46482 281118 46718
rect 281202 46482 281438 46718
rect 281522 46482 281758 46718
rect 281842 46482 282078 46718
rect 282162 46482 282398 46718
rect 282482 46482 282718 46718
rect 282802 46482 283038 46718
rect 283122 46482 283358 46718
rect 283442 46482 283678 46718
rect 283762 46482 283998 46718
rect 284082 46482 284318 46718
rect 284402 46482 284638 46718
rect 284722 46482 284958 46718
rect 44062 25822 44938 26378
rect 44062 5622 44938 6178
rect 47042 5282 47278 5518
rect 47362 5282 47598 5518
rect 47682 5282 47918 5518
rect 48002 5282 48238 5518
rect 48322 5282 48558 5518
rect 48642 5282 48878 5518
rect 48962 5282 49198 5518
rect 49282 5282 49518 5518
rect 49602 5282 49838 5518
rect 49922 5282 50158 5518
rect 50242 5282 50478 5518
rect 50562 5282 50798 5518
rect 50882 5282 51118 5518
rect 51202 5282 51438 5518
rect 51522 5282 51758 5518
rect 51842 5282 52078 5518
rect 52162 5282 52398 5518
rect 52482 5282 52718 5518
rect 52802 5282 53038 5518
rect 53122 5282 53358 5518
rect 53442 5282 53678 5518
rect 53762 5282 53998 5518
rect 54082 5282 54318 5518
rect 54402 5282 54638 5518
rect 54722 5282 54958 5518
rect 57042 5282 57278 5518
rect 57362 5282 57598 5518
rect 57682 5282 57918 5518
rect 58002 5282 58238 5518
rect 58322 5282 58558 5518
rect 58642 5282 58878 5518
rect 58962 5282 59198 5518
rect 59282 5282 59518 5518
rect 59602 5282 59838 5518
rect 59922 5282 60158 5518
rect 60242 5282 60478 5518
rect 60562 5282 60798 5518
rect 60882 5282 61118 5518
rect 61202 5282 61438 5518
rect 61522 5282 61758 5518
rect 61842 5282 62078 5518
rect 62162 5282 62398 5518
rect 62482 5282 62718 5518
rect 62802 5282 63038 5518
rect 63122 5282 63358 5518
rect 63442 5282 63678 5518
rect 63762 5282 63998 5518
rect 64082 5282 64318 5518
rect 64402 5282 64638 5518
rect 64722 5282 64958 5518
rect 67042 5282 67278 5518
rect 67362 5282 67598 5518
rect 67682 5282 67918 5518
rect 68002 5282 68238 5518
rect 68322 5282 68558 5518
rect 68642 5282 68878 5518
rect 68962 5282 69198 5518
rect 69282 5282 69518 5518
rect 69602 5282 69838 5518
rect 69922 5282 70158 5518
rect 70242 5282 70478 5518
rect 70562 5282 70798 5518
rect 70882 5282 71118 5518
rect 71202 5282 71438 5518
rect 71522 5282 71758 5518
rect 71842 5282 72078 5518
rect 72162 5282 72398 5518
rect 72482 5282 72718 5518
rect 72802 5282 73038 5518
rect 73122 5282 73358 5518
rect 73442 5282 73678 5518
rect 73762 5282 73998 5518
rect 74082 5282 74318 5518
rect 74402 5282 74638 5518
rect 74722 5282 74958 5518
rect 77042 5282 77278 5518
rect 77362 5282 77598 5518
rect 77682 5282 77918 5518
rect 78002 5282 78238 5518
rect 78322 5282 78558 5518
rect 78642 5282 78878 5518
rect 78962 5282 79198 5518
rect 79282 5282 79518 5518
rect 79602 5282 79838 5518
rect 79922 5282 80158 5518
rect 80242 5282 80478 5518
rect 80562 5282 80798 5518
rect 80882 5282 81118 5518
rect 81202 5282 81438 5518
rect 81522 5282 81758 5518
rect 81842 5282 82078 5518
rect 82162 5282 82398 5518
rect 82482 5282 82718 5518
rect 82802 5282 83038 5518
rect 83122 5282 83358 5518
rect 83442 5282 83678 5518
rect 83762 5282 83998 5518
rect 84082 5282 84318 5518
rect 84402 5282 84638 5518
rect 84722 5282 84958 5518
rect 87042 5282 87278 5518
rect 87362 5282 87598 5518
rect 87682 5282 87918 5518
rect 88002 5282 88238 5518
rect 88322 5282 88558 5518
rect 88642 5282 88878 5518
rect 88962 5282 89198 5518
rect 89282 5282 89518 5518
rect 89602 5282 89838 5518
rect 89922 5282 90158 5518
rect 90242 5282 90478 5518
rect 90562 5282 90798 5518
rect 90882 5282 91118 5518
rect 91202 5282 91438 5518
rect 91522 5282 91758 5518
rect 91842 5282 92078 5518
rect 92162 5282 92398 5518
rect 92482 5282 92718 5518
rect 92802 5282 93038 5518
rect 93122 5282 93358 5518
rect 93442 5282 93678 5518
rect 93762 5282 93998 5518
rect 94082 5282 94318 5518
rect 94402 5282 94638 5518
rect 94722 5282 94958 5518
rect 97042 5282 97278 5518
rect 97362 5282 97598 5518
rect 97682 5282 97918 5518
rect 98002 5282 98238 5518
rect 98322 5282 98558 5518
rect 98642 5282 98878 5518
rect 98962 5282 99198 5518
rect 99282 5282 99518 5518
rect 99602 5282 99838 5518
rect 99922 5282 100158 5518
rect 100242 5282 100478 5518
rect 100562 5282 100798 5518
rect 100882 5282 101118 5518
rect 101202 5282 101438 5518
rect 101522 5282 101758 5518
rect 101842 5282 102078 5518
rect 102162 5282 102398 5518
rect 102482 5282 102718 5518
rect 102802 5282 103038 5518
rect 103122 5282 103358 5518
rect 103442 5282 103678 5518
rect 103762 5282 103998 5518
rect 104082 5282 104318 5518
rect 104402 5282 104638 5518
rect 104722 5282 104958 5518
rect 107042 5282 107278 5518
rect 107362 5282 107598 5518
rect 107682 5282 107918 5518
rect 108002 5282 108238 5518
rect 108322 5282 108558 5518
rect 108642 5282 108878 5518
rect 108962 5282 109198 5518
rect 109282 5282 109518 5518
rect 109602 5282 109838 5518
rect 109922 5282 110158 5518
rect 110242 5282 110478 5518
rect 110562 5282 110798 5518
rect 110882 5282 111118 5518
rect 111202 5282 111438 5518
rect 111522 5282 111758 5518
rect 111842 5282 112078 5518
rect 112162 5282 112398 5518
rect 112482 5282 112718 5518
rect 112802 5282 113038 5518
rect 113122 5282 113358 5518
rect 113442 5282 113678 5518
rect 113762 5282 113998 5518
rect 114082 5282 114318 5518
rect 114402 5282 114638 5518
rect 114722 5282 114958 5518
rect 117042 5282 117278 5518
rect 117362 5282 117598 5518
rect 117682 5282 117918 5518
rect 118002 5282 118238 5518
rect 118322 5282 118558 5518
rect 118642 5282 118878 5518
rect 118962 5282 119198 5518
rect 119282 5282 119518 5518
rect 119602 5282 119838 5518
rect 119922 5282 120158 5518
rect 120242 5282 120478 5518
rect 120562 5282 120798 5518
rect 120882 5282 121118 5518
rect 121202 5282 121438 5518
rect 121522 5282 121758 5518
rect 121842 5282 122078 5518
rect 122162 5282 122398 5518
rect 122482 5282 122718 5518
rect 122802 5282 123038 5518
rect 123122 5282 123358 5518
rect 123442 5282 123678 5518
rect 123762 5282 123998 5518
rect 124082 5282 124318 5518
rect 124402 5282 124638 5518
rect 124722 5282 124958 5518
rect 127042 5282 127278 5518
rect 127362 5282 127598 5518
rect 127682 5282 127918 5518
rect 128002 5282 128238 5518
rect 128322 5282 128558 5518
rect 128642 5282 128878 5518
rect 128962 5282 129198 5518
rect 129282 5282 129518 5518
rect 129602 5282 129838 5518
rect 129922 5282 130158 5518
rect 130242 5282 130478 5518
rect 130562 5282 130798 5518
rect 130882 5282 131118 5518
rect 131202 5282 131438 5518
rect 131522 5282 131758 5518
rect 131842 5282 132078 5518
rect 132162 5282 132398 5518
rect 132482 5282 132718 5518
rect 132802 5282 133038 5518
rect 133122 5282 133358 5518
rect 133442 5282 133678 5518
rect 133762 5282 133998 5518
rect 134082 5282 134318 5518
rect 134402 5282 134638 5518
rect 134722 5282 134958 5518
rect 137042 5282 137278 5518
rect 137362 5282 137598 5518
rect 137682 5282 137918 5518
rect 138002 5282 138238 5518
rect 138322 5282 138558 5518
rect 138642 5282 138878 5518
rect 138962 5282 139198 5518
rect 139282 5282 139518 5518
rect 139602 5282 139838 5518
rect 139922 5282 140158 5518
rect 140242 5282 140478 5518
rect 140562 5282 140798 5518
rect 140882 5282 141118 5518
rect 141202 5282 141438 5518
rect 141522 5282 141758 5518
rect 141842 5282 142078 5518
rect 142162 5282 142398 5518
rect 142482 5282 142718 5518
rect 142802 5282 143038 5518
rect 143122 5282 143358 5518
rect 143442 5282 143678 5518
rect 143762 5282 143998 5518
rect 144082 5282 144318 5518
rect 144402 5282 144638 5518
rect 144722 5282 144958 5518
rect 147042 5282 147278 5518
rect 147362 5282 147598 5518
rect 147682 5282 147918 5518
rect 148002 5282 148238 5518
rect 148322 5282 148558 5518
rect 148642 5282 148878 5518
rect 148962 5282 149198 5518
rect 149282 5282 149518 5518
rect 149602 5282 149838 5518
rect 149922 5282 150158 5518
rect 150242 5282 150478 5518
rect 150562 5282 150798 5518
rect 150882 5282 151118 5518
rect 151202 5282 151438 5518
rect 151522 5282 151758 5518
rect 151842 5282 152078 5518
rect 152162 5282 152398 5518
rect 152482 5282 152718 5518
rect 152802 5282 153038 5518
rect 153122 5282 153358 5518
rect 153442 5282 153678 5518
rect 153762 5282 153998 5518
rect 154082 5282 154318 5518
rect 154402 5282 154638 5518
rect 154722 5282 154958 5518
rect 157042 5282 157278 5518
rect 157362 5282 157598 5518
rect 157682 5282 157918 5518
rect 158002 5282 158238 5518
rect 158322 5282 158558 5518
rect 158642 5282 158878 5518
rect 158962 5282 159198 5518
rect 159282 5282 159518 5518
rect 159602 5282 159838 5518
rect 159922 5282 160158 5518
rect 160242 5282 160478 5518
rect 160562 5282 160798 5518
rect 160882 5282 161118 5518
rect 161202 5282 161438 5518
rect 161522 5282 161758 5518
rect 161842 5282 162078 5518
rect 162162 5282 162398 5518
rect 162482 5282 162718 5518
rect 162802 5282 163038 5518
rect 163122 5282 163358 5518
rect 163442 5282 163678 5518
rect 163762 5282 163998 5518
rect 164082 5282 164318 5518
rect 164402 5282 164638 5518
rect 164722 5282 164958 5518
rect 167042 5282 167278 5518
rect 167362 5282 167598 5518
rect 167682 5282 167918 5518
rect 168002 5282 168238 5518
rect 168322 5282 168558 5518
rect 168642 5282 168878 5518
rect 168962 5282 169198 5518
rect 169282 5282 169518 5518
rect 169602 5282 169838 5518
rect 169922 5282 170158 5518
rect 170242 5282 170478 5518
rect 170562 5282 170798 5518
rect 170882 5282 171118 5518
rect 171202 5282 171438 5518
rect 171522 5282 171758 5518
rect 171842 5282 172078 5518
rect 172162 5282 172398 5518
rect 172482 5282 172718 5518
rect 172802 5282 173038 5518
rect 173122 5282 173358 5518
rect 173442 5282 173678 5518
rect 173762 5282 173998 5518
rect 174082 5282 174318 5518
rect 174402 5282 174638 5518
rect 174722 5282 174958 5518
rect 177042 5282 177278 5518
rect 177362 5282 177598 5518
rect 177682 5282 177918 5518
rect 178002 5282 178238 5518
rect 178322 5282 178558 5518
rect 178642 5282 178878 5518
rect 178962 5282 179198 5518
rect 179282 5282 179518 5518
rect 179602 5282 179838 5518
rect 179922 5282 180158 5518
rect 180242 5282 180478 5518
rect 180562 5282 180798 5518
rect 180882 5282 181118 5518
rect 181202 5282 181438 5518
rect 181522 5282 181758 5518
rect 181842 5282 182078 5518
rect 182162 5282 182398 5518
rect 182482 5282 182718 5518
rect 182802 5282 183038 5518
rect 183122 5282 183358 5518
rect 183442 5282 183678 5518
rect 183762 5282 183998 5518
rect 184082 5282 184318 5518
rect 184402 5282 184638 5518
rect 184722 5282 184958 5518
rect 187042 5282 187278 5518
rect 187362 5282 187598 5518
rect 187682 5282 187918 5518
rect 188002 5282 188238 5518
rect 188322 5282 188558 5518
rect 188642 5282 188878 5518
rect 188962 5282 189198 5518
rect 189282 5282 189518 5518
rect 189602 5282 189838 5518
rect 189922 5282 190158 5518
rect 190242 5282 190478 5518
rect 190562 5282 190798 5518
rect 190882 5282 191118 5518
rect 191202 5282 191438 5518
rect 191522 5282 191758 5518
rect 191842 5282 192078 5518
rect 192162 5282 192398 5518
rect 192482 5282 192718 5518
rect 192802 5282 193038 5518
rect 193122 5282 193358 5518
rect 193442 5282 193678 5518
rect 193762 5282 193998 5518
rect 194082 5282 194318 5518
rect 194402 5282 194638 5518
rect 194722 5282 194958 5518
rect 197042 5282 197278 5518
rect 197362 5282 197598 5518
rect 197682 5282 197918 5518
rect 198002 5282 198238 5518
rect 198322 5282 198558 5518
rect 198642 5282 198878 5518
rect 198962 5282 199198 5518
rect 199282 5282 199518 5518
rect 199602 5282 199838 5518
rect 199922 5282 200158 5518
rect 200242 5282 200478 5518
rect 200562 5282 200798 5518
rect 200882 5282 201118 5518
rect 201202 5282 201438 5518
rect 201522 5282 201758 5518
rect 201842 5282 202078 5518
rect 202162 5282 202398 5518
rect 202482 5282 202718 5518
rect 202802 5282 203038 5518
rect 203122 5282 203358 5518
rect 203442 5282 203678 5518
rect 203762 5282 203998 5518
rect 204082 5282 204318 5518
rect 204402 5282 204638 5518
rect 204722 5282 204958 5518
rect 207042 5282 207278 5518
rect 207362 5282 207598 5518
rect 207682 5282 207918 5518
rect 208002 5282 208238 5518
rect 208322 5282 208558 5518
rect 208642 5282 208878 5518
rect 208962 5282 209198 5518
rect 209282 5282 209518 5518
rect 209602 5282 209838 5518
rect 209922 5282 210158 5518
rect 210242 5282 210478 5518
rect 210562 5282 210798 5518
rect 210882 5282 211118 5518
rect 211202 5282 211438 5518
rect 211522 5282 211758 5518
rect 211842 5282 212078 5518
rect 212162 5282 212398 5518
rect 212482 5282 212718 5518
rect 212802 5282 213038 5518
rect 213122 5282 213358 5518
rect 213442 5282 213678 5518
rect 213762 5282 213998 5518
rect 214082 5282 214318 5518
rect 214402 5282 214638 5518
rect 214722 5282 214958 5518
rect 217042 5282 217278 5518
rect 217362 5282 217598 5518
rect 217682 5282 217918 5518
rect 218002 5282 218238 5518
rect 218322 5282 218558 5518
rect 218642 5282 218878 5518
rect 218962 5282 219198 5518
rect 219282 5282 219518 5518
rect 219602 5282 219838 5518
rect 219922 5282 220158 5518
rect 220242 5282 220478 5518
rect 220562 5282 220798 5518
rect 220882 5282 221118 5518
rect 221202 5282 221438 5518
rect 221522 5282 221758 5518
rect 221842 5282 222078 5518
rect 222162 5282 222398 5518
rect 222482 5282 222718 5518
rect 222802 5282 223038 5518
rect 223122 5282 223358 5518
rect 223442 5282 223678 5518
rect 223762 5282 223998 5518
rect 224082 5282 224318 5518
rect 224402 5282 224638 5518
rect 224722 5282 224958 5518
rect 227042 5282 227278 5518
rect 227362 5282 227598 5518
rect 227682 5282 227918 5518
rect 228002 5282 228238 5518
rect 228322 5282 228558 5518
rect 228642 5282 228878 5518
rect 228962 5282 229198 5518
rect 229282 5282 229518 5518
rect 229602 5282 229838 5518
rect 229922 5282 230158 5518
rect 230242 5282 230478 5518
rect 230562 5282 230798 5518
rect 230882 5282 231118 5518
rect 231202 5282 231438 5518
rect 231522 5282 231758 5518
rect 231842 5282 232078 5518
rect 232162 5282 232398 5518
rect 232482 5282 232718 5518
rect 232802 5282 233038 5518
rect 233122 5282 233358 5518
rect 233442 5282 233678 5518
rect 233762 5282 233998 5518
rect 234082 5282 234318 5518
rect 234402 5282 234638 5518
rect 234722 5282 234958 5518
rect 237042 5282 237278 5518
rect 237362 5282 237598 5518
rect 237682 5282 237918 5518
rect 238002 5282 238238 5518
rect 238322 5282 238558 5518
rect 238642 5282 238878 5518
rect 238962 5282 239198 5518
rect 239282 5282 239518 5518
rect 239602 5282 239838 5518
rect 239922 5282 240158 5518
rect 240242 5282 240478 5518
rect 240562 5282 240798 5518
rect 240882 5282 241118 5518
rect 241202 5282 241438 5518
rect 241522 5282 241758 5518
rect 241842 5282 242078 5518
rect 242162 5282 242398 5518
rect 242482 5282 242718 5518
rect 242802 5282 243038 5518
rect 243122 5282 243358 5518
rect 243442 5282 243678 5518
rect 243762 5282 243998 5518
rect 244082 5282 244318 5518
rect 244402 5282 244638 5518
rect 244722 5282 244958 5518
rect 247042 5282 247278 5518
rect 247362 5282 247598 5518
rect 247682 5282 247918 5518
rect 248002 5282 248238 5518
rect 248322 5282 248558 5518
rect 248642 5282 248878 5518
rect 248962 5282 249198 5518
rect 249282 5282 249518 5518
rect 249602 5282 249838 5518
rect 249922 5282 250158 5518
rect 250242 5282 250478 5518
rect 250562 5282 250798 5518
rect 250882 5282 251118 5518
rect 251202 5282 251438 5518
rect 251522 5282 251758 5518
rect 251842 5282 252078 5518
rect 252162 5282 252398 5518
rect 252482 5282 252718 5518
rect 252802 5282 253038 5518
rect 253122 5282 253358 5518
rect 253442 5282 253678 5518
rect 253762 5282 253998 5518
rect 254082 5282 254318 5518
rect 254402 5282 254638 5518
rect 254722 5282 254958 5518
rect 257042 5282 257278 5518
rect 257362 5282 257598 5518
rect 257682 5282 257918 5518
rect 258002 5282 258238 5518
rect 258322 5282 258558 5518
rect 258642 5282 258878 5518
rect 258962 5282 259198 5518
rect 259282 5282 259518 5518
rect 259602 5282 259838 5518
rect 259922 5282 260158 5518
rect 260242 5282 260478 5518
rect 260562 5282 260798 5518
rect 260882 5282 261118 5518
rect 261202 5282 261438 5518
rect 261522 5282 261758 5518
rect 261842 5282 262078 5518
rect 262162 5282 262398 5518
rect 262482 5282 262718 5518
rect 262802 5282 263038 5518
rect 263122 5282 263358 5518
rect 263442 5282 263678 5518
rect 263762 5282 263998 5518
rect 264082 5282 264318 5518
rect 264402 5282 264638 5518
rect 264722 5282 264958 5518
rect 267042 5282 267278 5518
rect 267362 5282 267598 5518
rect 267682 5282 267918 5518
rect 268002 5282 268238 5518
rect 268322 5282 268558 5518
rect 268642 5282 268878 5518
rect 268962 5282 269198 5518
rect 269282 5282 269518 5518
rect 269602 5282 269838 5518
rect 269922 5282 270158 5518
rect 270242 5282 270478 5518
rect 270562 5282 270798 5518
rect 270882 5282 271118 5518
rect 271202 5282 271438 5518
rect 271522 5282 271758 5518
rect 271842 5282 272078 5518
rect 272162 5282 272398 5518
rect 272482 5282 272718 5518
rect 272802 5282 273038 5518
rect 273122 5282 273358 5518
rect 273442 5282 273678 5518
rect 273762 5282 273998 5518
rect 274082 5282 274318 5518
rect 274402 5282 274638 5518
rect 274722 5282 274958 5518
rect 277042 5282 277278 5518
rect 277362 5282 277598 5518
rect 277682 5282 277918 5518
rect 278002 5282 278238 5518
rect 278322 5282 278558 5518
rect 278642 5282 278878 5518
rect 278962 5282 279198 5518
rect 279282 5282 279518 5518
rect 279602 5282 279838 5518
rect 279922 5282 280158 5518
rect 280242 5282 280478 5518
rect 280562 5282 280798 5518
rect 280882 5282 281118 5518
rect 281202 5282 281438 5518
rect 281522 5282 281758 5518
rect 281842 5282 282078 5518
rect 282162 5282 282398 5518
rect 282482 5282 282718 5518
rect 282802 5282 283038 5518
rect 283122 5282 283358 5518
rect 283442 5282 283678 5518
rect 283762 5282 283998 5518
rect 284082 5282 284318 5518
rect 284402 5282 284638 5518
rect 284722 5282 284958 5518
<< mimcap2 >>
rect 46040 45818 54360 45960
rect 46040 26382 46082 45818
rect 54318 26382 54360 45818
rect 46040 26240 54360 26382
rect 56040 45818 64360 45960
rect 56040 26382 56082 45818
rect 64318 26382 64360 45818
rect 56040 26240 64360 26382
rect 66040 45818 74360 45960
rect 66040 26382 66082 45818
rect 74318 26382 74360 45818
rect 66040 26240 74360 26382
rect 76040 45818 84360 45960
rect 76040 26382 76082 45818
rect 84318 26382 84360 45818
rect 76040 26240 84360 26382
rect 86040 45818 94360 45960
rect 86040 26382 86082 45818
rect 94318 26382 94360 45818
rect 86040 26240 94360 26382
rect 96040 45818 104360 45960
rect 96040 26382 96082 45818
rect 104318 26382 104360 45818
rect 96040 26240 104360 26382
rect 106040 45818 114360 45960
rect 106040 26382 106082 45818
rect 114318 26382 114360 45818
rect 106040 26240 114360 26382
rect 116040 45818 124360 45960
rect 116040 26382 116082 45818
rect 124318 26382 124360 45818
rect 116040 26240 124360 26382
rect 126040 45818 134360 45960
rect 126040 26382 126082 45818
rect 134318 26382 134360 45818
rect 126040 26240 134360 26382
rect 136040 45818 144360 45960
rect 136040 26382 136082 45818
rect 144318 26382 144360 45818
rect 136040 26240 144360 26382
rect 146040 45818 154360 45960
rect 146040 26382 146082 45818
rect 154318 26382 154360 45818
rect 146040 26240 154360 26382
rect 156040 45818 164360 45960
rect 156040 26382 156082 45818
rect 164318 26382 164360 45818
rect 156040 26240 164360 26382
rect 166040 45818 174360 45960
rect 166040 26382 166082 45818
rect 174318 26382 174360 45818
rect 166040 26240 174360 26382
rect 176040 45818 184360 45960
rect 176040 26382 176082 45818
rect 184318 26382 184360 45818
rect 176040 26240 184360 26382
rect 186040 45818 194360 45960
rect 186040 26382 186082 45818
rect 194318 26382 194360 45818
rect 186040 26240 194360 26382
rect 196040 45818 204360 45960
rect 196040 26382 196082 45818
rect 204318 26382 204360 45818
rect 196040 26240 204360 26382
rect 206040 45818 214360 45960
rect 206040 26382 206082 45818
rect 214318 26382 214360 45818
rect 206040 26240 214360 26382
rect 216040 45818 224360 45960
rect 216040 26382 216082 45818
rect 224318 26382 224360 45818
rect 216040 26240 224360 26382
rect 226040 45818 234360 45960
rect 226040 26382 226082 45818
rect 234318 26382 234360 45818
rect 226040 26240 234360 26382
rect 236040 45818 244360 45960
rect 236040 26382 236082 45818
rect 244318 26382 244360 45818
rect 236040 26240 244360 26382
rect 246040 45818 254360 45960
rect 246040 26382 246082 45818
rect 254318 26382 254360 45818
rect 246040 26240 254360 26382
rect 256040 45818 264360 45960
rect 256040 26382 256082 45818
rect 264318 26382 264360 45818
rect 256040 26240 264360 26382
rect 266040 45818 274360 45960
rect 266040 26382 266082 45818
rect 274318 26382 274360 45818
rect 266040 26240 274360 26382
rect 276040 45818 284360 45960
rect 276040 26382 276082 45818
rect 284318 26382 284360 45818
rect 276040 26240 284360 26382
rect 47640 25618 55960 25760
rect 47640 6182 47682 25618
rect 55918 6182 55960 25618
rect 47640 6040 55960 6182
rect 57640 25618 65960 25760
rect 57640 6182 57682 25618
rect 65918 6182 65960 25618
rect 57640 6040 65960 6182
rect 67640 25618 75960 25760
rect 67640 6182 67682 25618
rect 75918 6182 75960 25618
rect 67640 6040 75960 6182
rect 77640 25618 85960 25760
rect 77640 6182 77682 25618
rect 85918 6182 85960 25618
rect 77640 6040 85960 6182
rect 87640 25618 95960 25760
rect 87640 6182 87682 25618
rect 95918 6182 95960 25618
rect 87640 6040 95960 6182
rect 97640 25618 105960 25760
rect 97640 6182 97682 25618
rect 105918 6182 105960 25618
rect 97640 6040 105960 6182
rect 107640 25618 115960 25760
rect 107640 6182 107682 25618
rect 115918 6182 115960 25618
rect 107640 6040 115960 6182
rect 117640 25618 125960 25760
rect 117640 6182 117682 25618
rect 125918 6182 125960 25618
rect 117640 6040 125960 6182
rect 127640 25618 135960 25760
rect 127640 6182 127682 25618
rect 135918 6182 135960 25618
rect 127640 6040 135960 6182
rect 137640 25618 145960 25760
rect 137640 6182 137682 25618
rect 145918 6182 145960 25618
rect 137640 6040 145960 6182
rect 147640 25618 155960 25760
rect 147640 6182 147682 25618
rect 155918 6182 155960 25618
rect 147640 6040 155960 6182
rect 157640 25618 165960 25760
rect 157640 6182 157682 25618
rect 165918 6182 165960 25618
rect 157640 6040 165960 6182
rect 167640 25618 175960 25760
rect 167640 6182 167682 25618
rect 175918 6182 175960 25618
rect 167640 6040 175960 6182
rect 177640 25618 185960 25760
rect 177640 6182 177682 25618
rect 185918 6182 185960 25618
rect 177640 6040 185960 6182
rect 187640 25618 195960 25760
rect 187640 6182 187682 25618
rect 195918 6182 195960 25618
rect 187640 6040 195960 6182
rect 197640 25618 205960 25760
rect 197640 6182 197682 25618
rect 205918 6182 205960 25618
rect 197640 6040 205960 6182
rect 207640 25618 215960 25760
rect 207640 6182 207682 25618
rect 215918 6182 215960 25618
rect 207640 6040 215960 6182
rect 217640 25618 225960 25760
rect 217640 6182 217682 25618
rect 225918 6182 225960 25618
rect 217640 6040 225960 6182
rect 227640 25618 235960 25760
rect 227640 6182 227682 25618
rect 235918 6182 235960 25618
rect 227640 6040 235960 6182
rect 237640 25618 245960 25760
rect 237640 6182 237682 25618
rect 245918 6182 245960 25618
rect 237640 6040 245960 6182
rect 247640 25618 255960 25760
rect 247640 6182 247682 25618
rect 255918 6182 255960 25618
rect 247640 6040 255960 6182
rect 257640 25618 265960 25760
rect 257640 6182 257682 25618
rect 265918 6182 265960 25618
rect 257640 6040 265960 6182
rect 267640 25618 275960 25760
rect 267640 6182 267682 25618
rect 275918 6182 275960 25618
rect 267640 6040 275960 6182
rect 277640 25618 285960 25760
rect 277640 6182 277682 25618
rect 285918 6182 285960 25618
rect 277640 6040 285960 6182
<< mimcap2contact >>
rect 46082 26382 54318 45818
rect 56082 26382 64318 45818
rect 66082 26382 74318 45818
rect 76082 26382 84318 45818
rect 86082 26382 94318 45818
rect 96082 26382 104318 45818
rect 106082 26382 114318 45818
rect 116082 26382 124318 45818
rect 126082 26382 134318 45818
rect 136082 26382 144318 45818
rect 146082 26382 154318 45818
rect 156082 26382 164318 45818
rect 166082 26382 174318 45818
rect 176082 26382 184318 45818
rect 186082 26382 194318 45818
rect 196082 26382 204318 45818
rect 206082 26382 214318 45818
rect 216082 26382 224318 45818
rect 226082 26382 234318 45818
rect 236082 26382 244318 45818
rect 246082 26382 254318 45818
rect 256082 26382 264318 45818
rect 266082 26382 274318 45818
rect 276082 26382 284318 45818
rect 47682 6182 55918 25618
rect 57682 6182 65918 25618
rect 67682 6182 75918 25618
rect 77682 6182 85918 25618
rect 87682 6182 95918 25618
rect 97682 6182 105918 25618
rect 107682 6182 115918 25618
rect 117682 6182 125918 25618
rect 127682 6182 135918 25618
rect 137682 6182 145918 25618
rect 147682 6182 155918 25618
rect 157682 6182 165918 25618
rect 167682 6182 175918 25618
rect 177682 6182 185918 25618
rect 187682 6182 195918 25618
rect 197682 6182 205918 25618
rect 207682 6182 215918 25618
rect 217682 6182 225918 25618
rect 227682 6182 235918 25618
rect 237682 6182 245918 25618
rect 247682 6182 255918 25618
rect 257682 6182 265918 25618
rect 267682 6182 275918 25618
rect 277682 6182 285918 25618
<< metal5 >>
rect 46000 46718 286000 46800
rect 46000 46482 47042 46718
rect 47278 46482 47362 46718
rect 47598 46482 47682 46718
rect 47918 46482 48002 46718
rect 48238 46482 48322 46718
rect 48558 46482 48642 46718
rect 48878 46482 48962 46718
rect 49198 46482 49282 46718
rect 49518 46482 49602 46718
rect 49838 46482 49922 46718
rect 50158 46482 50242 46718
rect 50478 46482 50562 46718
rect 50798 46482 50882 46718
rect 51118 46482 51202 46718
rect 51438 46482 51522 46718
rect 51758 46482 51842 46718
rect 52078 46482 52162 46718
rect 52398 46482 52482 46718
rect 52718 46482 52802 46718
rect 53038 46482 53122 46718
rect 53358 46482 53442 46718
rect 53678 46482 53762 46718
rect 53998 46482 54082 46718
rect 54318 46482 54402 46718
rect 54638 46482 54722 46718
rect 54958 46482 57042 46718
rect 57278 46482 57362 46718
rect 57598 46482 57682 46718
rect 57918 46482 58002 46718
rect 58238 46482 58322 46718
rect 58558 46482 58642 46718
rect 58878 46482 58962 46718
rect 59198 46482 59282 46718
rect 59518 46482 59602 46718
rect 59838 46482 59922 46718
rect 60158 46482 60242 46718
rect 60478 46482 60562 46718
rect 60798 46482 60882 46718
rect 61118 46482 61202 46718
rect 61438 46482 61522 46718
rect 61758 46482 61842 46718
rect 62078 46482 62162 46718
rect 62398 46482 62482 46718
rect 62718 46482 62802 46718
rect 63038 46482 63122 46718
rect 63358 46482 63442 46718
rect 63678 46482 63762 46718
rect 63998 46482 64082 46718
rect 64318 46482 64402 46718
rect 64638 46482 64722 46718
rect 64958 46482 67042 46718
rect 67278 46482 67362 46718
rect 67598 46482 67682 46718
rect 67918 46482 68002 46718
rect 68238 46482 68322 46718
rect 68558 46482 68642 46718
rect 68878 46482 68962 46718
rect 69198 46482 69282 46718
rect 69518 46482 69602 46718
rect 69838 46482 69922 46718
rect 70158 46482 70242 46718
rect 70478 46482 70562 46718
rect 70798 46482 70882 46718
rect 71118 46482 71202 46718
rect 71438 46482 71522 46718
rect 71758 46482 71842 46718
rect 72078 46482 72162 46718
rect 72398 46482 72482 46718
rect 72718 46482 72802 46718
rect 73038 46482 73122 46718
rect 73358 46482 73442 46718
rect 73678 46482 73762 46718
rect 73998 46482 74082 46718
rect 74318 46482 74402 46718
rect 74638 46482 74722 46718
rect 74958 46482 77042 46718
rect 77278 46482 77362 46718
rect 77598 46482 77682 46718
rect 77918 46482 78002 46718
rect 78238 46482 78322 46718
rect 78558 46482 78642 46718
rect 78878 46482 78962 46718
rect 79198 46482 79282 46718
rect 79518 46482 79602 46718
rect 79838 46482 79922 46718
rect 80158 46482 80242 46718
rect 80478 46482 80562 46718
rect 80798 46482 80882 46718
rect 81118 46482 81202 46718
rect 81438 46482 81522 46718
rect 81758 46482 81842 46718
rect 82078 46482 82162 46718
rect 82398 46482 82482 46718
rect 82718 46482 82802 46718
rect 83038 46482 83122 46718
rect 83358 46482 83442 46718
rect 83678 46482 83762 46718
rect 83998 46482 84082 46718
rect 84318 46482 84402 46718
rect 84638 46482 84722 46718
rect 84958 46482 87042 46718
rect 87278 46482 87362 46718
rect 87598 46482 87682 46718
rect 87918 46482 88002 46718
rect 88238 46482 88322 46718
rect 88558 46482 88642 46718
rect 88878 46482 88962 46718
rect 89198 46482 89282 46718
rect 89518 46482 89602 46718
rect 89838 46482 89922 46718
rect 90158 46482 90242 46718
rect 90478 46482 90562 46718
rect 90798 46482 90882 46718
rect 91118 46482 91202 46718
rect 91438 46482 91522 46718
rect 91758 46482 91842 46718
rect 92078 46482 92162 46718
rect 92398 46482 92482 46718
rect 92718 46482 92802 46718
rect 93038 46482 93122 46718
rect 93358 46482 93442 46718
rect 93678 46482 93762 46718
rect 93998 46482 94082 46718
rect 94318 46482 94402 46718
rect 94638 46482 94722 46718
rect 94958 46482 97042 46718
rect 97278 46482 97362 46718
rect 97598 46482 97682 46718
rect 97918 46482 98002 46718
rect 98238 46482 98322 46718
rect 98558 46482 98642 46718
rect 98878 46482 98962 46718
rect 99198 46482 99282 46718
rect 99518 46482 99602 46718
rect 99838 46482 99922 46718
rect 100158 46482 100242 46718
rect 100478 46482 100562 46718
rect 100798 46482 100882 46718
rect 101118 46482 101202 46718
rect 101438 46482 101522 46718
rect 101758 46482 101842 46718
rect 102078 46482 102162 46718
rect 102398 46482 102482 46718
rect 102718 46482 102802 46718
rect 103038 46482 103122 46718
rect 103358 46482 103442 46718
rect 103678 46482 103762 46718
rect 103998 46482 104082 46718
rect 104318 46482 104402 46718
rect 104638 46482 104722 46718
rect 104958 46482 107042 46718
rect 107278 46482 107362 46718
rect 107598 46482 107682 46718
rect 107918 46482 108002 46718
rect 108238 46482 108322 46718
rect 108558 46482 108642 46718
rect 108878 46482 108962 46718
rect 109198 46482 109282 46718
rect 109518 46482 109602 46718
rect 109838 46482 109922 46718
rect 110158 46482 110242 46718
rect 110478 46482 110562 46718
rect 110798 46482 110882 46718
rect 111118 46482 111202 46718
rect 111438 46482 111522 46718
rect 111758 46482 111842 46718
rect 112078 46482 112162 46718
rect 112398 46482 112482 46718
rect 112718 46482 112802 46718
rect 113038 46482 113122 46718
rect 113358 46482 113442 46718
rect 113678 46482 113762 46718
rect 113998 46482 114082 46718
rect 114318 46482 114402 46718
rect 114638 46482 114722 46718
rect 114958 46482 117042 46718
rect 117278 46482 117362 46718
rect 117598 46482 117682 46718
rect 117918 46482 118002 46718
rect 118238 46482 118322 46718
rect 118558 46482 118642 46718
rect 118878 46482 118962 46718
rect 119198 46482 119282 46718
rect 119518 46482 119602 46718
rect 119838 46482 119922 46718
rect 120158 46482 120242 46718
rect 120478 46482 120562 46718
rect 120798 46482 120882 46718
rect 121118 46482 121202 46718
rect 121438 46482 121522 46718
rect 121758 46482 121842 46718
rect 122078 46482 122162 46718
rect 122398 46482 122482 46718
rect 122718 46482 122802 46718
rect 123038 46482 123122 46718
rect 123358 46482 123442 46718
rect 123678 46482 123762 46718
rect 123998 46482 124082 46718
rect 124318 46482 124402 46718
rect 124638 46482 124722 46718
rect 124958 46482 127042 46718
rect 127278 46482 127362 46718
rect 127598 46482 127682 46718
rect 127918 46482 128002 46718
rect 128238 46482 128322 46718
rect 128558 46482 128642 46718
rect 128878 46482 128962 46718
rect 129198 46482 129282 46718
rect 129518 46482 129602 46718
rect 129838 46482 129922 46718
rect 130158 46482 130242 46718
rect 130478 46482 130562 46718
rect 130798 46482 130882 46718
rect 131118 46482 131202 46718
rect 131438 46482 131522 46718
rect 131758 46482 131842 46718
rect 132078 46482 132162 46718
rect 132398 46482 132482 46718
rect 132718 46482 132802 46718
rect 133038 46482 133122 46718
rect 133358 46482 133442 46718
rect 133678 46482 133762 46718
rect 133998 46482 134082 46718
rect 134318 46482 134402 46718
rect 134638 46482 134722 46718
rect 134958 46482 137042 46718
rect 137278 46482 137362 46718
rect 137598 46482 137682 46718
rect 137918 46482 138002 46718
rect 138238 46482 138322 46718
rect 138558 46482 138642 46718
rect 138878 46482 138962 46718
rect 139198 46482 139282 46718
rect 139518 46482 139602 46718
rect 139838 46482 139922 46718
rect 140158 46482 140242 46718
rect 140478 46482 140562 46718
rect 140798 46482 140882 46718
rect 141118 46482 141202 46718
rect 141438 46482 141522 46718
rect 141758 46482 141842 46718
rect 142078 46482 142162 46718
rect 142398 46482 142482 46718
rect 142718 46482 142802 46718
rect 143038 46482 143122 46718
rect 143358 46482 143442 46718
rect 143678 46482 143762 46718
rect 143998 46482 144082 46718
rect 144318 46482 144402 46718
rect 144638 46482 144722 46718
rect 144958 46482 147042 46718
rect 147278 46482 147362 46718
rect 147598 46482 147682 46718
rect 147918 46482 148002 46718
rect 148238 46482 148322 46718
rect 148558 46482 148642 46718
rect 148878 46482 148962 46718
rect 149198 46482 149282 46718
rect 149518 46482 149602 46718
rect 149838 46482 149922 46718
rect 150158 46482 150242 46718
rect 150478 46482 150562 46718
rect 150798 46482 150882 46718
rect 151118 46482 151202 46718
rect 151438 46482 151522 46718
rect 151758 46482 151842 46718
rect 152078 46482 152162 46718
rect 152398 46482 152482 46718
rect 152718 46482 152802 46718
rect 153038 46482 153122 46718
rect 153358 46482 153442 46718
rect 153678 46482 153762 46718
rect 153998 46482 154082 46718
rect 154318 46482 154402 46718
rect 154638 46482 154722 46718
rect 154958 46482 157042 46718
rect 157278 46482 157362 46718
rect 157598 46482 157682 46718
rect 157918 46482 158002 46718
rect 158238 46482 158322 46718
rect 158558 46482 158642 46718
rect 158878 46482 158962 46718
rect 159198 46482 159282 46718
rect 159518 46482 159602 46718
rect 159838 46482 159922 46718
rect 160158 46482 160242 46718
rect 160478 46482 160562 46718
rect 160798 46482 160882 46718
rect 161118 46482 161202 46718
rect 161438 46482 161522 46718
rect 161758 46482 161842 46718
rect 162078 46482 162162 46718
rect 162398 46482 162482 46718
rect 162718 46482 162802 46718
rect 163038 46482 163122 46718
rect 163358 46482 163442 46718
rect 163678 46482 163762 46718
rect 163998 46482 164082 46718
rect 164318 46482 164402 46718
rect 164638 46482 164722 46718
rect 164958 46482 167042 46718
rect 167278 46482 167362 46718
rect 167598 46482 167682 46718
rect 167918 46482 168002 46718
rect 168238 46482 168322 46718
rect 168558 46482 168642 46718
rect 168878 46482 168962 46718
rect 169198 46482 169282 46718
rect 169518 46482 169602 46718
rect 169838 46482 169922 46718
rect 170158 46482 170242 46718
rect 170478 46482 170562 46718
rect 170798 46482 170882 46718
rect 171118 46482 171202 46718
rect 171438 46482 171522 46718
rect 171758 46482 171842 46718
rect 172078 46482 172162 46718
rect 172398 46482 172482 46718
rect 172718 46482 172802 46718
rect 173038 46482 173122 46718
rect 173358 46482 173442 46718
rect 173678 46482 173762 46718
rect 173998 46482 174082 46718
rect 174318 46482 174402 46718
rect 174638 46482 174722 46718
rect 174958 46482 177042 46718
rect 177278 46482 177362 46718
rect 177598 46482 177682 46718
rect 177918 46482 178002 46718
rect 178238 46482 178322 46718
rect 178558 46482 178642 46718
rect 178878 46482 178962 46718
rect 179198 46482 179282 46718
rect 179518 46482 179602 46718
rect 179838 46482 179922 46718
rect 180158 46482 180242 46718
rect 180478 46482 180562 46718
rect 180798 46482 180882 46718
rect 181118 46482 181202 46718
rect 181438 46482 181522 46718
rect 181758 46482 181842 46718
rect 182078 46482 182162 46718
rect 182398 46482 182482 46718
rect 182718 46482 182802 46718
rect 183038 46482 183122 46718
rect 183358 46482 183442 46718
rect 183678 46482 183762 46718
rect 183998 46482 184082 46718
rect 184318 46482 184402 46718
rect 184638 46482 184722 46718
rect 184958 46482 187042 46718
rect 187278 46482 187362 46718
rect 187598 46482 187682 46718
rect 187918 46482 188002 46718
rect 188238 46482 188322 46718
rect 188558 46482 188642 46718
rect 188878 46482 188962 46718
rect 189198 46482 189282 46718
rect 189518 46482 189602 46718
rect 189838 46482 189922 46718
rect 190158 46482 190242 46718
rect 190478 46482 190562 46718
rect 190798 46482 190882 46718
rect 191118 46482 191202 46718
rect 191438 46482 191522 46718
rect 191758 46482 191842 46718
rect 192078 46482 192162 46718
rect 192398 46482 192482 46718
rect 192718 46482 192802 46718
rect 193038 46482 193122 46718
rect 193358 46482 193442 46718
rect 193678 46482 193762 46718
rect 193998 46482 194082 46718
rect 194318 46482 194402 46718
rect 194638 46482 194722 46718
rect 194958 46482 197042 46718
rect 197278 46482 197362 46718
rect 197598 46482 197682 46718
rect 197918 46482 198002 46718
rect 198238 46482 198322 46718
rect 198558 46482 198642 46718
rect 198878 46482 198962 46718
rect 199198 46482 199282 46718
rect 199518 46482 199602 46718
rect 199838 46482 199922 46718
rect 200158 46482 200242 46718
rect 200478 46482 200562 46718
rect 200798 46482 200882 46718
rect 201118 46482 201202 46718
rect 201438 46482 201522 46718
rect 201758 46482 201842 46718
rect 202078 46482 202162 46718
rect 202398 46482 202482 46718
rect 202718 46482 202802 46718
rect 203038 46482 203122 46718
rect 203358 46482 203442 46718
rect 203678 46482 203762 46718
rect 203998 46482 204082 46718
rect 204318 46482 204402 46718
rect 204638 46482 204722 46718
rect 204958 46482 207042 46718
rect 207278 46482 207362 46718
rect 207598 46482 207682 46718
rect 207918 46482 208002 46718
rect 208238 46482 208322 46718
rect 208558 46482 208642 46718
rect 208878 46482 208962 46718
rect 209198 46482 209282 46718
rect 209518 46482 209602 46718
rect 209838 46482 209922 46718
rect 210158 46482 210242 46718
rect 210478 46482 210562 46718
rect 210798 46482 210882 46718
rect 211118 46482 211202 46718
rect 211438 46482 211522 46718
rect 211758 46482 211842 46718
rect 212078 46482 212162 46718
rect 212398 46482 212482 46718
rect 212718 46482 212802 46718
rect 213038 46482 213122 46718
rect 213358 46482 213442 46718
rect 213678 46482 213762 46718
rect 213998 46482 214082 46718
rect 214318 46482 214402 46718
rect 214638 46482 214722 46718
rect 214958 46482 217042 46718
rect 217278 46482 217362 46718
rect 217598 46482 217682 46718
rect 217918 46482 218002 46718
rect 218238 46482 218322 46718
rect 218558 46482 218642 46718
rect 218878 46482 218962 46718
rect 219198 46482 219282 46718
rect 219518 46482 219602 46718
rect 219838 46482 219922 46718
rect 220158 46482 220242 46718
rect 220478 46482 220562 46718
rect 220798 46482 220882 46718
rect 221118 46482 221202 46718
rect 221438 46482 221522 46718
rect 221758 46482 221842 46718
rect 222078 46482 222162 46718
rect 222398 46482 222482 46718
rect 222718 46482 222802 46718
rect 223038 46482 223122 46718
rect 223358 46482 223442 46718
rect 223678 46482 223762 46718
rect 223998 46482 224082 46718
rect 224318 46482 224402 46718
rect 224638 46482 224722 46718
rect 224958 46482 227042 46718
rect 227278 46482 227362 46718
rect 227598 46482 227682 46718
rect 227918 46482 228002 46718
rect 228238 46482 228322 46718
rect 228558 46482 228642 46718
rect 228878 46482 228962 46718
rect 229198 46482 229282 46718
rect 229518 46482 229602 46718
rect 229838 46482 229922 46718
rect 230158 46482 230242 46718
rect 230478 46482 230562 46718
rect 230798 46482 230882 46718
rect 231118 46482 231202 46718
rect 231438 46482 231522 46718
rect 231758 46482 231842 46718
rect 232078 46482 232162 46718
rect 232398 46482 232482 46718
rect 232718 46482 232802 46718
rect 233038 46482 233122 46718
rect 233358 46482 233442 46718
rect 233678 46482 233762 46718
rect 233998 46482 234082 46718
rect 234318 46482 234402 46718
rect 234638 46482 234722 46718
rect 234958 46482 237042 46718
rect 237278 46482 237362 46718
rect 237598 46482 237682 46718
rect 237918 46482 238002 46718
rect 238238 46482 238322 46718
rect 238558 46482 238642 46718
rect 238878 46482 238962 46718
rect 239198 46482 239282 46718
rect 239518 46482 239602 46718
rect 239838 46482 239922 46718
rect 240158 46482 240242 46718
rect 240478 46482 240562 46718
rect 240798 46482 240882 46718
rect 241118 46482 241202 46718
rect 241438 46482 241522 46718
rect 241758 46482 241842 46718
rect 242078 46482 242162 46718
rect 242398 46482 242482 46718
rect 242718 46482 242802 46718
rect 243038 46482 243122 46718
rect 243358 46482 243442 46718
rect 243678 46482 243762 46718
rect 243998 46482 244082 46718
rect 244318 46482 244402 46718
rect 244638 46482 244722 46718
rect 244958 46482 247042 46718
rect 247278 46482 247362 46718
rect 247598 46482 247682 46718
rect 247918 46482 248002 46718
rect 248238 46482 248322 46718
rect 248558 46482 248642 46718
rect 248878 46482 248962 46718
rect 249198 46482 249282 46718
rect 249518 46482 249602 46718
rect 249838 46482 249922 46718
rect 250158 46482 250242 46718
rect 250478 46482 250562 46718
rect 250798 46482 250882 46718
rect 251118 46482 251202 46718
rect 251438 46482 251522 46718
rect 251758 46482 251842 46718
rect 252078 46482 252162 46718
rect 252398 46482 252482 46718
rect 252718 46482 252802 46718
rect 253038 46482 253122 46718
rect 253358 46482 253442 46718
rect 253678 46482 253762 46718
rect 253998 46482 254082 46718
rect 254318 46482 254402 46718
rect 254638 46482 254722 46718
rect 254958 46482 257042 46718
rect 257278 46482 257362 46718
rect 257598 46482 257682 46718
rect 257918 46482 258002 46718
rect 258238 46482 258322 46718
rect 258558 46482 258642 46718
rect 258878 46482 258962 46718
rect 259198 46482 259282 46718
rect 259518 46482 259602 46718
rect 259838 46482 259922 46718
rect 260158 46482 260242 46718
rect 260478 46482 260562 46718
rect 260798 46482 260882 46718
rect 261118 46482 261202 46718
rect 261438 46482 261522 46718
rect 261758 46482 261842 46718
rect 262078 46482 262162 46718
rect 262398 46482 262482 46718
rect 262718 46482 262802 46718
rect 263038 46482 263122 46718
rect 263358 46482 263442 46718
rect 263678 46482 263762 46718
rect 263998 46482 264082 46718
rect 264318 46482 264402 46718
rect 264638 46482 264722 46718
rect 264958 46482 267042 46718
rect 267278 46482 267362 46718
rect 267598 46482 267682 46718
rect 267918 46482 268002 46718
rect 268238 46482 268322 46718
rect 268558 46482 268642 46718
rect 268878 46482 268962 46718
rect 269198 46482 269282 46718
rect 269518 46482 269602 46718
rect 269838 46482 269922 46718
rect 270158 46482 270242 46718
rect 270478 46482 270562 46718
rect 270798 46482 270882 46718
rect 271118 46482 271202 46718
rect 271438 46482 271522 46718
rect 271758 46482 271842 46718
rect 272078 46482 272162 46718
rect 272398 46482 272482 46718
rect 272718 46482 272802 46718
rect 273038 46482 273122 46718
rect 273358 46482 273442 46718
rect 273678 46482 273762 46718
rect 273998 46482 274082 46718
rect 274318 46482 274402 46718
rect 274638 46482 274722 46718
rect 274958 46482 277042 46718
rect 277278 46482 277362 46718
rect 277598 46482 277682 46718
rect 277918 46482 278002 46718
rect 278238 46482 278322 46718
rect 278558 46482 278642 46718
rect 278878 46482 278962 46718
rect 279198 46482 279282 46718
rect 279518 46482 279602 46718
rect 279838 46482 279922 46718
rect 280158 46482 280242 46718
rect 280478 46482 280562 46718
rect 280798 46482 280882 46718
rect 281118 46482 281202 46718
rect 281438 46482 281522 46718
rect 281758 46482 281842 46718
rect 282078 46482 282162 46718
rect 282398 46482 282482 46718
rect 282718 46482 282802 46718
rect 283038 46482 283122 46718
rect 283358 46482 283442 46718
rect 283678 46482 283762 46718
rect 283998 46482 284082 46718
rect 284318 46482 284402 46718
rect 284638 46482 284722 46718
rect 284958 46482 286000 46718
rect 46000 46000 286000 46482
rect 46000 45818 54400 46000
rect 43800 26378 45200 26600
rect 43800 25822 44062 26378
rect 44938 25822 45200 26378
rect 46000 26382 46082 45818
rect 54318 26382 54400 45818
rect 46000 26200 54400 26382
rect 56000 45818 64400 46000
rect 56000 26382 56082 45818
rect 64318 26382 64400 45818
rect 56000 26200 64400 26382
rect 66000 45818 74400 46000
rect 66000 26382 66082 45818
rect 74318 26382 74400 45818
rect 66000 26200 74400 26382
rect 76000 45818 84400 46000
rect 76000 26382 76082 45818
rect 84318 26382 84400 45818
rect 76000 26200 84400 26382
rect 86000 45818 94400 46000
rect 86000 26382 86082 45818
rect 94318 26382 94400 45818
rect 86000 26200 94400 26382
rect 96000 45818 104400 46000
rect 96000 26382 96082 45818
rect 104318 26382 104400 45818
rect 96000 26200 104400 26382
rect 106000 45818 114400 46000
rect 106000 26382 106082 45818
rect 114318 26382 114400 45818
rect 106000 26200 114400 26382
rect 116000 45818 124400 46000
rect 116000 26382 116082 45818
rect 124318 26382 124400 45818
rect 116000 26200 124400 26382
rect 126000 45818 134400 46000
rect 126000 26382 126082 45818
rect 134318 26382 134400 45818
rect 126000 26200 134400 26382
rect 136000 45818 144400 46000
rect 136000 26382 136082 45818
rect 144318 26382 144400 45818
rect 136000 26200 144400 26382
rect 146000 45818 154400 46000
rect 146000 26382 146082 45818
rect 154318 26382 154400 45818
rect 146000 26200 154400 26382
rect 156000 45818 164400 46000
rect 156000 26382 156082 45818
rect 164318 26382 164400 45818
rect 156000 26200 164400 26382
rect 166000 45818 174400 46000
rect 166000 26382 166082 45818
rect 174318 26382 174400 45818
rect 166000 26200 174400 26382
rect 176000 45818 184400 46000
rect 176000 26382 176082 45818
rect 184318 26382 184400 45818
rect 176000 26200 184400 26382
rect 186000 45818 194400 46000
rect 186000 26382 186082 45818
rect 194318 26382 194400 45818
rect 186000 26200 194400 26382
rect 196000 45818 204400 46000
rect 196000 26382 196082 45818
rect 204318 26382 204400 45818
rect 196000 26200 204400 26382
rect 206000 45818 214400 46000
rect 206000 26382 206082 45818
rect 214318 26382 214400 45818
rect 206000 26200 214400 26382
rect 216000 45818 224400 46000
rect 216000 26382 216082 45818
rect 224318 26382 224400 45818
rect 216000 26200 224400 26382
rect 226000 45818 234400 46000
rect 226000 26382 226082 45818
rect 234318 26382 234400 45818
rect 226000 26200 234400 26382
rect 236000 45818 244400 46000
rect 236000 26382 236082 45818
rect 244318 26382 244400 45818
rect 236000 26200 244400 26382
rect 246000 45818 254400 46000
rect 246000 26382 246082 45818
rect 254318 26382 254400 45818
rect 246000 26200 254400 26382
rect 256000 45818 264400 46000
rect 256000 26382 256082 45818
rect 264318 26382 264400 45818
rect 256000 26200 264400 26382
rect 266000 45818 274400 46000
rect 266000 26382 266082 45818
rect 274318 26382 274400 45818
rect 266000 26200 274400 26382
rect 276000 45818 284400 46000
rect 276000 26382 276082 45818
rect 284318 26382 284400 45818
rect 276000 26200 284400 26382
rect 43800 25600 45200 25822
rect 47600 25800 54400 26200
rect 57600 25800 64400 26200
rect 67600 25800 74400 26200
rect 77600 25800 84400 26200
rect 87600 25800 94400 26200
rect 97600 25800 104400 26200
rect 107600 25800 114400 26200
rect 117600 25800 124400 26200
rect 127600 25800 134400 26200
rect 137600 25800 144400 26200
rect 147600 25800 154400 26200
rect 157600 25800 164400 26200
rect 167600 25800 174400 26200
rect 177600 25800 184400 26200
rect 187600 25800 194400 26200
rect 197600 25800 204400 26200
rect 207600 25800 214400 26200
rect 217600 25800 224400 26200
rect 227600 25800 234400 26200
rect 237600 25800 244400 26200
rect 247600 25800 254400 26200
rect 257600 25800 264400 26200
rect 267600 25800 274400 26200
rect 277600 25800 284400 26200
rect 47600 25618 56000 25800
rect 43800 6178 45200 6400
rect 43800 5622 44062 6178
rect 44938 5622 45200 6178
rect 47600 6182 47682 25618
rect 55918 6182 56000 25618
rect 47600 6000 56000 6182
rect 57600 25618 66000 25800
rect 57600 6182 57682 25618
rect 65918 6182 66000 25618
rect 57600 6000 66000 6182
rect 67600 25618 76000 25800
rect 67600 6182 67682 25618
rect 75918 6182 76000 25618
rect 67600 6000 76000 6182
rect 77600 25618 86000 25800
rect 77600 6182 77682 25618
rect 85918 6182 86000 25618
rect 77600 6000 86000 6182
rect 87600 25618 96000 25800
rect 87600 6182 87682 25618
rect 95918 6182 96000 25618
rect 87600 6000 96000 6182
rect 97600 25618 106000 25800
rect 97600 6182 97682 25618
rect 105918 6182 106000 25618
rect 97600 6000 106000 6182
rect 107600 25618 116000 25800
rect 107600 6182 107682 25618
rect 115918 6182 116000 25618
rect 107600 6000 116000 6182
rect 117600 25618 126000 25800
rect 117600 6182 117682 25618
rect 125918 6182 126000 25618
rect 117600 6000 126000 6182
rect 127600 25618 136000 25800
rect 127600 6182 127682 25618
rect 135918 6182 136000 25618
rect 127600 6000 136000 6182
rect 137600 25618 146000 25800
rect 137600 6182 137682 25618
rect 145918 6182 146000 25618
rect 137600 6000 146000 6182
rect 147600 25618 156000 25800
rect 147600 6182 147682 25618
rect 155918 6182 156000 25618
rect 147600 6000 156000 6182
rect 157600 25618 166000 25800
rect 157600 6182 157682 25618
rect 165918 6182 166000 25618
rect 157600 6000 166000 6182
rect 167600 25618 176000 25800
rect 167600 6182 167682 25618
rect 175918 6182 176000 25618
rect 167600 6000 176000 6182
rect 177600 25618 186000 25800
rect 177600 6182 177682 25618
rect 185918 6182 186000 25618
rect 177600 6000 186000 6182
rect 187600 25618 196000 25800
rect 187600 6182 187682 25618
rect 195918 6182 196000 25618
rect 187600 6000 196000 6182
rect 197600 25618 206000 25800
rect 197600 6182 197682 25618
rect 205918 6182 206000 25618
rect 197600 6000 206000 6182
rect 207600 25618 216000 25800
rect 207600 6182 207682 25618
rect 215918 6182 216000 25618
rect 207600 6000 216000 6182
rect 217600 25618 226000 25800
rect 217600 6182 217682 25618
rect 225918 6182 226000 25618
rect 217600 6000 226000 6182
rect 227600 25618 236000 25800
rect 227600 6182 227682 25618
rect 235918 6182 236000 25618
rect 227600 6000 236000 6182
rect 237600 25618 246000 25800
rect 237600 6182 237682 25618
rect 245918 6182 246000 25618
rect 237600 6000 246000 6182
rect 247600 25618 256000 25800
rect 247600 6182 247682 25618
rect 255918 6182 256000 25618
rect 247600 6000 256000 6182
rect 257600 25618 266000 25800
rect 257600 6182 257682 25618
rect 265918 6182 266000 25618
rect 257600 6000 266000 6182
rect 267600 25618 276000 25800
rect 267600 6182 267682 25618
rect 275918 6182 276000 25618
rect 267600 6000 276000 6182
rect 277600 25618 286000 25800
rect 277600 6182 277682 25618
rect 285918 6182 286000 25618
rect 277600 6000 286000 6182
rect 43800 5400 45200 5622
rect 46000 5518 286000 6000
rect 46000 5282 47042 5518
rect 47278 5282 47362 5518
rect 47598 5282 47682 5518
rect 47918 5282 48002 5518
rect 48238 5282 48322 5518
rect 48558 5282 48642 5518
rect 48878 5282 48962 5518
rect 49198 5282 49282 5518
rect 49518 5282 49602 5518
rect 49838 5282 49922 5518
rect 50158 5282 50242 5518
rect 50478 5282 50562 5518
rect 50798 5282 50882 5518
rect 51118 5282 51202 5518
rect 51438 5282 51522 5518
rect 51758 5282 51842 5518
rect 52078 5282 52162 5518
rect 52398 5282 52482 5518
rect 52718 5282 52802 5518
rect 53038 5282 53122 5518
rect 53358 5282 53442 5518
rect 53678 5282 53762 5518
rect 53998 5282 54082 5518
rect 54318 5282 54402 5518
rect 54638 5282 54722 5518
rect 54958 5282 57042 5518
rect 57278 5282 57362 5518
rect 57598 5282 57682 5518
rect 57918 5282 58002 5518
rect 58238 5282 58322 5518
rect 58558 5282 58642 5518
rect 58878 5282 58962 5518
rect 59198 5282 59282 5518
rect 59518 5282 59602 5518
rect 59838 5282 59922 5518
rect 60158 5282 60242 5518
rect 60478 5282 60562 5518
rect 60798 5282 60882 5518
rect 61118 5282 61202 5518
rect 61438 5282 61522 5518
rect 61758 5282 61842 5518
rect 62078 5282 62162 5518
rect 62398 5282 62482 5518
rect 62718 5282 62802 5518
rect 63038 5282 63122 5518
rect 63358 5282 63442 5518
rect 63678 5282 63762 5518
rect 63998 5282 64082 5518
rect 64318 5282 64402 5518
rect 64638 5282 64722 5518
rect 64958 5282 67042 5518
rect 67278 5282 67362 5518
rect 67598 5282 67682 5518
rect 67918 5282 68002 5518
rect 68238 5282 68322 5518
rect 68558 5282 68642 5518
rect 68878 5282 68962 5518
rect 69198 5282 69282 5518
rect 69518 5282 69602 5518
rect 69838 5282 69922 5518
rect 70158 5282 70242 5518
rect 70478 5282 70562 5518
rect 70798 5282 70882 5518
rect 71118 5282 71202 5518
rect 71438 5282 71522 5518
rect 71758 5282 71842 5518
rect 72078 5282 72162 5518
rect 72398 5282 72482 5518
rect 72718 5282 72802 5518
rect 73038 5282 73122 5518
rect 73358 5282 73442 5518
rect 73678 5282 73762 5518
rect 73998 5282 74082 5518
rect 74318 5282 74402 5518
rect 74638 5282 74722 5518
rect 74958 5282 77042 5518
rect 77278 5282 77362 5518
rect 77598 5282 77682 5518
rect 77918 5282 78002 5518
rect 78238 5282 78322 5518
rect 78558 5282 78642 5518
rect 78878 5282 78962 5518
rect 79198 5282 79282 5518
rect 79518 5282 79602 5518
rect 79838 5282 79922 5518
rect 80158 5282 80242 5518
rect 80478 5282 80562 5518
rect 80798 5282 80882 5518
rect 81118 5282 81202 5518
rect 81438 5282 81522 5518
rect 81758 5282 81842 5518
rect 82078 5282 82162 5518
rect 82398 5282 82482 5518
rect 82718 5282 82802 5518
rect 83038 5282 83122 5518
rect 83358 5282 83442 5518
rect 83678 5282 83762 5518
rect 83998 5282 84082 5518
rect 84318 5282 84402 5518
rect 84638 5282 84722 5518
rect 84958 5282 87042 5518
rect 87278 5282 87362 5518
rect 87598 5282 87682 5518
rect 87918 5282 88002 5518
rect 88238 5282 88322 5518
rect 88558 5282 88642 5518
rect 88878 5282 88962 5518
rect 89198 5282 89282 5518
rect 89518 5282 89602 5518
rect 89838 5282 89922 5518
rect 90158 5282 90242 5518
rect 90478 5282 90562 5518
rect 90798 5282 90882 5518
rect 91118 5282 91202 5518
rect 91438 5282 91522 5518
rect 91758 5282 91842 5518
rect 92078 5282 92162 5518
rect 92398 5282 92482 5518
rect 92718 5282 92802 5518
rect 93038 5282 93122 5518
rect 93358 5282 93442 5518
rect 93678 5282 93762 5518
rect 93998 5282 94082 5518
rect 94318 5282 94402 5518
rect 94638 5282 94722 5518
rect 94958 5282 97042 5518
rect 97278 5282 97362 5518
rect 97598 5282 97682 5518
rect 97918 5282 98002 5518
rect 98238 5282 98322 5518
rect 98558 5282 98642 5518
rect 98878 5282 98962 5518
rect 99198 5282 99282 5518
rect 99518 5282 99602 5518
rect 99838 5282 99922 5518
rect 100158 5282 100242 5518
rect 100478 5282 100562 5518
rect 100798 5282 100882 5518
rect 101118 5282 101202 5518
rect 101438 5282 101522 5518
rect 101758 5282 101842 5518
rect 102078 5282 102162 5518
rect 102398 5282 102482 5518
rect 102718 5282 102802 5518
rect 103038 5282 103122 5518
rect 103358 5282 103442 5518
rect 103678 5282 103762 5518
rect 103998 5282 104082 5518
rect 104318 5282 104402 5518
rect 104638 5282 104722 5518
rect 104958 5282 107042 5518
rect 107278 5282 107362 5518
rect 107598 5282 107682 5518
rect 107918 5282 108002 5518
rect 108238 5282 108322 5518
rect 108558 5282 108642 5518
rect 108878 5282 108962 5518
rect 109198 5282 109282 5518
rect 109518 5282 109602 5518
rect 109838 5282 109922 5518
rect 110158 5282 110242 5518
rect 110478 5282 110562 5518
rect 110798 5282 110882 5518
rect 111118 5282 111202 5518
rect 111438 5282 111522 5518
rect 111758 5282 111842 5518
rect 112078 5282 112162 5518
rect 112398 5282 112482 5518
rect 112718 5282 112802 5518
rect 113038 5282 113122 5518
rect 113358 5282 113442 5518
rect 113678 5282 113762 5518
rect 113998 5282 114082 5518
rect 114318 5282 114402 5518
rect 114638 5282 114722 5518
rect 114958 5282 117042 5518
rect 117278 5282 117362 5518
rect 117598 5282 117682 5518
rect 117918 5282 118002 5518
rect 118238 5282 118322 5518
rect 118558 5282 118642 5518
rect 118878 5282 118962 5518
rect 119198 5282 119282 5518
rect 119518 5282 119602 5518
rect 119838 5282 119922 5518
rect 120158 5282 120242 5518
rect 120478 5282 120562 5518
rect 120798 5282 120882 5518
rect 121118 5282 121202 5518
rect 121438 5282 121522 5518
rect 121758 5282 121842 5518
rect 122078 5282 122162 5518
rect 122398 5282 122482 5518
rect 122718 5282 122802 5518
rect 123038 5282 123122 5518
rect 123358 5282 123442 5518
rect 123678 5282 123762 5518
rect 123998 5282 124082 5518
rect 124318 5282 124402 5518
rect 124638 5282 124722 5518
rect 124958 5282 127042 5518
rect 127278 5282 127362 5518
rect 127598 5282 127682 5518
rect 127918 5282 128002 5518
rect 128238 5282 128322 5518
rect 128558 5282 128642 5518
rect 128878 5282 128962 5518
rect 129198 5282 129282 5518
rect 129518 5282 129602 5518
rect 129838 5282 129922 5518
rect 130158 5282 130242 5518
rect 130478 5282 130562 5518
rect 130798 5282 130882 5518
rect 131118 5282 131202 5518
rect 131438 5282 131522 5518
rect 131758 5282 131842 5518
rect 132078 5282 132162 5518
rect 132398 5282 132482 5518
rect 132718 5282 132802 5518
rect 133038 5282 133122 5518
rect 133358 5282 133442 5518
rect 133678 5282 133762 5518
rect 133998 5282 134082 5518
rect 134318 5282 134402 5518
rect 134638 5282 134722 5518
rect 134958 5282 137042 5518
rect 137278 5282 137362 5518
rect 137598 5282 137682 5518
rect 137918 5282 138002 5518
rect 138238 5282 138322 5518
rect 138558 5282 138642 5518
rect 138878 5282 138962 5518
rect 139198 5282 139282 5518
rect 139518 5282 139602 5518
rect 139838 5282 139922 5518
rect 140158 5282 140242 5518
rect 140478 5282 140562 5518
rect 140798 5282 140882 5518
rect 141118 5282 141202 5518
rect 141438 5282 141522 5518
rect 141758 5282 141842 5518
rect 142078 5282 142162 5518
rect 142398 5282 142482 5518
rect 142718 5282 142802 5518
rect 143038 5282 143122 5518
rect 143358 5282 143442 5518
rect 143678 5282 143762 5518
rect 143998 5282 144082 5518
rect 144318 5282 144402 5518
rect 144638 5282 144722 5518
rect 144958 5282 147042 5518
rect 147278 5282 147362 5518
rect 147598 5282 147682 5518
rect 147918 5282 148002 5518
rect 148238 5282 148322 5518
rect 148558 5282 148642 5518
rect 148878 5282 148962 5518
rect 149198 5282 149282 5518
rect 149518 5282 149602 5518
rect 149838 5282 149922 5518
rect 150158 5282 150242 5518
rect 150478 5282 150562 5518
rect 150798 5282 150882 5518
rect 151118 5282 151202 5518
rect 151438 5282 151522 5518
rect 151758 5282 151842 5518
rect 152078 5282 152162 5518
rect 152398 5282 152482 5518
rect 152718 5282 152802 5518
rect 153038 5282 153122 5518
rect 153358 5282 153442 5518
rect 153678 5282 153762 5518
rect 153998 5282 154082 5518
rect 154318 5282 154402 5518
rect 154638 5282 154722 5518
rect 154958 5282 157042 5518
rect 157278 5282 157362 5518
rect 157598 5282 157682 5518
rect 157918 5282 158002 5518
rect 158238 5282 158322 5518
rect 158558 5282 158642 5518
rect 158878 5282 158962 5518
rect 159198 5282 159282 5518
rect 159518 5282 159602 5518
rect 159838 5282 159922 5518
rect 160158 5282 160242 5518
rect 160478 5282 160562 5518
rect 160798 5282 160882 5518
rect 161118 5282 161202 5518
rect 161438 5282 161522 5518
rect 161758 5282 161842 5518
rect 162078 5282 162162 5518
rect 162398 5282 162482 5518
rect 162718 5282 162802 5518
rect 163038 5282 163122 5518
rect 163358 5282 163442 5518
rect 163678 5282 163762 5518
rect 163998 5282 164082 5518
rect 164318 5282 164402 5518
rect 164638 5282 164722 5518
rect 164958 5282 167042 5518
rect 167278 5282 167362 5518
rect 167598 5282 167682 5518
rect 167918 5282 168002 5518
rect 168238 5282 168322 5518
rect 168558 5282 168642 5518
rect 168878 5282 168962 5518
rect 169198 5282 169282 5518
rect 169518 5282 169602 5518
rect 169838 5282 169922 5518
rect 170158 5282 170242 5518
rect 170478 5282 170562 5518
rect 170798 5282 170882 5518
rect 171118 5282 171202 5518
rect 171438 5282 171522 5518
rect 171758 5282 171842 5518
rect 172078 5282 172162 5518
rect 172398 5282 172482 5518
rect 172718 5282 172802 5518
rect 173038 5282 173122 5518
rect 173358 5282 173442 5518
rect 173678 5282 173762 5518
rect 173998 5282 174082 5518
rect 174318 5282 174402 5518
rect 174638 5282 174722 5518
rect 174958 5282 177042 5518
rect 177278 5282 177362 5518
rect 177598 5282 177682 5518
rect 177918 5282 178002 5518
rect 178238 5282 178322 5518
rect 178558 5282 178642 5518
rect 178878 5282 178962 5518
rect 179198 5282 179282 5518
rect 179518 5282 179602 5518
rect 179838 5282 179922 5518
rect 180158 5282 180242 5518
rect 180478 5282 180562 5518
rect 180798 5282 180882 5518
rect 181118 5282 181202 5518
rect 181438 5282 181522 5518
rect 181758 5282 181842 5518
rect 182078 5282 182162 5518
rect 182398 5282 182482 5518
rect 182718 5282 182802 5518
rect 183038 5282 183122 5518
rect 183358 5282 183442 5518
rect 183678 5282 183762 5518
rect 183998 5282 184082 5518
rect 184318 5282 184402 5518
rect 184638 5282 184722 5518
rect 184958 5282 187042 5518
rect 187278 5282 187362 5518
rect 187598 5282 187682 5518
rect 187918 5282 188002 5518
rect 188238 5282 188322 5518
rect 188558 5282 188642 5518
rect 188878 5282 188962 5518
rect 189198 5282 189282 5518
rect 189518 5282 189602 5518
rect 189838 5282 189922 5518
rect 190158 5282 190242 5518
rect 190478 5282 190562 5518
rect 190798 5282 190882 5518
rect 191118 5282 191202 5518
rect 191438 5282 191522 5518
rect 191758 5282 191842 5518
rect 192078 5282 192162 5518
rect 192398 5282 192482 5518
rect 192718 5282 192802 5518
rect 193038 5282 193122 5518
rect 193358 5282 193442 5518
rect 193678 5282 193762 5518
rect 193998 5282 194082 5518
rect 194318 5282 194402 5518
rect 194638 5282 194722 5518
rect 194958 5282 197042 5518
rect 197278 5282 197362 5518
rect 197598 5282 197682 5518
rect 197918 5282 198002 5518
rect 198238 5282 198322 5518
rect 198558 5282 198642 5518
rect 198878 5282 198962 5518
rect 199198 5282 199282 5518
rect 199518 5282 199602 5518
rect 199838 5282 199922 5518
rect 200158 5282 200242 5518
rect 200478 5282 200562 5518
rect 200798 5282 200882 5518
rect 201118 5282 201202 5518
rect 201438 5282 201522 5518
rect 201758 5282 201842 5518
rect 202078 5282 202162 5518
rect 202398 5282 202482 5518
rect 202718 5282 202802 5518
rect 203038 5282 203122 5518
rect 203358 5282 203442 5518
rect 203678 5282 203762 5518
rect 203998 5282 204082 5518
rect 204318 5282 204402 5518
rect 204638 5282 204722 5518
rect 204958 5282 207042 5518
rect 207278 5282 207362 5518
rect 207598 5282 207682 5518
rect 207918 5282 208002 5518
rect 208238 5282 208322 5518
rect 208558 5282 208642 5518
rect 208878 5282 208962 5518
rect 209198 5282 209282 5518
rect 209518 5282 209602 5518
rect 209838 5282 209922 5518
rect 210158 5282 210242 5518
rect 210478 5282 210562 5518
rect 210798 5282 210882 5518
rect 211118 5282 211202 5518
rect 211438 5282 211522 5518
rect 211758 5282 211842 5518
rect 212078 5282 212162 5518
rect 212398 5282 212482 5518
rect 212718 5282 212802 5518
rect 213038 5282 213122 5518
rect 213358 5282 213442 5518
rect 213678 5282 213762 5518
rect 213998 5282 214082 5518
rect 214318 5282 214402 5518
rect 214638 5282 214722 5518
rect 214958 5282 217042 5518
rect 217278 5282 217362 5518
rect 217598 5282 217682 5518
rect 217918 5282 218002 5518
rect 218238 5282 218322 5518
rect 218558 5282 218642 5518
rect 218878 5282 218962 5518
rect 219198 5282 219282 5518
rect 219518 5282 219602 5518
rect 219838 5282 219922 5518
rect 220158 5282 220242 5518
rect 220478 5282 220562 5518
rect 220798 5282 220882 5518
rect 221118 5282 221202 5518
rect 221438 5282 221522 5518
rect 221758 5282 221842 5518
rect 222078 5282 222162 5518
rect 222398 5282 222482 5518
rect 222718 5282 222802 5518
rect 223038 5282 223122 5518
rect 223358 5282 223442 5518
rect 223678 5282 223762 5518
rect 223998 5282 224082 5518
rect 224318 5282 224402 5518
rect 224638 5282 224722 5518
rect 224958 5282 227042 5518
rect 227278 5282 227362 5518
rect 227598 5282 227682 5518
rect 227918 5282 228002 5518
rect 228238 5282 228322 5518
rect 228558 5282 228642 5518
rect 228878 5282 228962 5518
rect 229198 5282 229282 5518
rect 229518 5282 229602 5518
rect 229838 5282 229922 5518
rect 230158 5282 230242 5518
rect 230478 5282 230562 5518
rect 230798 5282 230882 5518
rect 231118 5282 231202 5518
rect 231438 5282 231522 5518
rect 231758 5282 231842 5518
rect 232078 5282 232162 5518
rect 232398 5282 232482 5518
rect 232718 5282 232802 5518
rect 233038 5282 233122 5518
rect 233358 5282 233442 5518
rect 233678 5282 233762 5518
rect 233998 5282 234082 5518
rect 234318 5282 234402 5518
rect 234638 5282 234722 5518
rect 234958 5282 237042 5518
rect 237278 5282 237362 5518
rect 237598 5282 237682 5518
rect 237918 5282 238002 5518
rect 238238 5282 238322 5518
rect 238558 5282 238642 5518
rect 238878 5282 238962 5518
rect 239198 5282 239282 5518
rect 239518 5282 239602 5518
rect 239838 5282 239922 5518
rect 240158 5282 240242 5518
rect 240478 5282 240562 5518
rect 240798 5282 240882 5518
rect 241118 5282 241202 5518
rect 241438 5282 241522 5518
rect 241758 5282 241842 5518
rect 242078 5282 242162 5518
rect 242398 5282 242482 5518
rect 242718 5282 242802 5518
rect 243038 5282 243122 5518
rect 243358 5282 243442 5518
rect 243678 5282 243762 5518
rect 243998 5282 244082 5518
rect 244318 5282 244402 5518
rect 244638 5282 244722 5518
rect 244958 5282 247042 5518
rect 247278 5282 247362 5518
rect 247598 5282 247682 5518
rect 247918 5282 248002 5518
rect 248238 5282 248322 5518
rect 248558 5282 248642 5518
rect 248878 5282 248962 5518
rect 249198 5282 249282 5518
rect 249518 5282 249602 5518
rect 249838 5282 249922 5518
rect 250158 5282 250242 5518
rect 250478 5282 250562 5518
rect 250798 5282 250882 5518
rect 251118 5282 251202 5518
rect 251438 5282 251522 5518
rect 251758 5282 251842 5518
rect 252078 5282 252162 5518
rect 252398 5282 252482 5518
rect 252718 5282 252802 5518
rect 253038 5282 253122 5518
rect 253358 5282 253442 5518
rect 253678 5282 253762 5518
rect 253998 5282 254082 5518
rect 254318 5282 254402 5518
rect 254638 5282 254722 5518
rect 254958 5282 257042 5518
rect 257278 5282 257362 5518
rect 257598 5282 257682 5518
rect 257918 5282 258002 5518
rect 258238 5282 258322 5518
rect 258558 5282 258642 5518
rect 258878 5282 258962 5518
rect 259198 5282 259282 5518
rect 259518 5282 259602 5518
rect 259838 5282 259922 5518
rect 260158 5282 260242 5518
rect 260478 5282 260562 5518
rect 260798 5282 260882 5518
rect 261118 5282 261202 5518
rect 261438 5282 261522 5518
rect 261758 5282 261842 5518
rect 262078 5282 262162 5518
rect 262398 5282 262482 5518
rect 262718 5282 262802 5518
rect 263038 5282 263122 5518
rect 263358 5282 263442 5518
rect 263678 5282 263762 5518
rect 263998 5282 264082 5518
rect 264318 5282 264402 5518
rect 264638 5282 264722 5518
rect 264958 5282 267042 5518
rect 267278 5282 267362 5518
rect 267598 5282 267682 5518
rect 267918 5282 268002 5518
rect 268238 5282 268322 5518
rect 268558 5282 268642 5518
rect 268878 5282 268962 5518
rect 269198 5282 269282 5518
rect 269518 5282 269602 5518
rect 269838 5282 269922 5518
rect 270158 5282 270242 5518
rect 270478 5282 270562 5518
rect 270798 5282 270882 5518
rect 271118 5282 271202 5518
rect 271438 5282 271522 5518
rect 271758 5282 271842 5518
rect 272078 5282 272162 5518
rect 272398 5282 272482 5518
rect 272718 5282 272802 5518
rect 273038 5282 273122 5518
rect 273358 5282 273442 5518
rect 273678 5282 273762 5518
rect 273998 5282 274082 5518
rect 274318 5282 274402 5518
rect 274638 5282 274722 5518
rect 274958 5282 277042 5518
rect 277278 5282 277362 5518
rect 277598 5282 277682 5518
rect 277918 5282 278002 5518
rect 278238 5282 278322 5518
rect 278558 5282 278642 5518
rect 278878 5282 278962 5518
rect 279198 5282 279282 5518
rect 279518 5282 279602 5518
rect 279838 5282 279922 5518
rect 280158 5282 280242 5518
rect 280478 5282 280562 5518
rect 280798 5282 280882 5518
rect 281118 5282 281202 5518
rect 281438 5282 281522 5518
rect 281758 5282 281842 5518
rect 282078 5282 282162 5518
rect 282398 5282 282482 5518
rect 282718 5282 282802 5518
rect 283038 5282 283122 5518
rect 283358 5282 283442 5518
rect 283678 5282 283762 5518
rect 283998 5282 284082 5518
rect 284318 5282 284402 5518
rect 284638 5282 284722 5518
rect 284958 5282 286000 5518
rect 46000 5200 286000 5282
use sky130_fd_pr__res_xhigh_po_0p35_FE9J4G  sky130_fd_pr__res_xhigh_po_0p35_FE9J4G_0
timestamp 1672341375
transform -1 0 45401 0 -1 15998
box -191 -10588 191 10588
<< labels >>
rlabel metal5 s 43800 25600 43990 26600 4 A
port 1 se
rlabel metal5 s 43800 5400 43990 6400 4 B
port 3 se
rlabel metal4 s 45040 15750 45160 16750 4 VLO
port 2 se
<< end >>
