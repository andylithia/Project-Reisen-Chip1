magic
tech sky130A
magscale 1 2
timestamp 1672030875
<< metal3 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46000 286000 46240
rect 46000 26200 54400 46000
rect 56000 26200 64400 46000
rect 66000 26200 74400 46000
rect 76000 26200 84400 46000
rect 86000 26200 94400 46000
rect 96000 26200 104400 46000
rect 106000 26200 114400 46000
rect 116000 26200 124400 46000
rect 126000 26200 134400 46000
rect 136000 26200 144400 46000
rect 146000 26200 154400 46000
rect 156000 26200 164400 46000
rect 166000 26200 174400 46000
rect 176000 26200 184400 46000
rect 186000 26200 194400 46000
rect 196000 26200 204400 46000
rect 206000 26200 214400 46000
rect 216000 26200 224400 46000
rect 226000 26200 234400 46000
rect 236000 26200 244400 46000
rect 246000 26200 254400 46000
rect 256000 26200 264400 46000
rect 266000 26200 274400 46000
rect 276000 26200 284400 46000
rect 47600 25800 54400 26200
rect 57600 25800 64400 26200
rect 67600 25800 74400 26200
rect 77600 25800 84400 26200
rect 87600 25800 94400 26200
rect 97600 25800 104400 26200
rect 107600 25800 114400 26200
rect 117600 25800 124400 26200
rect 127600 25800 134400 26200
rect 137600 25800 144400 26200
rect 147600 25800 154400 26200
rect 157600 25800 164400 26200
rect 167600 25800 174400 26200
rect 177600 25800 184400 26200
rect 187600 25800 194400 26200
rect 197600 25800 204400 26200
rect 207600 25800 214400 26200
rect 217600 25800 224400 26200
rect 227600 25800 234400 26200
rect 237600 25800 244400 26200
rect 247600 25800 254400 26200
rect 257600 25800 264400 26200
rect 267600 25800 274400 26200
rect 277600 25800 284400 26200
rect 47600 6000 56000 25800
rect 57600 6000 66000 25800
rect 67600 6000 76000 25800
rect 77600 6000 86000 25800
rect 87600 6000 96000 25800
rect 97600 6000 106000 25800
rect 107600 6000 116000 25800
rect 117600 6000 126000 25800
rect 127600 6000 136000 25800
rect 137600 6000 146000 25800
rect 147600 6000 156000 25800
rect 157600 6000 166000 25800
rect 167600 6000 176000 25800
rect 177600 6000 186000 25800
rect 187600 6000 196000 25800
rect 197600 6000 206000 25800
rect 207600 6000 216000 25800
rect 217600 6000 226000 25800
rect 227600 6000 236000 25800
rect 237600 6000 246000 25800
rect 247600 6000 256000 25800
rect 257600 6000 266000 25800
rect 267600 6000 276000 25800
rect 277600 6000 286000 25800
rect 46000 5760 286000 6000
rect 46000 5440 47000 5760
rect 55960 5440 57000 5760
rect 65960 5440 67000 5760
rect 75960 5440 77000 5760
rect 85960 5440 87000 5760
rect 95960 5440 97000 5760
rect 105960 5440 107000 5760
rect 115960 5440 117000 5760
rect 125960 5440 127000 5760
rect 135960 5440 137000 5760
rect 145960 5440 147000 5760
rect 155960 5440 157000 5760
rect 165960 5440 167000 5760
rect 175960 5440 177000 5760
rect 185960 5440 187000 5760
rect 195960 5440 197000 5760
rect 205960 5440 207000 5760
rect 215960 5440 217000 5760
rect 225960 5440 227000 5760
rect 235960 5440 237000 5760
rect 245960 5440 247000 5760
rect 255960 5440 257000 5760
rect 265960 5440 267000 5760
rect 275960 5440 277000 5760
rect 285960 5440 286000 5760
rect 46000 5400 286000 5440
<< via3 >>
rect 47000 46240 55000 46560
rect 57000 46240 65000 46560
rect 67000 46240 75000 46560
rect 77000 46240 85000 46560
rect 87000 46240 95000 46560
rect 97000 46240 105000 46560
rect 107000 46240 115000 46560
rect 117000 46240 125000 46560
rect 127000 46240 135000 46560
rect 137000 46240 145000 46560
rect 147000 46240 155000 46560
rect 157000 46240 165000 46560
rect 167000 46240 175000 46560
rect 177000 46240 185000 46560
rect 187000 46240 195000 46560
rect 197000 46240 205000 46560
rect 207000 46240 215000 46560
rect 217000 46240 225000 46560
rect 227000 46240 235000 46560
rect 237000 46240 245000 46560
rect 247000 46240 255000 46560
rect 257000 46240 265000 46560
rect 267000 46240 275000 46560
rect 277000 46240 285000 46560
rect 47000 5440 55960 5760
rect 57000 5440 65960 5760
rect 67000 5440 75960 5760
rect 77000 5440 85960 5760
rect 87000 5440 95960 5760
rect 97000 5440 105960 5760
rect 107000 5440 115960 5760
rect 117000 5440 125960 5760
rect 127000 5440 135960 5760
rect 137000 5440 145960 5760
rect 147000 5440 155960 5760
rect 157000 5440 165960 5760
rect 167000 5440 175960 5760
rect 177000 5440 185960 5760
rect 187000 5440 195960 5760
rect 197000 5440 205960 5760
rect 207000 5440 215960 5760
rect 217000 5440 225960 5760
rect 227000 5440 235960 5760
rect 237000 5440 245960 5760
rect 247000 5440 255960 5760
rect 257000 5440 265960 5760
rect 267000 5440 275960 5760
rect 277000 5440 285960 5760
<< mimcap >>
rect 46040 45940 54360 45960
rect 46040 26260 46060 45940
rect 54340 26260 54360 45940
rect 46040 26240 54360 26260
rect 56040 45940 64360 45960
rect 56040 26260 56060 45940
rect 64340 26260 64360 45940
rect 56040 26240 64360 26260
rect 66040 45940 74360 45960
rect 66040 26260 66060 45940
rect 74340 26260 74360 45940
rect 66040 26240 74360 26260
rect 76040 45940 84360 45960
rect 76040 26260 76060 45940
rect 84340 26260 84360 45940
rect 76040 26240 84360 26260
rect 86040 45940 94360 45960
rect 86040 26260 86060 45940
rect 94340 26260 94360 45940
rect 86040 26240 94360 26260
rect 96040 45940 104360 45960
rect 96040 26260 96060 45940
rect 104340 26260 104360 45940
rect 96040 26240 104360 26260
rect 106040 45940 114360 45960
rect 106040 26260 106060 45940
rect 114340 26260 114360 45940
rect 106040 26240 114360 26260
rect 116040 45940 124360 45960
rect 116040 26260 116060 45940
rect 124340 26260 124360 45940
rect 116040 26240 124360 26260
rect 126040 45940 134360 45960
rect 126040 26260 126060 45940
rect 134340 26260 134360 45940
rect 126040 26240 134360 26260
rect 136040 45940 144360 45960
rect 136040 26260 136060 45940
rect 144340 26260 144360 45940
rect 136040 26240 144360 26260
rect 146040 45940 154360 45960
rect 146040 26260 146060 45940
rect 154340 26260 154360 45940
rect 146040 26240 154360 26260
rect 156040 45940 164360 45960
rect 156040 26260 156060 45940
rect 164340 26260 164360 45940
rect 156040 26240 164360 26260
rect 166040 45940 174360 45960
rect 166040 26260 166060 45940
rect 174340 26260 174360 45940
rect 166040 26240 174360 26260
rect 176040 45940 184360 45960
rect 176040 26260 176060 45940
rect 184340 26260 184360 45940
rect 176040 26240 184360 26260
rect 186040 45940 194360 45960
rect 186040 26260 186060 45940
rect 194340 26260 194360 45940
rect 186040 26240 194360 26260
rect 196040 45940 204360 45960
rect 196040 26260 196060 45940
rect 204340 26260 204360 45940
rect 196040 26240 204360 26260
rect 206040 45940 214360 45960
rect 206040 26260 206060 45940
rect 214340 26260 214360 45940
rect 206040 26240 214360 26260
rect 216040 45940 224360 45960
rect 216040 26260 216060 45940
rect 224340 26260 224360 45940
rect 216040 26240 224360 26260
rect 226040 45940 234360 45960
rect 226040 26260 226060 45940
rect 234340 26260 234360 45940
rect 226040 26240 234360 26260
rect 236040 45940 244360 45960
rect 236040 26260 236060 45940
rect 244340 26260 244360 45940
rect 236040 26240 244360 26260
rect 246040 45940 254360 45960
rect 246040 26260 246060 45940
rect 254340 26260 254360 45940
rect 246040 26240 254360 26260
rect 256040 45940 264360 45960
rect 256040 26260 256060 45940
rect 264340 26260 264360 45940
rect 256040 26240 264360 26260
rect 266040 45940 274360 45960
rect 266040 26260 266060 45940
rect 274340 26260 274360 45940
rect 266040 26240 274360 26260
rect 276040 45940 284360 45960
rect 276040 26260 276060 45940
rect 284340 26260 284360 45940
rect 276040 26240 284360 26260
rect 47640 25740 55960 25760
rect 47640 6060 47660 25740
rect 55940 6060 55960 25740
rect 47640 6040 55960 6060
rect 57640 25740 65960 25760
rect 57640 6060 57660 25740
rect 65940 6060 65960 25740
rect 57640 6040 65960 6060
rect 67640 25740 75960 25760
rect 67640 6060 67660 25740
rect 75940 6060 75960 25740
rect 67640 6040 75960 6060
rect 77640 25740 85960 25760
rect 77640 6060 77660 25740
rect 85940 6060 85960 25740
rect 77640 6040 85960 6060
rect 87640 25740 95960 25760
rect 87640 6060 87660 25740
rect 95940 6060 95960 25740
rect 87640 6040 95960 6060
rect 97640 25740 105960 25760
rect 97640 6060 97660 25740
rect 105940 6060 105960 25740
rect 97640 6040 105960 6060
rect 107640 25740 115960 25760
rect 107640 6060 107660 25740
rect 115940 6060 115960 25740
rect 107640 6040 115960 6060
rect 117640 25740 125960 25760
rect 117640 6060 117660 25740
rect 125940 6060 125960 25740
rect 117640 6040 125960 6060
rect 127640 25740 135960 25760
rect 127640 6060 127660 25740
rect 135940 6060 135960 25740
rect 127640 6040 135960 6060
rect 137640 25740 145960 25760
rect 137640 6060 137660 25740
rect 145940 6060 145960 25740
rect 137640 6040 145960 6060
rect 147640 25740 155960 25760
rect 147640 6060 147660 25740
rect 155940 6060 155960 25740
rect 147640 6040 155960 6060
rect 157640 25740 165960 25760
rect 157640 6060 157660 25740
rect 165940 6060 165960 25740
rect 157640 6040 165960 6060
rect 167640 25740 175960 25760
rect 167640 6060 167660 25740
rect 175940 6060 175960 25740
rect 167640 6040 175960 6060
rect 177640 25740 185960 25760
rect 177640 6060 177660 25740
rect 185940 6060 185960 25740
rect 177640 6040 185960 6060
rect 187640 25740 195960 25760
rect 187640 6060 187660 25740
rect 195940 6060 195960 25740
rect 187640 6040 195960 6060
rect 197640 25740 205960 25760
rect 197640 6060 197660 25740
rect 205940 6060 205960 25740
rect 197640 6040 205960 6060
rect 207640 25740 215960 25760
rect 207640 6060 207660 25740
rect 215940 6060 215960 25740
rect 207640 6040 215960 6060
rect 217640 25740 225960 25760
rect 217640 6060 217660 25740
rect 225940 6060 225960 25740
rect 217640 6040 225960 6060
rect 227640 25740 235960 25760
rect 227640 6060 227660 25740
rect 235940 6060 235960 25740
rect 227640 6040 235960 6060
rect 237640 25740 245960 25760
rect 237640 6060 237660 25740
rect 245940 6060 245960 25740
rect 237640 6040 245960 6060
rect 247640 25740 255960 25760
rect 247640 6060 247660 25740
rect 255940 6060 255960 25740
rect 247640 6040 255960 6060
rect 257640 25740 265960 25760
rect 257640 6060 257660 25740
rect 265940 6060 265960 25740
rect 257640 6040 265960 6060
rect 267640 25740 275960 25760
rect 267640 6060 267660 25740
rect 275940 6060 275960 25740
rect 267640 6040 275960 6060
rect 277640 25740 285960 25760
rect 277640 6060 277660 25740
rect 285940 6060 285960 25740
rect 277640 6040 285960 6060
<< mimcapcontact >>
rect 46060 26260 54340 45940
rect 56060 26260 64340 45940
rect 66060 26260 74340 45940
rect 76060 26260 84340 45940
rect 86060 26260 94340 45940
rect 96060 26260 104340 45940
rect 106060 26260 114340 45940
rect 116060 26260 124340 45940
rect 126060 26260 134340 45940
rect 136060 26260 144340 45940
rect 146060 26260 154340 45940
rect 156060 26260 164340 45940
rect 166060 26260 174340 45940
rect 176060 26260 184340 45940
rect 186060 26260 194340 45940
rect 196060 26260 204340 45940
rect 206060 26260 214340 45940
rect 216060 26260 224340 45940
rect 226060 26260 234340 45940
rect 236060 26260 244340 45940
rect 246060 26260 254340 45940
rect 256060 26260 264340 45940
rect 266060 26260 274340 45940
rect 276060 26260 284340 45940
rect 47660 6060 55940 25740
rect 57660 6060 65940 25740
rect 67660 6060 75940 25740
rect 77660 6060 85940 25740
rect 87660 6060 95940 25740
rect 97660 6060 105940 25740
rect 107660 6060 115940 25740
rect 117660 6060 125940 25740
rect 127660 6060 135940 25740
rect 137660 6060 145940 25740
rect 147660 6060 155940 25740
rect 157660 6060 165940 25740
rect 167660 6060 175940 25740
rect 177660 6060 185940 25740
rect 187660 6060 195940 25740
rect 197660 6060 205940 25740
rect 207660 6060 215940 25740
rect 217660 6060 225940 25740
rect 227660 6060 235940 25740
rect 237660 6060 245940 25740
rect 247660 6060 255940 25740
rect 257660 6060 265940 25740
rect 267660 6060 275940 25740
rect 277660 6060 285940 25740
<< metal4 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46200 286000 46240
rect 46000 45940 54400 46200
rect 46000 26260 46060 45940
rect 54340 26260 54400 45940
rect 46000 26200 54400 26260
rect 56000 45940 64400 46200
rect 56000 26260 56060 45940
rect 64340 26260 64400 45940
rect 56000 26200 64400 26260
rect 66000 45940 74400 46200
rect 66000 26260 66060 45940
rect 74340 26260 74400 45940
rect 66000 26200 74400 26260
rect 76000 45940 84400 46200
rect 76000 26260 76060 45940
rect 84340 26260 84400 45940
rect 76000 26200 84400 26260
rect 86000 45940 94400 46200
rect 86000 26260 86060 45940
rect 94340 26260 94400 45940
rect 86000 26200 94400 26260
rect 96000 45940 104400 46200
rect 96000 26260 96060 45940
rect 104340 26260 104400 45940
rect 96000 26200 104400 26260
rect 106000 45940 114400 46200
rect 106000 26260 106060 45940
rect 114340 26260 114400 45940
rect 106000 26200 114400 26260
rect 116000 45940 124400 46200
rect 116000 26260 116060 45940
rect 124340 26260 124400 45940
rect 116000 26200 124400 26260
rect 126000 45940 134400 46200
rect 126000 26260 126060 45940
rect 134340 26260 134400 45940
rect 126000 26200 134400 26260
rect 136000 45940 144400 46200
rect 136000 26260 136060 45940
rect 144340 26260 144400 45940
rect 136000 26200 144400 26260
rect 146000 45940 154400 46200
rect 146000 26260 146060 45940
rect 154340 26260 154400 45940
rect 146000 26200 154400 26260
rect 156000 45940 164400 46200
rect 156000 26260 156060 45940
rect 164340 26260 164400 45940
rect 156000 26200 164400 26260
rect 166000 45940 174400 46200
rect 166000 26260 166060 45940
rect 174340 26260 174400 45940
rect 166000 26200 174400 26260
rect 176000 45940 184400 46200
rect 176000 26260 176060 45940
rect 184340 26260 184400 45940
rect 176000 26200 184400 26260
rect 186000 45940 194400 46200
rect 186000 26260 186060 45940
rect 194340 26260 194400 45940
rect 186000 26200 194400 26260
rect 196000 45940 204400 46200
rect 196000 26260 196060 45940
rect 204340 26260 204400 45940
rect 196000 26200 204400 26260
rect 206000 45940 214400 46200
rect 206000 26260 206060 45940
rect 214340 26260 214400 45940
rect 206000 26200 214400 26260
rect 216000 45940 224400 46200
rect 216000 26260 216060 45940
rect 224340 26260 224400 45940
rect 216000 26200 224400 26260
rect 226000 45940 234400 46200
rect 226000 26260 226060 45940
rect 234340 26260 234400 45940
rect 226000 26200 234400 26260
rect 236000 45940 244400 46200
rect 236000 26260 236060 45940
rect 244340 26260 244400 45940
rect 236000 26200 244400 26260
rect 246000 45940 254400 46200
rect 246000 26260 246060 45940
rect 254340 26260 254400 45940
rect 246000 26200 254400 26260
rect 256000 45940 264400 46200
rect 256000 26260 256060 45940
rect 264340 26260 264400 45940
rect 256000 26200 264400 26260
rect 266000 45940 274400 46200
rect 266000 26260 266060 45940
rect 274340 26260 274400 45940
rect 266000 26200 274400 26260
rect 276000 45940 284400 46200
rect 276000 26260 276060 45940
rect 284340 26260 284400 45940
rect 276000 26200 284400 26260
rect 47600 25800 54400 26200
rect 57600 25800 64400 26200
rect 67600 25800 74400 26200
rect 77600 25800 84400 26200
rect 87600 25800 94400 26200
rect 97600 25800 104400 26200
rect 107600 25800 114400 26200
rect 117600 25800 124400 26200
rect 127600 25800 134400 26200
rect 137600 25800 144400 26200
rect 147600 25800 154400 26200
rect 157600 25800 164400 26200
rect 167600 25800 174400 26200
rect 177600 25800 184400 26200
rect 187600 25800 194400 26200
rect 197600 25800 204400 26200
rect 207600 25800 214400 26200
rect 217600 25800 224400 26200
rect 227600 25800 234400 26200
rect 237600 25800 244400 26200
rect 247600 25800 254400 26200
rect 257600 25800 264400 26200
rect 267600 25800 274400 26200
rect 277600 25800 284400 26200
rect 47600 25740 56000 25800
rect 47600 6060 47660 25740
rect 55940 6060 56000 25740
rect 47600 6000 56000 6060
rect 57600 25740 66000 25800
rect 57600 6060 57660 25740
rect 65940 6060 66000 25740
rect 57600 6000 66000 6060
rect 67600 25740 76000 25800
rect 67600 6060 67660 25740
rect 75940 6060 76000 25740
rect 67600 6000 76000 6060
rect 77600 25740 86000 25800
rect 77600 6060 77660 25740
rect 85940 6060 86000 25740
rect 77600 6000 86000 6060
rect 87600 25740 96000 25800
rect 87600 6060 87660 25740
rect 95940 6060 96000 25740
rect 87600 6000 96000 6060
rect 97600 25740 106000 25800
rect 97600 6060 97660 25740
rect 105940 6060 106000 25740
rect 97600 6000 106000 6060
rect 107600 25740 116000 25800
rect 107600 6060 107660 25740
rect 115940 6060 116000 25740
rect 107600 6000 116000 6060
rect 117600 25740 126000 25800
rect 117600 6060 117660 25740
rect 125940 6060 126000 25740
rect 117600 6000 126000 6060
rect 127600 25740 136000 25800
rect 127600 6060 127660 25740
rect 135940 6060 136000 25740
rect 127600 6000 136000 6060
rect 137600 25740 146000 25800
rect 137600 6060 137660 25740
rect 145940 6060 146000 25740
rect 137600 6000 146000 6060
rect 147600 25740 156000 25800
rect 147600 6060 147660 25740
rect 155940 6060 156000 25740
rect 147600 6000 156000 6060
rect 157600 25740 166000 25800
rect 157600 6060 157660 25740
rect 165940 6060 166000 25740
rect 157600 6000 166000 6060
rect 167600 25740 176000 25800
rect 167600 6060 167660 25740
rect 175940 6060 176000 25740
rect 167600 6000 176000 6060
rect 177600 25740 186000 25800
rect 177600 6060 177660 25740
rect 185940 6060 186000 25740
rect 177600 6000 186000 6060
rect 187600 25740 196000 25800
rect 187600 6060 187660 25740
rect 195940 6060 196000 25740
rect 187600 6000 196000 6060
rect 197600 25740 206000 25800
rect 197600 6060 197660 25740
rect 205940 6060 206000 25740
rect 197600 6000 206000 6060
rect 207600 25740 216000 25800
rect 207600 6060 207660 25740
rect 215940 6060 216000 25740
rect 207600 6000 216000 6060
rect 217600 25740 226000 25800
rect 217600 6060 217660 25740
rect 225940 6060 226000 25740
rect 217600 6000 226000 6060
rect 227600 25740 236000 25800
rect 227600 6060 227660 25740
rect 235940 6060 236000 25740
rect 227600 6000 236000 6060
rect 237600 25740 246000 25800
rect 237600 6060 237660 25740
rect 245940 6060 246000 25740
rect 237600 6000 246000 6060
rect 247600 25740 256000 25800
rect 247600 6060 247660 25740
rect 255940 6060 256000 25740
rect 247600 6000 256000 6060
rect 257600 25740 266000 25800
rect 257600 6060 257660 25740
rect 265940 6060 266000 25740
rect 257600 6000 266000 6060
rect 267600 25740 276000 25800
rect 267600 6060 267660 25740
rect 275940 6060 276000 25740
rect 267600 6000 276000 6060
rect 277600 25740 286000 25800
rect 277600 6060 277660 25740
rect 285940 6060 286000 25740
rect 277600 6000 286000 6060
rect 46000 5760 286000 5800
rect 46000 5440 47000 5760
rect 55960 5440 57000 5760
rect 65960 5440 67000 5760
rect 75960 5440 77000 5760
rect 85960 5440 87000 5760
rect 95960 5440 97000 5760
rect 105960 5440 107000 5760
rect 115960 5440 117000 5760
rect 125960 5440 127000 5760
rect 135960 5440 137000 5760
rect 145960 5440 147000 5760
rect 155960 5440 157000 5760
rect 165960 5440 167000 5760
rect 175960 5440 177000 5760
rect 185960 5440 187000 5760
rect 195960 5440 197000 5760
rect 205960 5440 207000 5760
rect 215960 5440 217000 5760
rect 225960 5440 227000 5760
rect 235960 5440 237000 5760
rect 245960 5440 247000 5760
rect 255960 5440 257000 5760
rect 265960 5440 267000 5760
rect 275960 5440 277000 5760
rect 285960 5440 286000 5760
rect 46000 5400 286000 5440
<< via4 >>
rect 47000 46240 55000 46560
rect 57000 46240 65000 46560
rect 67000 46240 75000 46560
rect 77000 46240 85000 46560
rect 87000 46240 95000 46560
rect 97000 46240 105000 46560
rect 107000 46240 115000 46560
rect 117000 46240 125000 46560
rect 127000 46240 135000 46560
rect 137000 46240 145000 46560
rect 147000 46240 155000 46560
rect 157000 46240 165000 46560
rect 167000 46240 175000 46560
rect 177000 46240 185000 46560
rect 187000 46240 195000 46560
rect 197000 46240 205000 46560
rect 207000 46240 215000 46560
rect 217000 46240 225000 46560
rect 227000 46240 235000 46560
rect 237000 46240 245000 46560
rect 247000 46240 255000 46560
rect 257000 46240 265000 46560
rect 267000 46240 275000 46560
rect 277000 46240 285000 46560
rect 47000 5440 55000 5760
rect 57000 5440 65000 5760
rect 67000 5440 75000 5760
rect 77000 5440 85000 5760
rect 87000 5440 95000 5760
rect 97000 5440 105000 5760
rect 107000 5440 115000 5760
rect 117000 5440 125000 5760
rect 127000 5440 135000 5760
rect 137000 5440 145000 5760
rect 147000 5440 155000 5760
rect 157000 5440 165000 5760
rect 167000 5440 175000 5760
rect 177000 5440 185000 5760
rect 187000 5440 195000 5760
rect 197000 5440 205000 5760
rect 207000 5440 215000 5760
rect 217000 5440 225000 5760
rect 227000 5440 235000 5760
rect 237000 5440 245000 5760
rect 247000 5440 255000 5760
rect 257000 5440 265000 5760
rect 267000 5440 275000 5760
rect 277000 5440 285000 5760
<< mimcap2 >>
rect 46040 45940 54360 45960
rect 46040 26260 46060 45940
rect 54340 26260 54360 45940
rect 46040 26240 54360 26260
rect 56040 45940 64360 45960
rect 56040 26260 56060 45940
rect 64340 26260 64360 45940
rect 56040 26240 64360 26260
rect 66040 45940 74360 45960
rect 66040 26260 66060 45940
rect 74340 26260 74360 45940
rect 66040 26240 74360 26260
rect 76040 45940 84360 45960
rect 76040 26260 76060 45940
rect 84340 26260 84360 45940
rect 76040 26240 84360 26260
rect 86040 45940 94360 45960
rect 86040 26260 86060 45940
rect 94340 26260 94360 45940
rect 86040 26240 94360 26260
rect 96040 45940 104360 45960
rect 96040 26260 96060 45940
rect 104340 26260 104360 45940
rect 96040 26240 104360 26260
rect 106040 45940 114360 45960
rect 106040 26260 106060 45940
rect 114340 26260 114360 45940
rect 106040 26240 114360 26260
rect 116040 45940 124360 45960
rect 116040 26260 116060 45940
rect 124340 26260 124360 45940
rect 116040 26240 124360 26260
rect 126040 45940 134360 45960
rect 126040 26260 126060 45940
rect 134340 26260 134360 45940
rect 126040 26240 134360 26260
rect 136040 45940 144360 45960
rect 136040 26260 136060 45940
rect 144340 26260 144360 45940
rect 136040 26240 144360 26260
rect 146040 45940 154360 45960
rect 146040 26260 146060 45940
rect 154340 26260 154360 45940
rect 146040 26240 154360 26260
rect 156040 45940 164360 45960
rect 156040 26260 156060 45940
rect 164340 26260 164360 45940
rect 156040 26240 164360 26260
rect 166040 45940 174360 45960
rect 166040 26260 166060 45940
rect 174340 26260 174360 45940
rect 166040 26240 174360 26260
rect 176040 45940 184360 45960
rect 176040 26260 176060 45940
rect 184340 26260 184360 45940
rect 176040 26240 184360 26260
rect 186040 45940 194360 45960
rect 186040 26260 186060 45940
rect 194340 26260 194360 45940
rect 186040 26240 194360 26260
rect 196040 45940 204360 45960
rect 196040 26260 196060 45940
rect 204340 26260 204360 45940
rect 196040 26240 204360 26260
rect 206040 45940 214360 45960
rect 206040 26260 206060 45940
rect 214340 26260 214360 45940
rect 206040 26240 214360 26260
rect 216040 45940 224360 45960
rect 216040 26260 216060 45940
rect 224340 26260 224360 45940
rect 216040 26240 224360 26260
rect 226040 45940 234360 45960
rect 226040 26260 226060 45940
rect 234340 26260 234360 45940
rect 226040 26240 234360 26260
rect 236040 45940 244360 45960
rect 236040 26260 236060 45940
rect 244340 26260 244360 45940
rect 236040 26240 244360 26260
rect 246040 45940 254360 45960
rect 246040 26260 246060 45940
rect 254340 26260 254360 45940
rect 246040 26240 254360 26260
rect 256040 45940 264360 45960
rect 256040 26260 256060 45940
rect 264340 26260 264360 45940
rect 256040 26240 264360 26260
rect 266040 45940 274360 45960
rect 266040 26260 266060 45940
rect 274340 26260 274360 45940
rect 266040 26240 274360 26260
rect 276040 45940 284360 45960
rect 276040 26260 276060 45940
rect 284340 26260 284360 45940
rect 276040 26240 284360 26260
rect 47640 25740 55960 25760
rect 47640 6060 47660 25740
rect 55940 6060 55960 25740
rect 47640 6040 55960 6060
rect 57640 25740 65960 25760
rect 57640 6060 57660 25740
rect 65940 6060 65960 25740
rect 57640 6040 65960 6060
rect 67640 25740 75960 25760
rect 67640 6060 67660 25740
rect 75940 6060 75960 25740
rect 67640 6040 75960 6060
rect 77640 25740 85960 25760
rect 77640 6060 77660 25740
rect 85940 6060 85960 25740
rect 77640 6040 85960 6060
rect 87640 25740 95960 25760
rect 87640 6060 87660 25740
rect 95940 6060 95960 25740
rect 87640 6040 95960 6060
rect 97640 25740 105960 25760
rect 97640 6060 97660 25740
rect 105940 6060 105960 25740
rect 97640 6040 105960 6060
rect 107640 25740 115960 25760
rect 107640 6060 107660 25740
rect 115940 6060 115960 25740
rect 107640 6040 115960 6060
rect 117640 25740 125960 25760
rect 117640 6060 117660 25740
rect 125940 6060 125960 25740
rect 117640 6040 125960 6060
rect 127640 25740 135960 25760
rect 127640 6060 127660 25740
rect 135940 6060 135960 25740
rect 127640 6040 135960 6060
rect 137640 25740 145960 25760
rect 137640 6060 137660 25740
rect 145940 6060 145960 25740
rect 137640 6040 145960 6060
rect 147640 25740 155960 25760
rect 147640 6060 147660 25740
rect 155940 6060 155960 25740
rect 147640 6040 155960 6060
rect 157640 25740 165960 25760
rect 157640 6060 157660 25740
rect 165940 6060 165960 25740
rect 157640 6040 165960 6060
rect 167640 25740 175960 25760
rect 167640 6060 167660 25740
rect 175940 6060 175960 25740
rect 167640 6040 175960 6060
rect 177640 25740 185960 25760
rect 177640 6060 177660 25740
rect 185940 6060 185960 25740
rect 177640 6040 185960 6060
rect 187640 25740 195960 25760
rect 187640 6060 187660 25740
rect 195940 6060 195960 25740
rect 187640 6040 195960 6060
rect 197640 25740 205960 25760
rect 197640 6060 197660 25740
rect 205940 6060 205960 25740
rect 197640 6040 205960 6060
rect 207640 25740 215960 25760
rect 207640 6060 207660 25740
rect 215940 6060 215960 25740
rect 207640 6040 215960 6060
rect 217640 25740 225960 25760
rect 217640 6060 217660 25740
rect 225940 6060 225960 25740
rect 217640 6040 225960 6060
rect 227640 25740 235960 25760
rect 227640 6060 227660 25740
rect 235940 6060 235960 25740
rect 227640 6040 235960 6060
rect 237640 25740 245960 25760
rect 237640 6060 237660 25740
rect 245940 6060 245960 25740
rect 237640 6040 245960 6060
rect 247640 25740 255960 25760
rect 247640 6060 247660 25740
rect 255940 6060 255960 25740
rect 247640 6040 255960 6060
rect 257640 25740 265960 25760
rect 257640 6060 257660 25740
rect 265940 6060 265960 25740
rect 257640 6040 265960 6060
rect 267640 25740 275960 25760
rect 267640 6060 267660 25740
rect 275940 6060 275960 25740
rect 267640 6040 275960 6060
rect 277640 25740 285960 25760
rect 277640 6060 277660 25740
rect 285940 6060 285960 25740
rect 277640 6040 285960 6060
<< mimcap2contact >>
rect 46060 26260 54340 45940
rect 56060 26260 64340 45940
rect 66060 26260 74340 45940
rect 76060 26260 84340 45940
rect 86060 26260 94340 45940
rect 96060 26260 104340 45940
rect 106060 26260 114340 45940
rect 116060 26260 124340 45940
rect 126060 26260 134340 45940
rect 136060 26260 144340 45940
rect 146060 26260 154340 45940
rect 156060 26260 164340 45940
rect 166060 26260 174340 45940
rect 176060 26260 184340 45940
rect 186060 26260 194340 45940
rect 196060 26260 204340 45940
rect 206060 26260 214340 45940
rect 216060 26260 224340 45940
rect 226060 26260 234340 45940
rect 236060 26260 244340 45940
rect 246060 26260 254340 45940
rect 256060 26260 264340 45940
rect 266060 26260 274340 45940
rect 276060 26260 284340 45940
rect 47660 6060 55940 25740
rect 57660 6060 65940 25740
rect 67660 6060 75940 25740
rect 77660 6060 85940 25740
rect 87660 6060 95940 25740
rect 97660 6060 105940 25740
rect 107660 6060 115940 25740
rect 117660 6060 125940 25740
rect 127660 6060 135940 25740
rect 137660 6060 145940 25740
rect 147660 6060 155940 25740
rect 157660 6060 165940 25740
rect 167660 6060 175940 25740
rect 177660 6060 185940 25740
rect 187660 6060 195940 25740
rect 197660 6060 205940 25740
rect 207660 6060 215940 25740
rect 217660 6060 225940 25740
rect 227660 6060 235940 25740
rect 237660 6060 245940 25740
rect 247660 6060 255940 25740
rect 257660 6060 265940 25740
rect 267660 6060 275940 25740
rect 277660 6060 285940 25740
<< metal5 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46000 286000 46240
rect 46000 45940 54400 46000
rect 46000 26260 46060 45940
rect 54340 26260 54400 45940
rect 46000 26200 54400 26260
rect 56000 45940 64400 46000
rect 56000 26260 56060 45940
rect 64340 26260 64400 45940
rect 56000 26200 64400 26260
rect 66000 45940 74400 46000
rect 66000 26260 66060 45940
rect 74340 26260 74400 45940
rect 66000 26200 74400 26260
rect 76000 45940 84400 46000
rect 76000 26260 76060 45940
rect 84340 26260 84400 45940
rect 76000 26200 84400 26260
rect 86000 45940 94400 46000
rect 86000 26260 86060 45940
rect 94340 26260 94400 45940
rect 86000 26200 94400 26260
rect 96000 45940 104400 46000
rect 96000 26260 96060 45940
rect 104340 26260 104400 45940
rect 96000 26200 104400 26260
rect 106000 45940 114400 46000
rect 106000 26260 106060 45940
rect 114340 26260 114400 45940
rect 106000 26200 114400 26260
rect 116000 45940 124400 46000
rect 116000 26260 116060 45940
rect 124340 26260 124400 45940
rect 116000 26200 124400 26260
rect 126000 45940 134400 46000
rect 126000 26260 126060 45940
rect 134340 26260 134400 45940
rect 126000 26200 134400 26260
rect 136000 45940 144400 46000
rect 136000 26260 136060 45940
rect 144340 26260 144400 45940
rect 136000 26200 144400 26260
rect 146000 45940 154400 46000
rect 146000 26260 146060 45940
rect 154340 26260 154400 45940
rect 146000 26200 154400 26260
rect 156000 45940 164400 46000
rect 156000 26260 156060 45940
rect 164340 26260 164400 45940
rect 156000 26200 164400 26260
rect 166000 45940 174400 46000
rect 166000 26260 166060 45940
rect 174340 26260 174400 45940
rect 166000 26200 174400 26260
rect 176000 45940 184400 46000
rect 176000 26260 176060 45940
rect 184340 26260 184400 45940
rect 176000 26200 184400 26260
rect 186000 45940 194400 46000
rect 186000 26260 186060 45940
rect 194340 26260 194400 45940
rect 186000 26200 194400 26260
rect 196000 45940 204400 46000
rect 196000 26260 196060 45940
rect 204340 26260 204400 45940
rect 196000 26200 204400 26260
rect 206000 45940 214400 46000
rect 206000 26260 206060 45940
rect 214340 26260 214400 45940
rect 206000 26200 214400 26260
rect 216000 45940 224400 46000
rect 216000 26260 216060 45940
rect 224340 26260 224400 45940
rect 216000 26200 224400 26260
rect 226000 45940 234400 46000
rect 226000 26260 226060 45940
rect 234340 26260 234400 45940
rect 226000 26200 234400 26260
rect 236000 45940 244400 46000
rect 236000 26260 236060 45940
rect 244340 26260 244400 45940
rect 236000 26200 244400 26260
rect 246000 45940 254400 46000
rect 246000 26260 246060 45940
rect 254340 26260 254400 45940
rect 246000 26200 254400 26260
rect 256000 45940 264400 46000
rect 256000 26260 256060 45940
rect 264340 26260 264400 45940
rect 256000 26200 264400 26260
rect 266000 45940 274400 46000
rect 266000 26260 266060 45940
rect 274340 26260 274400 45940
rect 266000 26200 274400 26260
rect 276000 45940 284400 46000
rect 276000 26260 276060 45940
rect 284340 26260 284400 45940
rect 276000 26200 284400 26260
rect 47600 25800 54400 26200
rect 57600 25800 64400 26200
rect 67600 25800 74400 26200
rect 77600 25800 84400 26200
rect 87600 25800 94400 26200
rect 97600 25800 104400 26200
rect 107600 25800 114400 26200
rect 117600 25800 124400 26200
rect 127600 25800 134400 26200
rect 137600 25800 144400 26200
rect 147600 25800 154400 26200
rect 157600 25800 164400 26200
rect 167600 25800 174400 26200
rect 177600 25800 184400 26200
rect 187600 25800 194400 26200
rect 197600 25800 204400 26200
rect 207600 25800 214400 26200
rect 217600 25800 224400 26200
rect 227600 25800 234400 26200
rect 237600 25800 244400 26200
rect 247600 25800 254400 26200
rect 257600 25800 264400 26200
rect 267600 25800 274400 26200
rect 277600 25800 284400 26200
rect 47600 25740 56000 25800
rect 47600 6060 47660 25740
rect 55940 6060 56000 25740
rect 47600 6000 56000 6060
rect 57600 25740 66000 25800
rect 57600 6060 57660 25740
rect 65940 6060 66000 25740
rect 57600 6000 66000 6060
rect 67600 25740 76000 25800
rect 67600 6060 67660 25740
rect 75940 6060 76000 25740
rect 67600 6000 76000 6060
rect 77600 25740 86000 25800
rect 77600 6060 77660 25740
rect 85940 6060 86000 25740
rect 77600 6000 86000 6060
rect 87600 25740 96000 25800
rect 87600 6060 87660 25740
rect 95940 6060 96000 25740
rect 87600 6000 96000 6060
rect 97600 25740 106000 25800
rect 97600 6060 97660 25740
rect 105940 6060 106000 25740
rect 97600 6000 106000 6060
rect 107600 25740 116000 25800
rect 107600 6060 107660 25740
rect 115940 6060 116000 25740
rect 107600 6000 116000 6060
rect 117600 25740 126000 25800
rect 117600 6060 117660 25740
rect 125940 6060 126000 25740
rect 117600 6000 126000 6060
rect 127600 25740 136000 25800
rect 127600 6060 127660 25740
rect 135940 6060 136000 25740
rect 127600 6000 136000 6060
rect 137600 25740 146000 25800
rect 137600 6060 137660 25740
rect 145940 6060 146000 25740
rect 137600 6000 146000 6060
rect 147600 25740 156000 25800
rect 147600 6060 147660 25740
rect 155940 6060 156000 25740
rect 147600 6000 156000 6060
rect 157600 25740 166000 25800
rect 157600 6060 157660 25740
rect 165940 6060 166000 25740
rect 157600 6000 166000 6060
rect 167600 25740 176000 25800
rect 167600 6060 167660 25740
rect 175940 6060 176000 25740
rect 167600 6000 176000 6060
rect 177600 25740 186000 25800
rect 177600 6060 177660 25740
rect 185940 6060 186000 25740
rect 177600 6000 186000 6060
rect 187600 25740 196000 25800
rect 187600 6060 187660 25740
rect 195940 6060 196000 25740
rect 187600 6000 196000 6060
rect 197600 25740 206000 25800
rect 197600 6060 197660 25740
rect 205940 6060 206000 25740
rect 197600 6000 206000 6060
rect 207600 25740 216000 25800
rect 207600 6060 207660 25740
rect 215940 6060 216000 25740
rect 207600 6000 216000 6060
rect 217600 25740 226000 25800
rect 217600 6060 217660 25740
rect 225940 6060 226000 25740
rect 217600 6000 226000 6060
rect 227600 25740 236000 25800
rect 227600 6060 227660 25740
rect 235940 6060 236000 25740
rect 227600 6000 236000 6060
rect 237600 25740 246000 25800
rect 237600 6060 237660 25740
rect 245940 6060 246000 25740
rect 237600 6000 246000 6060
rect 247600 25740 256000 25800
rect 247600 6060 247660 25740
rect 255940 6060 256000 25740
rect 247600 6000 256000 6060
rect 257600 25740 266000 25800
rect 257600 6060 257660 25740
rect 265940 6060 266000 25740
rect 257600 6000 266000 6060
rect 267600 25740 276000 25800
rect 267600 6060 267660 25740
rect 275940 6060 276000 25740
rect 267600 6000 276000 6060
rect 277600 25740 286000 25800
rect 277600 6060 277660 25740
rect 285940 6060 286000 25740
rect 277600 6000 286000 6060
rect 46000 5760 286000 6000
rect 46000 5440 47000 5760
rect 55000 5440 57000 5760
rect 65000 5440 67000 5760
rect 75000 5440 77000 5760
rect 85000 5440 87000 5760
rect 95000 5440 97000 5760
rect 105000 5440 107000 5760
rect 115000 5440 117000 5760
rect 125000 5440 127000 5760
rect 135000 5440 137000 5760
rect 145000 5440 147000 5760
rect 155000 5440 157000 5760
rect 165000 5440 167000 5760
rect 175000 5440 177000 5760
rect 185000 5440 187000 5760
rect 195000 5440 197000 5760
rect 205000 5440 207000 5760
rect 215000 5440 217000 5760
rect 225000 5440 227000 5760
rect 235000 5440 237000 5760
rect 245000 5440 247000 5760
rect 255000 5440 257000 5760
rect 265000 5440 267000 5760
rect 275000 5440 277000 5760
rect 285000 5440 286000 5760
rect 46000 5400 286000 5440
use sky130_fd_pr__res_xhigh_po_0p35_FE9J4G  sky130_fd_pr__res_xhigh_po_0p35_FE9J4G_0
timestamp 1672019510
transform 0 1 56598 -1 0 48201
box -201 -10598 201 10598
<< end >>
