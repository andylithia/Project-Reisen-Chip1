magic
tech sky130A
magscale 1 2
timestamp 1672475812
<< metal2 >>
rect -1504 32 188 88
rect -1504 -1258 -1448 32
rect 312 -12 368 88
rect -1228 -68 368 -12
rect -1228 -1268 -1172 -68
rect 552 -112 608 88
rect -952 -168 608 -112
rect -952 -1288 -896 -168
rect 732 -212 788 88
rect 972 -72 1028 88
rect -676 -268 788 -212
rect 832 -128 1028 -72
rect -676 -1208 -620 -268
rect 832 -312 888 -128
rect 1152 -192 1208 68
rect 1412 -52 1468 108
rect -400 -368 888 -312
rect 952 -248 1208 -192
rect 1252 -108 1468 -52
rect -400 -1288 -344 -368
rect 952 -412 1008 -248
rect 1252 -312 1308 -108
rect 1572 -152 1628 88
rect 1832 -52 1888 68
rect -124 -468 1008 -412
rect 1052 -368 1308 -312
rect 1352 -208 1628 -152
rect 1672 -108 1888 -52
rect -124 -1208 -68 -468
rect 1052 -512 1108 -368
rect 1352 -432 1408 -208
rect 1672 -252 1728 -108
rect 1992 -152 2048 88
rect 2252 -32 2308 68
rect 152 -568 1108 -512
rect 1152 -488 1408 -432
rect 1472 -308 1728 -252
rect 1772 -208 2048 -152
rect 2092 -88 2308 -32
rect 152 -1288 208 -568
rect 1152 -612 1208 -488
rect 1472 -532 1528 -308
rect 1772 -352 1828 -208
rect 2092 -252 2148 -88
rect 2412 -132 2468 108
rect 428 -668 1208 -612
rect 1272 -588 1528 -532
rect 1572 -408 1828 -352
rect 1872 -308 2148 -252
rect 2192 -188 2468 -132
rect 428 -1228 484 -668
rect 1272 -732 1328 -588
rect 1572 -632 1628 -408
rect 1872 -472 1928 -308
rect 2192 -352 2248 -188
rect 2672 -232 2728 88
rect 704 -788 1328 -732
rect 1372 -688 1628 -632
rect 1692 -528 1928 -472
rect 1972 -408 2248 -352
rect 2292 -288 2728 -232
rect 704 -1208 760 -788
rect 1372 -832 1428 -688
rect 1692 -732 1748 -528
rect 1972 -572 2028 -408
rect 2292 -452 2348 -288
rect 2832 -332 2888 88
rect 980 -888 1428 -832
rect 1492 -788 1748 -732
rect 1792 -628 2028 -572
rect 2072 -508 2348 -452
rect 2392 -388 2888 -332
rect 980 -1248 1036 -888
rect 1492 -932 1548 -788
rect 1792 -832 1848 -628
rect 2072 -672 2128 -508
rect 2392 -552 2448 -388
rect 3072 -432 3128 88
rect 2552 -488 3128 -432
rect 1256 -988 1548 -932
rect 1632 -888 1848 -832
rect 1892 -728 2128 -672
rect 2172 -608 2468 -552
rect 1256 -1188 1312 -988
rect 1632 -1072 1688 -888
rect 1892 -932 1948 -728
rect 2172 -772 2228 -608
rect 2552 -672 2608 -488
rect 3252 -532 3308 88
rect 3512 -112 3568 88
rect 1532 -1128 1688 -1072
rect 1808 -988 1948 -932
rect 2084 -828 2228 -772
rect 2360 -728 2608 -672
rect 2712 -588 3308 -532
rect 3352 -168 3568 -112
rect 1808 -1128 1864 -988
rect 2084 -1128 2140 -828
rect 2360 -1148 2416 -728
rect 2712 -772 2768 -588
rect 3352 -672 3408 -168
rect 3672 -232 3728 68
rect 3932 -32 3988 88
rect 2636 -828 2768 -772
rect 2912 -728 3408 -672
rect 3452 -288 3728 -232
rect 3772 -88 3988 -32
rect 2636 -1148 2692 -828
rect 2912 -1128 2968 -728
rect 3452 -792 3508 -288
rect 3772 -332 3828 -88
rect 4092 -152 4148 88
rect 4352 -52 4408 108
rect 3188 -848 3508 -792
rect 3572 -388 3828 -332
rect 3872 -208 4148 -152
rect 4232 -108 4408 -52
rect 3188 -1148 3244 -848
rect 3572 -912 3628 -388
rect 3872 -452 3928 -208
rect 4232 -252 4288 -108
rect 4512 -152 4568 68
rect 4772 -32 4828 88
rect 3464 -968 3628 -912
rect 3740 -508 3928 -452
rect 4016 -308 4288 -252
rect 4332 -208 4568 -152
rect 4652 -88 4828 -32
rect 3464 -1148 3520 -968
rect 3740 -1168 3796 -508
rect 4016 -1308 4072 -308
rect 4332 -392 4388 -208
rect 4652 -252 4708 -88
rect 4932 -132 4988 68
rect 5212 -132 5268 88
rect 4292 -448 4388 -392
rect 4568 -308 4708 -252
rect 4844 -188 4988 -132
rect 5120 -188 5268 -132
rect 4292 -1228 4348 -448
rect 4568 -1148 4624 -308
rect 4844 -1168 4900 -188
rect 5120 -1188 5176 -188
rect 5396 -1168 5452 68
rect 5592 -372 5648 88
rect 5592 -428 5728 -372
rect 5672 -1188 5728 -428
rect 5792 -892 5848 88
rect 6032 -792 6088 88
rect 6172 -692 6228 88
rect 6172 -748 6556 -692
rect 6032 -848 6280 -792
rect 5792 -948 6004 -892
rect 5948 -1108 6004 -948
rect 6224 -1188 6280 -848
rect 6500 -1188 6556 -748
rect 7292 -952 7348 68
rect 7452 -872 7508 88
rect 8532 -12 8588 88
rect 7880 -68 8588 -12
rect 7452 -928 7660 -872
rect 7292 -1008 7384 -952
rect 7328 -1248 7384 -1008
rect 7604 -1168 7660 -928
rect 7880 -1148 7936 -68
rect 8712 -132 8768 88
rect 9812 -32 9868 88
rect 8156 -188 8768 -132
rect 8832 -88 9868 -32
rect 8156 -1148 8212 -188
rect 8832 -252 8888 -88
rect 9992 -132 10048 68
rect 11072 -32 11128 108
rect 8432 -308 8888 -252
rect 8932 -188 10048 -132
rect 10332 -88 11128 -32
rect 8432 -1148 8488 -308
rect 8932 -352 8988 -188
rect 10332 -232 10388 -88
rect 11232 -132 11288 88
rect 12332 -32 12388 88
rect 8708 -408 8988 -352
rect 9072 -288 10388 -232
rect 10432 -188 11288 -132
rect 11472 -88 12388 -32
rect 8708 -1128 8764 -408
rect 9072 -472 9128 -288
rect 10432 -352 10488 -188
rect 11472 -232 11528 -88
rect 12492 -132 12548 68
rect 13592 -52 13648 88
rect 8984 -528 9128 -472
rect 9260 -408 10488 -352
rect 10552 -288 11528 -232
rect 11572 -188 12548 -132
rect 12872 -108 13648 -52
rect 8984 -1148 9040 -528
rect 9260 -1168 9316 -408
rect 10552 -452 10608 -288
rect 11572 -332 11628 -188
rect 12872 -232 12928 -108
rect 13772 -172 13828 68
rect 9536 -508 10608 -452
rect 10672 -388 11628 -332
rect 11712 -288 12928 -232
rect 12992 -228 13828 -172
rect 9536 -1228 9592 -508
rect 10672 -572 10728 -388
rect 11712 -452 11768 -288
rect 12992 -332 13048 -228
rect 14012 -272 14068 48
rect 9812 -628 10728 -572
rect 10792 -508 11768 -452
rect 11812 -388 13048 -332
rect 13112 -328 14068 -272
rect 9812 -1128 9868 -628
rect 10792 -672 10848 -508
rect 11812 -572 11868 -388
rect 13112 -452 13168 -328
rect 14172 -372 14228 88
rect 10088 -728 10848 -672
rect 10932 -628 11868 -572
rect 11912 -508 13168 -452
rect 13212 -428 14228 -372
rect 10088 -1148 10144 -728
rect 10932 -792 10988 -628
rect 11912 -692 11968 -508
rect 13212 -552 13268 -428
rect 10364 -848 10988 -792
rect 11112 -748 11968 -692
rect 12032 -608 13268 -552
rect 10364 -1248 10420 -848
rect 11112 -912 11168 -748
rect 12032 -792 12088 -608
rect 10640 -968 11168 -912
rect 11272 -848 12088 -792
rect 10640 -1168 10696 -968
rect 11272 -1052 11328 -848
rect 10916 -1108 11328 -1052
rect -2540 -31060 -2440 -30240
rect -1440 -31060 -1340 -30240
rect -340 -31060 -240 -30240
rect 780 -31060 880 -30240
rect 1880 -31060 1980 -30240
rect 2980 -31060 3080 -30240
rect 4080 -31060 4180 -30240
rect 5180 -31060 5280 -30240
rect 6300 -31060 6400 -30240
rect 7400 -31060 7500 -30240
rect 8500 -31060 8600 -30240
rect 9600 -31060 9700 -30240
rect 10720 -31060 10820 -30240
rect 11820 -31060 11920 -30240
<< metal3 >>
rect -1180 2910 -20 3020
rect -1180 2840 30 2910
rect -30 2830 30 2840
rect -860 2760 -100 2780
rect -860 2620 -840 2760
rect -560 2740 -100 2760
rect -560 2660 30 2740
rect -560 2620 -100 2660
rect -860 2600 -100 2620
rect -1180 2160 -40 2220
rect -1180 2080 30 2160
rect -1180 2040 -40 2080
rect -1180 1400 -40 1480
rect -1180 1320 30 1400
rect -1180 1300 -40 1320
rect 140 -10 220 30
rect 310 -10 390 30
rect 560 -10 640 30
<< via3 >>
rect -840 2620 -560 2760
<< metal4 >>
rect -1180 2760 -540 2780
rect -1180 2620 -840 2760
rect -560 2620 -540 2760
rect -1180 2320 -540 2620
rect -860 -2220 -540 2320
rect -860 -2240 8274 -2220
rect -860 -2540 11701 -2240
rect 1100 -5960 1420 -2540
rect 4527 -5480 4847 -2540
rect 7954 -2560 11701 -2540
rect 7954 -3818 8274 -2560
rect 11381 -3760 11701 -2560
rect -613 -29440 -293 -27540
rect 2814 -29440 3134 -28440
rect 6241 -29440 6561 -28440
rect 9668 -29440 9988 -27978
rect -2700 -29760 9988 -29440
use dac_2r_1  dac_2r_1_0
timestamp 1672475742
transform 1 0 2720 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_1
timestamp 1672475742
transform 1 0 -1060 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_2
timestamp 1672475742
transform 1 0 -640 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_3
timestamp 1672475742
transform 1 0 -220 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_4
timestamp 1672475742
transform 1 0 200 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_5
timestamp 1672475742
transform 1 0 620 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_6
timestamp 1672475742
transform 1 0 1040 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_7
timestamp 1672475742
transform 1 0 1460 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_8
timestamp 1672475742
transform 1 0 1880 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_9
timestamp 1672475742
transform 1 0 2300 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_11
timestamp 1672475742
transform 1 0 3140 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_12
timestamp 1672475742
transform 1 0 3560 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_13
timestamp 1672475742
transform 1 0 3980 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_14
timestamp 1672475742
transform 1 0 4400 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_15
timestamp 1672475742
transform 1 0 4820 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_16
timestamp 1672475742
transform 1 0 7340 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_17
timestamp 1672475742
transform 1 0 6080 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_18
timestamp 1672475742
transform 1 0 8600 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_19
timestamp 1672475742
transform 1 0 9860 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_20
timestamp 1672475742
transform 1 0 11120 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_21
timestamp 1672475742
transform 1 0 12800 0 1 -460
box 1060 450 1590 3370
use dac_2r_1  dac_2r_1_22
timestamp 1672475742
transform 1 0 12380 0 1 -460
box 1060 450 1590 3370
use dac_con  dac_con_0
timestamp 1672474575
transform 1 0 -3270 0 1 -31050
box 750 0 15166 30000
use dac_r_1  dac_r_1_0
timestamp 1672468680
transform 1 0 6500 0 1 -460
box 1060 558 2010 3370
use dac_r_1  dac_r_1_1
timestamp 1672468680
transform 1 0 5240 0 1 -460
box 1060 558 2010 3370
use dac_r_1  dac_r_1_2
timestamp 1672468680
transform 1 0 7760 0 1 -460
box 1060 558 2010 3370
use dac_r_1  dac_r_1_3
timestamp 1672468680
transform 1 0 9020 0 1 -460
box 1060 558 2010 3370
use dac_r_1  dac_r_1_4
timestamp 1672468680
transform 1 0 10280 0 1 -460
box 1060 558 2010 3370
use dac_r_1  dac_r_1_5
timestamp 1672468680
transform 1 0 11540 0 1 -460
box 1060 558 2010 3370
<< labels >>
rlabel metal3 -30 2830 30 2910 1 IOUT
port 1 n
rlabel metal3 -30 2660 30 2740 1 VSUB
port 2 n
rlabel metal3 -30 2080 30 2160 1 VHI
port 3 n
rlabel metal3 140 -10 220 30 1 SG15
port 4 n
rlabel metal3 310 -10 390 30 1 SO15
port 5 n
rlabel metal3 560 -10 640 30 1 SG14
port 6 n
rlabel metal4 -1180 2320 -860 2780 1 VLO
port 7 n
rlabel metal3 -1180 2840 -860 3020 1 IOUT
port 1 n
rlabel metal3 -1180 2040 -860 2220 1 VREF
port 8 n
rlabel metal4 -2700 -29760 -2540 -29440 1 VHI
port 3 n
rlabel metal2 -2540 -31060 -2440 -30240 1 TEST_MODE
port 9 n
rlabel metal2 -1440 -31060 -1340 -30240 1 RST_N
port 10 n
rlabel metal2 -340 -31060 -240 -30240 1 CLK
port 11 n
rlabel metal2 780 -31060 880 -30240 1 DIN9
port 12 n
rlabel metal2 1880 -31060 1980 -30240 1 DIN8
port 13 n
rlabel metal2 2980 -31060 3080 -30240 1 DIN7
port 14 n
rlabel metal2 4080 -31060 4180 -30240 1 DIN6
port 15 n
rlabel metal2 5180 -31060 5280 -30240 1 DIN5
port 16 n
rlabel metal2 6300 -31060 6400 -30240 1 DIN4
port 17 n
rlabel metal2 7400 -31060 7500 -30240 1 DIN3
port 18 n
rlabel metal2 8500 -31060 8600 -30240 1 DIN2
port 19 n
rlabel metal2 9600 -31060 9700 -30240 1 DIN1
port 20 n
rlabel metal2 10720 -31060 10820 -30240 1 DIN0
port 21 n
rlabel metal2 11820 -31060 11920 -30240 1 DUMMY
port 22 n
rlabel metal3 -1180 1300 -860 1480 1 VMID
port 23 n
<< end >>
