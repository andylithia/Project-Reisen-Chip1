magic
tech sky130B
magscale 1 2
timestamp 1668746166
<< metal1 >>
rect 207 569 259 585
rect 541 569 593 585
rect 359 501 441 507
rect 359 449 373 501
rect 425 449 441 501
rect 359 443 441 449
rect 319 395 379 415
rect 319 343 327 395
rect 319 323 379 343
rect 421 395 481 415
rect 473 343 481 395
rect 421 323 481 343
rect 207 249 259 265
rect 541 249 593 265
rect 207 197 275 249
rect 525 197 593 249
<< via1 >>
rect 207 265 259 569
rect 373 449 425 501
rect 327 343 379 395
rect 421 343 473 395
rect 541 265 593 569
rect 275 197 525 249
<< metal2 >>
rect 207 569 259 585
rect 541 569 593 585
rect 359 525 441 527
rect 359 469 371 525
rect 427 469 441 525
rect 359 449 373 469
rect 425 449 441 469
rect 359 443 441 449
rect 319 397 379 415
rect 319 341 323 397
rect 319 323 379 341
rect 421 397 481 415
rect 477 341 481 397
rect 421 323 481 341
rect 207 249 259 265
rect 541 249 593 265
rect 207 241 275 249
rect 525 241 593 249
rect 207 185 217 241
rect 583 185 593 241
rect 207 177 593 185
<< via2 >>
rect 371 501 427 525
rect 371 469 373 501
rect 373 469 425 501
rect 425 469 427 501
rect 323 395 379 397
rect 323 343 327 395
rect 327 343 379 395
rect 323 341 379 343
rect 421 395 477 397
rect 421 343 473 395
rect 473 343 477 395
rect 421 341 477 343
rect 217 197 275 241
rect 275 197 525 241
rect 525 197 583 241
rect 217 185 583 197
<< metal3 >>
rect 359 525 441 607
rect 359 469 371 525
rect 427 469 441 525
rect 359 463 441 469
rect 317 397 483 403
rect 317 341 323 397
rect 379 341 421 397
rect 477 341 483 397
rect 317 323 483 341
rect 207 241 593 249
rect 207 185 217 241
rect 583 185 593 241
rect 207 177 593 185
<< comment >>
rect 225 569 259 585
rect 541 569 575 585
rect 225 249 259 265
rect 541 249 575 265
rect 259 215 275 249
rect 525 215 541 249
use sky130_fd_pr__nfet_01v8_DA57K3  sky130_fd_pr__nfet_01v8_DA57K3_0
timestamp 1668741270
transform 1 0 400 0 1 400
box -211 -221 211 221
<< end >>
