magic
tech sky130A
magscale 1 2
timestamp 1671203110
<< viali >>
rect -128 -624 -94 -224
rect 1280 -624 1314 -224
rect 3885 -624 3919 -224
rect 5293 -624 5327 -224
rect 1553 -1740 1587 -1340
rect 3613 -1740 3647 -1340
rect -128 -2224 -94 -1824
rect 1280 -2224 1314 -1824
rect 3885 -2224 3919 -1824
rect 5293 -2224 5327 -1824
rect 1553 -3340 1587 -2940
rect 3613 -3340 3647 -2940
<< metal1 >>
rect 331 -42 383 -36
rect 331 -146 383 -94
rect 567 -42 619 -36
rect 567 -146 619 -94
rect 803 -42 855 -36
rect 803 -146 855 -94
rect 4344 -42 4396 -36
rect 4344 -146 4396 -94
rect 4580 -42 4632 -36
rect 4580 -146 4632 -94
rect 4816 -42 4868 -36
rect 4816 -146 4868 -94
rect -23 -192 91 -146
rect 151 -192 1035 -146
rect 1095 -192 1209 -146
rect -134 -224 -88 -212
rect -23 -224 29 -192
rect 1157 -224 1209 -192
rect 3990 -192 4104 -146
rect 4164 -192 5048 -146
rect 5108 -192 5222 -146
rect 1300 -212 1400 -200
rect 1274 -224 1400 -212
rect -134 -624 -128 -224
rect -94 -236 29 -224
rect -94 -624 -23 -236
rect -134 -636 -88 -624
rect -134 -1824 -88 -1812
rect -134 -2224 -128 -1824
rect -94 -2212 -23 -1824
rect -94 -2224 29 -2212
rect 95 -236 147 -224
rect 95 -2224 147 -2212
rect 213 -236 265 -224
rect 213 -2224 265 -2212
rect 331 -236 383 -224
rect 331 -2224 383 -2212
rect 449 -236 501 -224
rect 449 -2224 501 -2212
rect 567 -236 619 -224
rect 567 -2224 619 -2212
rect 685 -236 737 -224
rect 685 -2224 737 -2212
rect 803 -236 855 -224
rect 803 -2224 855 -2212
rect 921 -236 973 -224
rect 921 -2224 973 -2212
rect 1039 -236 1091 -224
rect 1039 -2224 1091 -2212
rect 1157 -236 1280 -224
rect 1209 -624 1280 -236
rect 1314 -300 1400 -224
rect 3800 -212 3900 -200
rect 3800 -224 3925 -212
rect 3990 -224 4042 -192
rect 5170 -224 5222 -192
rect 5287 -224 5333 -212
rect 3800 -300 3885 -224
rect 1314 -624 1560 -300
rect 1274 -636 1560 -624
rect 1300 -800 1560 -636
rect 1400 -1200 1560 -800
rect 3640 -624 3885 -300
rect 3919 -236 4042 -224
rect 3919 -624 3990 -236
rect 3640 -636 3925 -624
rect 3640 -800 3900 -636
rect 1400 -1340 1600 -1200
rect 1672 -1308 3483 -1262
rect 3640 -1328 3800 -800
rect 3607 -1340 3800 -1328
rect 1400 -1700 1553 -1340
rect 1300 -1740 1553 -1700
rect 1587 -1352 1710 -1340
rect 1587 -1740 1658 -1352
rect 1300 -1800 1600 -1740
rect 1300 -1812 1560 -1800
rect 1274 -1824 1560 -1812
rect 1209 -2212 1280 -1824
rect 1157 -2224 1280 -2212
rect 1314 -2224 1560 -1824
rect -134 -2236 -88 -2224
rect -23 -2256 29 -2224
rect 1157 -2256 1209 -2224
rect 1274 -2236 1560 -2224
rect -23 -2302 91 -2256
rect 151 -2302 1035 -2256
rect 1095 -2302 1209 -2256
rect 1300 -2300 1560 -2236
rect 1400 -2360 1560 -2300
rect 1400 -3580 1420 -2360
rect 1480 -2928 1560 -2360
rect 1480 -2940 1593 -2928
rect 1480 -3340 1553 -2940
rect 1587 -3328 1658 -2940
rect 1587 -3340 1710 -3328
rect 2116 -1352 2168 -1340
rect 2116 -3340 2168 -3328
rect 2574 -1352 2626 -1340
rect 2574 -3340 2626 -3328
rect 3032 -1352 3084 -1340
rect 3032 -3340 3084 -3328
rect 3490 -1352 3613 -1340
rect 3542 -1740 3613 -1352
rect 3647 -1700 3800 -1340
rect 3647 -1740 3900 -1700
rect 3607 -1752 3900 -1740
rect 3640 -1812 3900 -1752
rect 3640 -1824 3925 -1812
rect 3640 -2224 3885 -1824
rect 3919 -2212 3990 -1824
rect 3919 -2224 4042 -2212
rect 4108 -236 4160 -224
rect 4108 -2224 4160 -2212
rect 4226 -236 4278 -224
rect 4226 -2224 4278 -2212
rect 4344 -236 4396 -224
rect 4344 -2224 4396 -2212
rect 4462 -236 4514 -224
rect 4462 -2224 4514 -2212
rect 4580 -236 4632 -224
rect 4580 -2224 4632 -2212
rect 4698 -236 4750 -224
rect 4698 -2224 4750 -2212
rect 4816 -236 4868 -224
rect 4816 -2224 4868 -2212
rect 4934 -236 4986 -224
rect 4934 -2224 4986 -2212
rect 5052 -236 5104 -224
rect 5052 -2224 5104 -2212
rect 5170 -236 5293 -224
rect 5222 -624 5293 -236
rect 5327 -624 5333 -224
rect 5287 -636 5333 -624
rect 5287 -1824 5333 -1812
rect 5222 -2212 5293 -1824
rect 5170 -2224 5293 -2212
rect 5327 -2224 5333 -1824
rect 3640 -2236 3925 -2224
rect 3640 -2300 3900 -2236
rect 3990 -2256 4042 -2224
rect 5170 -2256 5222 -2224
rect 5287 -2236 5333 -2224
rect 3640 -2360 3800 -2300
rect 3990 -2302 4104 -2256
rect 4164 -2302 5048 -2256
rect 5108 -2302 5222 -2256
rect 3640 -2928 3720 -2360
rect 3607 -2940 3720 -2928
rect 3542 -3328 3613 -2940
rect 3490 -3340 3613 -3328
rect 3647 -3340 3720 -2940
rect 1480 -3352 1593 -3340
rect 3607 -3352 3720 -3340
rect 1480 -3580 1560 -3352
rect 1717 -3418 3483 -3372
rect 1400 -3600 1560 -3580
rect 3640 -3580 3720 -3352
rect 3780 -3580 3800 -2360
rect 3640 -3600 3800 -3580
<< via1 >>
rect 331 -94 383 -42
rect 567 -94 619 -42
rect 803 -94 855 -42
rect 4344 -94 4396 -42
rect 4580 -94 4632 -42
rect 4816 -94 4868 -42
rect -23 -2212 29 -236
rect 95 -2212 147 -236
rect 213 -2212 265 -236
rect 331 -2212 383 -236
rect 449 -2212 501 -236
rect 567 -2212 619 -236
rect 685 -2212 737 -236
rect 803 -2212 855 -236
rect 921 -2212 973 -236
rect 1039 -2212 1091 -236
rect 1157 -2212 1209 -236
rect 1420 -3580 1480 -2360
rect 1658 -3328 1710 -1352
rect 2116 -3328 2168 -1352
rect 2574 -3328 2626 -1352
rect 3032 -3328 3084 -1352
rect 3490 -3328 3542 -1352
rect 3990 -2212 4042 -236
rect 4108 -2212 4160 -236
rect 4226 -2212 4278 -236
rect 4344 -2212 4396 -236
rect 4462 -2212 4514 -236
rect 4580 -2212 4632 -236
rect 4698 -2212 4750 -236
rect 4816 -2212 4868 -236
rect 4934 -2212 4986 -236
rect 5052 -2212 5104 -236
rect 5170 -2212 5222 -236
rect 3720 -3580 3780 -2360
<< metal2 >>
rect 0 2600 5200 2800
rect 0 2500 100 2600
rect 400 2500 500 2600
rect 800 2500 900 2600
rect 1200 2500 1300 2600
rect 1600 2500 1700 2600
rect 2000 2500 2100 2600
rect 2400 2500 2500 2600
rect 2700 2500 2800 2600
rect 3100 2500 3200 2600
rect 3500 2500 3600 2600
rect 3900 2500 4000 2600
rect 4300 2500 4400 2600
rect 4700 2500 4800 2600
rect 5100 2500 5200 2600
rect 213 34 974 136
rect 213 -31 265 34
rect 449 -31 501 34
rect 685 -31 737 34
rect 921 -31 973 34
rect 213 -40 973 -31
rect 213 -96 329 -40
rect 385 -96 565 -40
rect 621 -96 801 -40
rect 857 -96 973 -40
rect 213 -105 973 -96
rect -23 -236 29 -224
rect -23 -2364 29 -2212
rect 95 -236 147 -224
rect 95 -2364 147 -2212
rect 213 -236 265 -105
rect 213 -2224 265 -2212
rect 331 -236 383 -224
rect 331 -2364 383 -2212
rect 449 -236 501 -105
rect 449 -2224 501 -2212
rect 567 -236 619 -224
rect 567 -2364 619 -2212
rect 685 -236 737 -105
rect 685 -2224 737 -2212
rect 803 -236 855 -224
rect 803 -2364 855 -2212
rect 921 -236 973 -105
rect 921 -2224 973 -2212
rect 1039 -236 1091 -224
rect 1039 -2340 1091 -2212
rect 1157 -236 1209 -224
rect 2220 -255 2324 105
rect 2876 102 2928 105
rect 2876 -255 2980 102
rect 4226 34 4986 136
rect 3990 -236 4042 -224
rect 1805 -1216 1859 -1057
rect 1997 -1216 2051 -1057
rect 2189 -1216 2243 -1057
rect 2381 -1216 2435 -1057
rect 2573 -1216 2627 -1057
rect 2765 -1216 2819 -1057
rect 2957 -1216 3011 -1057
rect 3149 -1216 3203 -1057
rect 3341 -1216 3395 -1057
rect 1805 -1308 3395 -1216
rect 1157 -2340 1209 -2212
rect 1658 -1352 1710 -1340
rect 1039 -2360 1500 -2340
rect 1039 -2364 1420 -2360
rect -23 -2434 1420 -2364
rect 0 -2600 100 -2434
rect 200 -2600 300 -2434
rect 400 -2600 500 -2434
rect 600 -2600 700 -2434
rect 800 -2600 900 -2434
rect 1000 -2440 1420 -2434
rect 1000 -2600 1100 -2440
rect 1200 -2600 1300 -2440
rect 1400 -2600 1420 -2440
rect 0 -2800 1420 -2600
rect 1100 -3100 1300 -2800
rect 1400 -3100 1420 -2800
rect 1100 -3200 1420 -3100
rect 1100 -3500 1300 -3200
rect 1400 -3500 1420 -3200
rect 1100 -3580 1420 -3500
rect 1480 -3500 1500 -2360
rect 1658 -3480 1710 -3328
rect 2116 -1352 2168 -1308
rect 2116 -3340 2168 -3328
rect 2574 -1352 2626 -1340
rect 2574 -3480 2626 -3328
rect 3032 -1352 3084 -1308
rect 3032 -3340 3084 -3328
rect 3490 -1352 3542 -1340
rect 3990 -2340 4042 -2212
rect 4108 -236 4160 -224
rect 4108 -2340 4160 -2212
rect 4226 -236 4278 34
rect 4339 -40 4400 -31
rect 4339 -96 4342 -40
rect 4398 -96 4400 -40
rect 4339 -105 4400 -96
rect 4226 -2224 4278 -2212
rect 4344 -236 4396 -224
rect 3490 -3480 3542 -3328
rect 1658 -3500 3542 -3480
rect 3700 -2360 4160 -2340
rect 3700 -3500 3720 -2360
rect 1480 -3580 3720 -3500
rect 3780 -2364 4160 -2360
rect 4344 -2364 4396 -2212
rect 4462 -236 4514 34
rect 4575 -40 4636 -31
rect 4575 -96 4578 -40
rect 4634 -96 4636 -40
rect 4575 -105 4636 -96
rect 4462 -2224 4514 -2212
rect 4580 -236 4632 -224
rect 4580 -2364 4632 -2212
rect 4698 -236 4750 34
rect 4811 -40 4872 -31
rect 4811 -96 4814 -40
rect 4870 -96 4872 -40
rect 4811 -105 4872 -96
rect 4698 -2224 4750 -2212
rect 4816 -236 4868 -224
rect 4816 -2364 4868 -2212
rect 4934 -236 4986 34
rect 4934 -2224 4986 -2212
rect 5052 -236 5104 -224
rect 5052 -2364 5104 -2212
rect 5170 -236 5222 -224
rect 5170 -2364 5222 -2212
rect 3780 -2434 5222 -2364
rect 3780 -2440 4200 -2434
rect 3780 -2700 3800 -2440
rect 3900 -2600 4000 -2440
rect 4100 -2600 4200 -2440
rect 4300 -2600 4400 -2434
rect 4500 -2600 4600 -2434
rect 4700 -2600 4800 -2434
rect 4900 -2600 5000 -2434
rect 5100 -2600 5200 -2434
rect 3900 -2700 5200 -2600
rect 3780 -2800 5200 -2700
rect 3780 -3100 3800 -2800
rect 3900 -3100 4100 -2800
rect 3780 -3200 4100 -3100
rect 3780 -3500 3800 -3200
rect 3900 -3500 4100 -3200
rect 3780 -3580 4100 -3500
rect 1100 -3800 4100 -3580
<< via2 >>
rect 329 -42 385 -40
rect 329 -94 331 -42
rect 331 -94 383 -42
rect 383 -94 385 -42
rect 329 -96 385 -94
rect 565 -42 621 -40
rect 565 -94 567 -42
rect 567 -94 619 -42
rect 619 -94 621 -42
rect 565 -96 621 -94
rect 801 -42 857 -40
rect 801 -94 803 -42
rect 803 -94 855 -42
rect 855 -94 857 -42
rect 801 -96 857 -94
rect 4342 -42 4398 -40
rect 4342 -94 4344 -42
rect 4344 -94 4396 -42
rect 4396 -94 4398 -42
rect 4342 -96 4398 -94
rect 4578 -42 4634 -40
rect 4578 -94 4580 -42
rect 4580 -94 4632 -42
rect 4632 -94 4634 -42
rect 4578 -96 4634 -94
rect 4814 -42 4870 -40
rect 4814 -94 4816 -42
rect 4816 -94 4868 -42
rect 4868 -94 4870 -42
rect 4814 -96 4870 -94
<< metal3 >>
rect 324 -40 4875 -31
rect 324 -96 329 -40
rect 385 -96 565 -40
rect 621 -96 801 -40
rect 857 -96 4342 -40
rect 4398 -96 4578 -40
rect 4634 -96 4814 -40
rect 4870 -96 4875 -40
rect 324 -105 4875 -96
rect 860 -136 4339 -105
rect 1900 -1010 1960 -950
rect 3240 -1010 3300 -950
<< comment >>
rect 2600 -1900 2603 2640
use imirror_pfb_1_8  imirror_pfb_1_8_0
timestamp 1671169241
transform 1 0 1275 0 1 -4606
box -1438 4640 4088 7142
use inputpair_0p15_2p5x8_lvt  inputpair_0p15_2p5x8_lvt_0
timestamp 1671154469
transform 1 0 9487 0 -1 4842
box -8014 5032 -5760 5972
use sky130_fd_pr__nfet_01v8_C44ETF  sky130_fd_pr__nfet_01v8_C44ETF_0
timestamp 1671166957
transform 1 0 4606 0 1 -1224
box -757 -1210 757 1210
use sky130_fd_pr__nfet_01v8_C44ETF  sky130_fd_pr__nfet_01v8_C44ETF_1
timestamp 1671166957
transform -1 0 593 0 1 -1224
box -757 -1210 757 1210
use sky130_fd_pr__nfet_01v8_CA7RJ6  sky130_fd_pr__nfet_01v8_CA7RJ6_0
timestamp 1671167000
transform 1 0 2600 0 1 -2340
box -1083 -1210 1083 1210
<< labels >>
rlabel metal2 0 2700 200 2800 1 VHI
rlabel metal2 1100 -3700 1300 -3600 1 VLO
rlabel metal3 1900 -1010 1960 -950 1 VIN
rlabel metal3 3240 -1010 3300 -950 1 VIP
rlabel metal2 4940 -10 4980 30 1 VOP
rlabel metal1 1672 -1308 1697 -1262 1 VREF
<< end >>
