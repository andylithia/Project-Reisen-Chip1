magic
tech sky130A
timestamp 1671388962
<< nwell >>
rect -1459 832 2467 1018
rect -1459 314 2467 500
rect -883 166 2467 314
<< pwell >>
rect -944 1776 -733 1841
rect -944 1749 -854 1776
rect -827 1749 -733 1776
rect -944 1419 -733 1749
rect -944 1392 -854 1419
rect -827 1392 -733 1419
rect -944 1074 -733 1392
rect -553 1776 -342 1841
rect -553 1749 -459 1776
rect -432 1749 -342 1776
rect -553 1419 -342 1749
rect -553 1392 -459 1419
rect -432 1392 -342 1419
rect -553 1074 -342 1392
rect -1402 690 -1297 790
rect -718 690 -581 790
rect -568 690 -259 763
rect 2 690 93 793
rect 104 690 412 763
rect 440 690 748 763
rect 776 690 1084 763
rect 1112 690 1420 763
rect 1448 690 1756 763
rect 1784 690 2092 763
rect 2120 690 2301 763
rect -1440 641 2448 690
rect -1402 542 -1297 641
rect -718 542 -581 641
rect -575 542 -145 641
rect -142 542 -1 641
rect 2 538 93 641
rect 99 570 1919 641
rect 99 557 1132 570
rect 99 551 1085 557
rect 427 548 1085 551
rect 427 530 609 548
rect 819 535 1085 548
rect 1269 542 1919 570
rect 1920 542 2015 641
rect 2016 542 2447 641
rect 1467 521 1561 542
rect -826 24 -721 124
rect -142 24 -5 124
rect 2 24 93 127
rect 427 117 609 136
rect 819 117 1085 130
rect 1467 124 1561 145
rect 427 114 1085 117
rect 99 109 1085 114
rect 99 96 1132 109
rect 1269 96 1919 124
rect 99 24 1919 96
rect 1920 24 2015 124
rect 2016 24 2447 136
rect -864 0 2448 24
rect -769 -109 -558 -44
rect -769 -135 -675 -109
rect -648 -135 -558 -109
rect -769 -466 -558 -135
rect -769 -492 -675 -466
rect -648 -492 -558 -466
rect -769 -811 -558 -492
<< nmos >>
rect -846 1536 -831 1736
rect -846 1179 -831 1379
rect -455 1536 -440 1736
rect -455 1179 -440 1379
rect -671 -349 -656 -149
rect -671 -706 -656 -506
<< scpmos >>
rect -1355 850 -1340 962
rect -678 850 -663 962
rect -633 850 -618 962
rect -535 862 -435 962
rect -407 862 -307 962
rect 137 862 237 962
rect 264 862 364 962
rect 473 862 573 962
rect 600 862 700 962
rect 809 862 909 962
rect 936 862 1036 962
rect 1145 862 1245 962
rect 1272 862 1372 962
rect 1481 862 1581 962
rect 1608 862 1708 962
rect 1817 862 1917 962
rect 1944 862 2044 962
rect 2153 862 2253 962
rect -1355 370 -1340 482
rect -678 370 -663 482
rect -633 370 -618 482
rect -533 398 -518 482
rect -479 382 -464 482
rect -383 382 -368 482
rect -329 382 -314 482
rect -272 382 -257 482
rect -210 370 -195 482
rect -102 370 -87 482
rect -57 370 -42 482
rect 139 370 154 434
rect 184 370 199 434
rect 223 370 238 434
rect 268 370 283 434
rect 369 370 384 434
rect 470 370 485 482
rect 515 370 530 482
rect 616 392 631 434
rect 658 392 673 434
rect 711 370 726 434
rect 877 370 892 454
rect 919 370 934 454
rect 973 370 988 454
rect 1074 370 1089 454
rect 1113 370 1128 454
rect 1166 370 1181 412
rect 1205 370 1220 412
rect 1308 370 1323 470
rect 1359 370 1374 470
rect 1401 370 1416 470
rect 1502 402 1517 466
rect 1620 370 1635 482
rect 1665 370 1680 482
rect 1764 374 1779 474
rect 1817 370 1832 482
rect 1862 370 1877 482
rect 2059 370 2074 482
rect 2185 370 2200 482
rect 2235 370 2250 482
rect 2385 370 2400 482
rect -779 184 -764 296
rect -102 184 -87 296
rect -57 184 -42 296
rect 139 232 154 296
rect 184 232 199 296
rect 223 232 238 296
rect 268 232 283 296
rect 369 232 384 296
rect 470 184 485 296
rect 515 184 530 296
rect 616 232 631 274
rect 658 232 673 274
rect 711 232 726 296
rect 877 212 892 296
rect 919 212 934 296
rect 973 212 988 296
rect 1074 212 1089 296
rect 1113 212 1128 296
rect 1166 254 1181 296
rect 1205 254 1220 296
rect 1308 196 1323 296
rect 1359 196 1374 296
rect 1401 196 1416 296
rect 1502 199 1517 263
rect 1620 184 1635 296
rect 1665 184 1680 296
rect 1764 192 1779 292
rect 1817 184 1832 296
rect 1862 184 1877 296
rect 2059 204 2074 288
rect 2104 204 2119 288
rect 2152 204 2167 288
rect 2199 204 2214 288
rect 2253 184 2268 296
rect 2300 184 2315 296
rect 2345 184 2360 296
rect 2390 184 2405 296
<< nmoslvt >>
rect -1354 703 -1339 777
rect -676 703 -661 777
rect -637 703 -622 777
rect -528 708 -428 750
rect -400 708 -300 750
rect 143 708 243 750
rect 271 708 371 750
rect 479 708 579 750
rect 607 708 707 750
rect 815 708 915 750
rect 943 708 1043 750
rect 1151 708 1251 750
rect 1279 708 1379 750
rect 1487 708 1587 750
rect 1615 708 1715 750
rect 1823 708 1923 750
rect 1951 708 2051 750
rect 2159 708 2259 750
rect -1354 555 -1339 629
rect -676 555 -661 629
rect -637 555 -622 629
rect -534 555 -519 610
rect -478 555 -463 629
rect -439 555 -424 629
rect -369 555 -354 629
rect -273 555 -258 629
rect -202 555 -187 629
rect -100 555 -85 629
rect -57 555 -42 629
rect 140 564 155 606
rect 179 564 194 606
rect 262 564 277 606
rect 301 564 316 606
rect 369 564 384 606
rect 468 543 483 617
rect 552 543 567 617
rect 673 561 688 603
rect 709 561 724 603
rect 755 561 770 603
rect 878 548 893 603
rect 921 548 936 603
rect 982 548 997 603
rect 1032 548 1047 603
rect 1079 570 1094 625
rect 1204 583 1219 625
rect 1243 583 1258 625
rect 1307 555 1322 629
rect 1359 555 1374 629
rect 1402 555 1417 629
rect 1508 534 1523 576
rect 1611 555 1626 629
rect 1654 555 1669 629
rect 1760 555 1775 619
rect 1820 555 1835 629
rect 1863 555 1878 629
rect 2058 555 2073 629
rect 2101 555 2116 629
rect 2144 555 2159 629
rect 2187 555 2202 629
rect 2234 555 2249 629
rect 2280 555 2295 629
rect 2330 555 2345 629
rect 2386 555 2401 629
rect -778 37 -763 111
rect -100 37 -85 111
rect -61 37 -46 111
rect 140 59 155 101
rect 179 59 194 101
rect 262 59 277 101
rect 301 59 316 101
rect 369 59 384 101
rect 468 49 483 123
rect 552 49 567 123
rect 673 62 688 104
rect 709 62 724 104
rect 755 62 770 104
rect 878 62 893 117
rect 921 62 936 117
rect 982 62 997 117
rect 1032 62 1047 117
rect 1079 41 1094 96
rect 1204 41 1219 83
rect 1243 41 1258 83
rect 1307 37 1322 111
rect 1359 37 1374 111
rect 1402 37 1417 111
rect 1508 90 1523 132
rect 1611 37 1626 111
rect 1654 37 1669 111
rect 1760 47 1775 111
rect 1820 37 1835 111
rect 1863 37 1878 111
rect 2058 59 2073 123
rect 2103 59 2118 123
rect 2150 59 2165 123
rect 2196 59 2211 123
rect 2247 49 2262 123
rect 2305 49 2320 123
rect 2348 49 2363 123
rect 2391 49 2406 123
<< ndiff >>
rect -875 1730 -846 1736
rect -875 1542 -869 1730
rect -852 1542 -846 1730
rect -875 1536 -846 1542
rect -831 1730 -802 1736
rect -831 1542 -825 1730
rect -808 1542 -802 1730
rect -831 1536 -802 1542
rect -875 1373 -846 1379
rect -875 1185 -869 1373
rect -852 1185 -846 1373
rect -875 1179 -846 1185
rect -831 1373 -802 1379
rect -831 1185 -825 1373
rect -808 1185 -802 1373
rect -831 1179 -802 1185
rect -484 1730 -455 1736
rect -484 1542 -478 1730
rect -461 1542 -455 1730
rect -484 1536 -455 1542
rect -440 1730 -411 1736
rect -440 1542 -434 1730
rect -417 1542 -411 1730
rect -440 1536 -411 1542
rect -484 1373 -455 1379
rect -484 1185 -478 1373
rect -461 1185 -455 1373
rect -484 1179 -455 1185
rect -440 1373 -411 1379
rect -440 1185 -434 1373
rect -417 1185 -411 1373
rect -440 1179 -411 1185
rect -1389 771 -1354 777
rect -1389 754 -1383 771
rect -1366 754 -1354 771
rect -1389 726 -1354 754
rect -1389 709 -1383 726
rect -1366 709 -1354 726
rect -1389 703 -1354 709
rect -1339 771 -1310 777
rect -1339 754 -1333 771
rect -1316 754 -1310 771
rect -1339 726 -1310 754
rect -705 767 -676 777
rect -705 750 -699 767
rect -682 750 -676 767
rect -1339 709 -1333 726
rect -1316 709 -1310 726
rect -1339 703 -1310 709
rect -705 726 -676 750
rect -705 709 -699 726
rect -682 709 -676 726
rect -705 703 -676 709
rect -661 703 -637 777
rect -622 767 -594 777
rect -622 750 -617 767
rect -600 750 -594 767
rect -622 726 -594 750
rect -622 709 -617 726
rect -600 709 -594 726
rect -622 703 -594 709
rect -555 738 -528 750
rect -555 721 -551 738
rect -534 721 -528 738
rect -555 708 -528 721
rect -428 738 -400 750
rect -428 721 -423 738
rect -406 721 -400 738
rect -428 708 -400 721
rect -300 738 -272 750
rect -300 721 -295 738
rect -278 721 -272 738
rect -300 708 -272 721
rect 117 738 143 750
rect 117 721 121 738
rect 138 721 143 738
rect 117 708 143 721
rect 243 738 271 750
rect 243 721 249 738
rect 266 721 271 738
rect 243 708 271 721
rect 371 738 399 750
rect 371 721 377 738
rect 394 721 399 738
rect 371 708 399 721
rect 453 738 479 750
rect 453 721 457 738
rect 474 721 479 738
rect 453 708 479 721
rect 579 738 607 750
rect 579 721 585 738
rect 602 721 607 738
rect 579 708 607 721
rect 707 738 735 750
rect 707 721 713 738
rect 730 721 735 738
rect 707 708 735 721
rect 789 738 815 750
rect 789 721 793 738
rect 810 721 815 738
rect 789 708 815 721
rect 915 738 943 750
rect 915 721 921 738
rect 938 721 943 738
rect 915 708 943 721
rect 1043 738 1071 750
rect 1043 721 1049 738
rect 1066 721 1071 738
rect 1043 708 1071 721
rect 1125 738 1151 750
rect 1125 721 1129 738
rect 1146 721 1151 738
rect 1125 708 1151 721
rect 1251 738 1279 750
rect 1251 721 1257 738
rect 1274 721 1279 738
rect 1251 708 1279 721
rect 1379 738 1407 750
rect 1379 721 1385 738
rect 1402 721 1407 738
rect 1379 708 1407 721
rect 1461 738 1487 750
rect 1461 721 1465 738
rect 1482 721 1487 738
rect 1461 708 1487 721
rect 1587 738 1615 750
rect 1587 721 1593 738
rect 1610 721 1615 738
rect 1587 708 1615 721
rect 1715 738 1743 750
rect 1715 721 1721 738
rect 1738 721 1743 738
rect 1715 708 1743 721
rect 1797 738 1823 750
rect 1797 721 1801 738
rect 1818 721 1823 738
rect 1797 708 1823 721
rect 1923 738 1951 750
rect 1923 721 1929 738
rect 1946 721 1951 738
rect 1923 708 1951 721
rect 2051 738 2079 750
rect 2051 721 2057 738
rect 2074 721 2079 738
rect 2051 708 2079 721
rect 2133 738 2159 750
rect 2133 721 2137 738
rect 2154 721 2159 738
rect 2133 708 2159 721
rect 2259 738 2288 750
rect 2259 721 2265 738
rect 2282 721 2288 738
rect 2259 708 2288 721
rect -1389 623 -1354 629
rect -1389 606 -1383 623
rect -1366 606 -1354 623
rect -1389 578 -1354 606
rect -1389 561 -1383 578
rect -1366 561 -1354 578
rect -1389 555 -1354 561
rect -1339 623 -1310 629
rect -1339 606 -1333 623
rect -1316 606 -1310 623
rect -1339 578 -1310 606
rect -705 623 -676 629
rect -705 606 -699 623
rect -682 606 -676 623
rect -1339 561 -1333 578
rect -1316 561 -1310 578
rect -1339 555 -1310 561
rect -705 582 -676 606
rect -705 565 -699 582
rect -682 565 -676 582
rect -705 555 -676 565
rect -661 555 -637 629
rect -622 623 -594 629
rect -511 623 -478 629
rect -622 606 -617 623
rect -600 606 -594 623
rect -511 610 -503 623
rect -622 582 -594 606
rect -622 565 -617 582
rect -600 565 -594 582
rect -622 555 -594 565
rect -562 591 -534 610
rect -562 574 -556 591
rect -539 574 -534 591
rect -562 555 -534 574
rect -519 606 -503 610
rect -486 606 -478 623
rect -519 578 -478 606
rect -519 561 -512 578
rect -495 561 -478 578
rect -519 555 -478 561
rect -463 555 -439 629
rect -424 619 -369 629
rect -424 602 -405 619
rect -388 602 -369 619
rect -424 555 -369 602
rect -354 555 -273 629
rect -258 610 -202 629
rect -258 593 -238 610
rect -221 593 -202 610
rect -258 555 -202 593
rect -187 623 -158 629
rect -187 606 -181 623
rect -164 606 -158 623
rect -187 578 -158 606
rect -187 561 -181 578
rect -164 561 -158 578
rect -187 555 -158 561
rect -129 623 -100 629
rect -129 606 -123 623
rect -106 606 -100 623
rect -129 578 -100 606
rect -129 561 -123 578
rect -106 561 -100 578
rect -129 555 -100 561
rect -85 623 -57 629
rect -85 606 -80 623
rect -63 606 -57 623
rect -85 578 -57 606
rect -85 561 -80 578
rect -63 561 -57 578
rect -85 555 -57 561
rect -42 623 -14 629
rect -42 606 -37 623
rect -20 606 -14 623
rect -42 578 -14 606
rect -42 561 -37 578
rect -20 561 -14 578
rect -42 555 -14 561
rect 491 642 520 648
rect 491 625 497 642
rect 514 625 520 642
rect 491 617 520 625
rect 635 624 666 630
rect 112 598 140 606
rect 112 581 118 598
rect 135 581 140 598
rect 112 564 140 581
rect 155 564 179 606
rect 194 595 262 606
rect 194 578 200 595
rect 217 578 240 595
rect 257 578 262 595
rect 194 564 262 578
rect 277 564 301 606
rect 316 598 369 606
rect 316 581 322 598
rect 339 581 369 598
rect 316 564 369 581
rect 384 593 413 606
rect 384 576 390 593
rect 407 576 413 593
rect 384 564 413 576
rect 440 566 468 617
rect 440 549 446 566
rect 463 549 468 566
rect 440 543 468 549
rect 483 543 552 617
rect 567 598 596 617
rect 567 581 573 598
rect 590 581 596 598
rect 567 564 596 581
rect 567 547 573 564
rect 590 547 596 564
rect 635 607 642 624
rect 659 607 666 624
rect 635 603 666 607
rect 832 623 871 629
rect 1266 640 1299 646
rect 1266 625 1274 640
rect 832 606 843 623
rect 860 606 871 623
rect 832 603 871 606
rect 1054 603 1079 625
rect 635 561 673 603
rect 688 561 709 603
rect 724 591 755 603
rect 724 574 732 591
rect 749 574 755 591
rect 724 561 755 574
rect 770 593 805 603
rect 770 576 782 593
rect 799 576 805 593
rect 770 561 805 576
rect 567 543 596 547
rect 832 548 878 603
rect 893 588 921 603
rect 893 571 899 588
rect 916 571 921 588
rect 893 548 921 571
rect 936 597 982 603
rect 936 580 954 597
rect 971 580 982 597
rect 936 548 982 580
rect 997 597 1032 603
rect 997 580 1009 597
rect 1026 580 1032 597
rect 997 548 1032 580
rect 1047 570 1079 603
rect 1094 606 1204 625
rect 1094 589 1100 606
rect 1117 589 1141 606
rect 1158 589 1182 606
rect 1199 589 1204 606
rect 1094 583 1204 589
rect 1219 583 1243 625
rect 1258 623 1274 625
rect 1291 629 1299 640
rect 1424 633 1453 639
rect 1424 629 1430 633
rect 1291 623 1307 629
rect 1258 583 1307 623
rect 1094 570 1119 583
rect 1047 548 1072 570
rect 1282 555 1307 583
rect 1322 623 1359 629
rect 1322 606 1332 623
rect 1349 606 1359 623
rect 1322 555 1359 606
rect 1374 597 1402 629
rect 1374 580 1379 597
rect 1396 580 1402 597
rect 1374 555 1402 580
rect 1417 616 1430 629
rect 1447 616 1453 633
rect 1417 555 1453 616
rect 1585 623 1611 629
rect 1585 606 1589 623
rect 1606 606 1611 623
rect 1585 578 1611 606
rect 1585 576 1589 578
rect 1480 557 1508 576
rect 1480 540 1486 557
rect 1503 540 1508 557
rect 1480 534 1508 540
rect 1523 561 1589 576
rect 1606 561 1611 578
rect 1523 555 1611 561
rect 1626 623 1654 629
rect 1626 606 1632 623
rect 1649 606 1654 623
rect 1626 578 1654 606
rect 1626 561 1632 578
rect 1649 561 1654 578
rect 1626 555 1654 561
rect 1669 623 1700 629
rect 1669 606 1675 623
rect 1692 606 1700 623
rect 1785 623 1820 629
rect 1785 619 1791 623
rect 1669 578 1700 606
rect 1669 561 1675 578
rect 1692 561 1700 578
rect 1669 555 1700 561
rect 1732 610 1760 619
rect 1732 593 1738 610
rect 1755 593 1760 610
rect 1732 576 1760 593
rect 1732 559 1738 576
rect 1755 559 1760 576
rect 1732 555 1760 559
rect 1775 606 1791 619
rect 1808 606 1820 623
rect 1775 586 1820 606
rect 1775 569 1791 586
rect 1808 569 1820 586
rect 1775 555 1820 569
rect 1835 623 1863 629
rect 1835 606 1841 623
rect 1858 606 1863 623
rect 1835 586 1863 606
rect 1835 569 1841 586
rect 1858 569 1863 586
rect 1835 555 1863 569
rect 1878 623 1906 629
rect 1878 606 1884 623
rect 1901 606 1906 623
rect 1878 578 1906 606
rect 1878 561 1884 578
rect 1901 561 1906 578
rect 1878 555 1906 561
rect 1933 625 2002 629
rect 1933 608 1941 625
rect 1958 608 1977 625
rect 1994 608 2002 625
rect 1933 555 2002 608
rect 2029 623 2058 629
rect 2029 606 2035 623
rect 2052 606 2058 623
rect 2029 578 2058 606
rect 2029 561 2035 578
rect 2052 561 2058 578
rect 2029 555 2058 561
rect 2073 612 2101 629
rect 2073 595 2078 612
rect 2095 595 2101 612
rect 2073 555 2101 595
rect 2116 623 2144 629
rect 2116 606 2121 623
rect 2138 606 2144 623
rect 2116 578 2144 606
rect 2116 561 2121 578
rect 2138 561 2144 578
rect 2116 555 2144 561
rect 2159 612 2187 629
rect 2159 595 2164 612
rect 2181 595 2187 612
rect 2159 555 2187 595
rect 2202 623 2234 629
rect 2202 606 2207 623
rect 2224 606 2234 623
rect 2202 578 2234 606
rect 2202 561 2207 578
rect 2224 561 2234 578
rect 2202 555 2234 561
rect 2249 596 2280 629
rect 2249 579 2257 596
rect 2274 579 2280 596
rect 2249 555 2280 579
rect 2295 612 2330 629
rect 2295 595 2307 612
rect 2324 595 2330 612
rect 2295 555 2330 595
rect 2345 596 2386 629
rect 2345 579 2359 596
rect 2376 579 2386 596
rect 2345 555 2386 579
rect 2401 612 2434 629
rect 2401 595 2411 612
rect 2428 595 2434 612
rect 2401 555 2434 595
rect 1523 534 1548 555
rect -813 105 -778 111
rect -813 88 -807 105
rect -790 88 -778 105
rect -813 60 -778 88
rect -813 43 -807 60
rect -790 43 -778 60
rect -813 37 -778 43
rect -763 105 -734 111
rect -763 88 -757 105
rect -740 88 -734 105
rect -763 60 -734 88
rect -129 101 -100 111
rect -129 84 -123 101
rect -106 84 -100 101
rect -763 43 -757 60
rect -740 43 -734 60
rect -763 37 -734 43
rect -129 60 -100 84
rect -129 43 -123 60
rect -106 43 -100 60
rect -129 37 -100 43
rect -85 37 -61 111
rect -46 101 -18 111
rect -46 84 -41 101
rect -24 84 -18 101
rect -46 60 -18 84
rect -46 43 -41 60
rect -24 43 -18 60
rect -46 37 -18 43
rect 440 117 468 123
rect 112 85 140 101
rect 112 68 118 85
rect 135 68 140 85
rect 112 59 140 68
rect 155 59 179 101
rect 194 87 262 101
rect 194 70 200 87
rect 217 70 240 87
rect 257 70 262 87
rect 194 59 262 70
rect 277 59 301 101
rect 316 84 369 101
rect 316 67 322 84
rect 339 67 369 84
rect 316 59 369 67
rect 384 90 413 101
rect 384 73 390 90
rect 407 73 413 90
rect 384 59 413 73
rect 440 100 446 117
rect 463 100 468 117
rect 440 49 468 100
rect 483 49 552 123
rect 567 118 596 123
rect 567 101 573 118
rect 590 101 596 118
rect 567 84 596 101
rect 567 67 573 84
rect 590 67 596 84
rect 567 49 596 67
rect 635 62 673 104
rect 688 62 709 104
rect 724 92 755 104
rect 724 75 732 92
rect 749 75 755 92
rect 724 62 755 75
rect 770 89 805 104
rect 770 72 782 89
rect 799 72 805 89
rect 770 62 805 72
rect 832 62 878 117
rect 893 94 921 117
rect 893 77 899 94
rect 916 77 921 94
rect 893 62 921 77
rect 936 85 982 117
rect 936 68 954 85
rect 971 68 982 85
rect 936 62 982 68
rect 997 85 1032 117
rect 997 68 1009 85
rect 1026 68 1032 85
rect 997 62 1032 68
rect 1047 96 1072 117
rect 1047 62 1079 96
rect 635 59 666 62
rect 491 41 520 49
rect 491 24 497 41
rect 514 24 520 41
rect 491 18 520 24
rect 635 42 642 59
rect 659 42 666 59
rect 635 36 666 42
rect 832 59 871 62
rect 832 42 843 59
rect 860 42 871 59
rect 832 36 871 42
rect 1054 41 1079 62
rect 1094 83 1119 96
rect 1480 125 1508 132
rect 1282 83 1307 111
rect 1094 77 1204 83
rect 1094 60 1100 77
rect 1117 60 1141 77
rect 1158 60 1182 77
rect 1199 60 1204 77
rect 1094 41 1204 60
rect 1219 41 1243 83
rect 1258 43 1307 83
rect 1258 41 1274 43
rect 1266 26 1274 41
rect 1291 37 1307 43
rect 1322 60 1359 111
rect 1322 43 1332 60
rect 1349 43 1359 60
rect 1322 37 1359 43
rect 1374 86 1402 111
rect 1374 69 1379 86
rect 1396 69 1402 86
rect 1374 37 1402 69
rect 1417 49 1453 111
rect 1480 108 1486 125
rect 1503 108 1508 125
rect 1480 90 1508 108
rect 1523 111 1548 132
rect 2029 117 2058 123
rect 1523 105 1611 111
rect 1523 90 1589 105
rect 1585 88 1589 90
rect 1606 88 1611 105
rect 1417 37 1430 49
rect 1291 26 1299 37
rect 1266 20 1299 26
rect 1424 32 1430 37
rect 1447 32 1453 49
rect 1585 60 1611 88
rect 1585 43 1589 60
rect 1606 43 1611 60
rect 1585 37 1611 43
rect 1626 105 1654 111
rect 1626 88 1632 105
rect 1649 88 1654 105
rect 1626 60 1654 88
rect 1626 43 1632 60
rect 1649 43 1654 60
rect 1626 37 1654 43
rect 1669 105 1700 111
rect 1669 88 1675 105
rect 1692 88 1700 105
rect 1669 60 1700 88
rect 1669 43 1675 60
rect 1692 43 1700 60
rect 1732 107 1760 111
rect 1732 90 1738 107
rect 1755 90 1760 107
rect 1732 73 1760 90
rect 1732 56 1738 73
rect 1755 56 1760 73
rect 1732 47 1760 56
rect 1775 97 1820 111
rect 1775 80 1791 97
rect 1808 80 1820 97
rect 1775 60 1820 80
rect 1775 47 1791 60
rect 1669 37 1700 43
rect 1424 26 1453 32
rect 1785 43 1791 47
rect 1808 43 1820 60
rect 1785 37 1820 43
rect 1835 97 1863 111
rect 1835 80 1841 97
rect 1858 80 1863 97
rect 1835 60 1863 80
rect 1835 43 1841 60
rect 1858 43 1863 60
rect 1835 37 1863 43
rect 1878 105 1906 111
rect 1878 88 1884 105
rect 1901 88 1906 105
rect 1878 60 1906 88
rect 1878 43 1884 60
rect 1901 43 1906 60
rect 1878 37 1906 43
rect 1933 58 2002 111
rect 2029 100 2035 117
rect 2052 100 2058 117
rect 2029 82 2058 100
rect 2029 65 2035 82
rect 2052 65 2058 82
rect 2029 59 2058 65
rect 2073 84 2103 123
rect 2073 67 2080 84
rect 2097 67 2103 84
rect 2073 59 2103 67
rect 2118 119 2150 123
rect 2118 102 2123 119
rect 2140 102 2150 119
rect 2118 80 2150 102
rect 2118 63 2123 80
rect 2140 63 2150 80
rect 2118 59 2150 63
rect 2165 114 2196 123
rect 2165 97 2173 114
rect 2190 97 2196 114
rect 2165 80 2196 97
rect 2165 63 2173 80
rect 2190 63 2196 80
rect 2165 59 2196 63
rect 2211 117 2247 123
rect 2211 100 2224 117
rect 2241 100 2247 117
rect 2211 78 2247 100
rect 2211 61 2224 78
rect 2241 61 2247 78
rect 2211 59 2247 61
rect 1933 41 1941 58
rect 1958 41 1977 58
rect 1994 41 2002 58
rect 1933 37 2002 41
rect 2218 49 2247 59
rect 2262 109 2305 123
rect 2262 92 2275 109
rect 2292 92 2305 109
rect 2262 72 2305 92
rect 2262 55 2275 72
rect 2292 55 2305 72
rect 2262 49 2305 55
rect 2320 75 2348 123
rect 2320 58 2325 75
rect 2342 58 2348 75
rect 2320 49 2348 58
rect 2363 117 2391 123
rect 2363 100 2368 117
rect 2385 100 2391 117
rect 2363 72 2391 100
rect 2363 55 2368 72
rect 2385 55 2391 72
rect 2363 49 2391 55
rect 2406 117 2434 123
rect 2406 100 2411 117
rect 2428 100 2434 117
rect 2406 72 2434 100
rect 2406 55 2411 72
rect 2428 55 2434 72
rect 2406 49 2434 55
rect -700 -155 -671 -149
rect -700 -343 -694 -155
rect -677 -343 -671 -155
rect -700 -349 -671 -343
rect -656 -155 -627 -149
rect -656 -343 -650 -155
rect -633 -343 -627 -155
rect -656 -349 -627 -343
rect -700 -512 -671 -506
rect -700 -700 -694 -512
rect -677 -700 -671 -512
rect -700 -706 -671 -700
rect -656 -512 -627 -506
rect -656 -700 -650 -512
rect -633 -700 -627 -512
rect -656 -706 -627 -700
<< pdiff >>
rect -1389 956 -1355 962
rect -1389 939 -1383 956
rect -1366 939 -1355 956
rect -1389 921 -1355 939
rect -1389 904 -1383 921
rect -1366 904 -1355 921
rect -1389 886 -1355 904
rect -1389 869 -1383 886
rect -1366 869 -1355 886
rect -1389 850 -1355 869
rect -1340 956 -1310 962
rect -1340 939 -1333 956
rect -1316 939 -1310 956
rect -1340 914 -1310 939
rect -1340 897 -1333 914
rect -1316 897 -1310 914
rect -1340 873 -1310 897
rect -706 956 -678 962
rect -706 939 -701 956
rect -684 939 -678 956
rect -706 914 -678 939
rect -706 897 -701 914
rect -684 897 -678 914
rect -1340 856 -1333 873
rect -1316 856 -1310 873
rect -1340 850 -1310 856
rect -706 873 -678 897
rect -706 856 -701 873
rect -684 856 -678 873
rect -706 850 -678 856
rect -663 956 -633 962
rect -663 939 -656 956
rect -639 939 -633 956
rect -663 914 -633 939
rect -663 897 -656 914
rect -639 897 -633 914
rect -663 873 -633 897
rect -663 856 -656 873
rect -639 856 -633 873
rect -663 850 -633 856
rect -618 956 -589 962
rect -618 939 -611 956
rect -594 939 -589 956
rect -618 914 -589 939
rect -618 897 -611 914
rect -594 897 -589 914
rect -618 873 -589 897
rect -618 856 -611 873
rect -594 856 -589 873
rect -562 956 -535 962
rect -562 939 -558 956
rect -541 939 -535 956
rect -562 920 -535 939
rect -562 903 -558 920
rect -541 903 -535 920
rect -562 885 -535 903
rect -562 868 -558 885
rect -541 868 -535 885
rect -562 862 -535 868
rect -435 956 -407 962
rect -435 939 -429 956
rect -412 939 -407 956
rect -435 920 -407 939
rect -435 903 -429 920
rect -412 903 -407 920
rect -435 885 -407 903
rect -435 868 -429 885
rect -412 868 -407 885
rect -435 862 -407 868
rect -307 956 -279 962
rect -307 939 -302 956
rect -285 939 -279 956
rect -307 920 -279 939
rect -307 903 -302 920
rect -285 903 -279 920
rect -307 885 -279 903
rect -307 868 -302 885
rect -285 868 -279 885
rect 109 956 137 962
rect 109 939 113 956
rect 130 939 137 956
rect 109 920 137 939
rect 109 903 113 920
rect 130 903 137 920
rect 109 885 137 903
rect -307 862 -279 868
rect 109 868 113 885
rect 130 868 137 885
rect 109 862 137 868
rect 237 956 264 962
rect 237 939 242 956
rect 259 939 264 956
rect 237 920 264 939
rect 237 903 242 920
rect 259 903 264 920
rect 237 885 264 903
rect 237 868 242 885
rect 259 868 264 885
rect 237 862 264 868
rect 364 956 393 962
rect 364 939 370 956
rect 387 939 393 956
rect 364 920 393 939
rect 364 903 370 920
rect 387 903 393 920
rect 364 885 393 903
rect 364 868 370 885
rect 387 868 393 885
rect 364 862 393 868
rect 445 956 473 962
rect 445 939 449 956
rect 466 939 473 956
rect 445 920 473 939
rect 445 903 449 920
rect 466 903 473 920
rect 445 885 473 903
rect 445 868 449 885
rect 466 868 473 885
rect 445 862 473 868
rect 573 956 600 962
rect 573 939 578 956
rect 595 939 600 956
rect 573 920 600 939
rect 573 903 578 920
rect 595 903 600 920
rect 573 885 600 903
rect 573 868 578 885
rect 595 868 600 885
rect 573 862 600 868
rect 700 956 729 962
rect 700 939 706 956
rect 723 939 729 956
rect 700 920 729 939
rect 700 903 706 920
rect 723 903 729 920
rect 700 885 729 903
rect 700 868 706 885
rect 723 868 729 885
rect 700 862 729 868
rect 781 956 809 962
rect 781 939 785 956
rect 802 939 809 956
rect 781 920 809 939
rect 781 903 785 920
rect 802 903 809 920
rect 781 885 809 903
rect 781 868 785 885
rect 802 868 809 885
rect 781 862 809 868
rect 909 956 936 962
rect 909 939 914 956
rect 931 939 936 956
rect 909 920 936 939
rect 909 903 914 920
rect 931 903 936 920
rect 909 885 936 903
rect 909 868 914 885
rect 931 868 936 885
rect 909 862 936 868
rect 1036 956 1065 962
rect 1036 939 1042 956
rect 1059 939 1065 956
rect 1036 920 1065 939
rect 1036 903 1042 920
rect 1059 903 1065 920
rect 1036 885 1065 903
rect 1036 868 1042 885
rect 1059 868 1065 885
rect 1036 862 1065 868
rect 1117 956 1145 962
rect 1117 939 1121 956
rect 1138 939 1145 956
rect 1117 920 1145 939
rect 1117 903 1121 920
rect 1138 903 1145 920
rect 1117 885 1145 903
rect 1117 868 1121 885
rect 1138 868 1145 885
rect 1117 862 1145 868
rect 1245 956 1272 962
rect 1245 939 1250 956
rect 1267 939 1272 956
rect 1245 920 1272 939
rect 1245 903 1250 920
rect 1267 903 1272 920
rect 1245 885 1272 903
rect 1245 868 1250 885
rect 1267 868 1272 885
rect 1245 862 1272 868
rect 1372 956 1401 962
rect 1372 939 1378 956
rect 1395 939 1401 956
rect 1372 920 1401 939
rect 1372 903 1378 920
rect 1395 903 1401 920
rect 1372 885 1401 903
rect 1372 868 1378 885
rect 1395 868 1401 885
rect 1372 862 1401 868
rect 1453 956 1481 962
rect 1453 939 1457 956
rect 1474 939 1481 956
rect 1453 920 1481 939
rect 1453 903 1457 920
rect 1474 903 1481 920
rect 1453 885 1481 903
rect 1453 868 1457 885
rect 1474 868 1481 885
rect 1453 862 1481 868
rect 1581 956 1608 962
rect 1581 939 1586 956
rect 1603 939 1608 956
rect 1581 920 1608 939
rect 1581 903 1586 920
rect 1603 903 1608 920
rect 1581 885 1608 903
rect 1581 868 1586 885
rect 1603 868 1608 885
rect 1581 862 1608 868
rect 1708 956 1737 962
rect 1708 939 1714 956
rect 1731 939 1737 956
rect 1708 920 1737 939
rect 1708 903 1714 920
rect 1731 903 1737 920
rect 1708 885 1737 903
rect 1708 868 1714 885
rect 1731 868 1737 885
rect 1708 862 1737 868
rect 1789 956 1817 962
rect 1789 939 1793 956
rect 1810 939 1817 956
rect 1789 920 1817 939
rect 1789 903 1793 920
rect 1810 903 1817 920
rect 1789 885 1817 903
rect 1789 868 1793 885
rect 1810 868 1817 885
rect 1789 862 1817 868
rect 1917 956 1944 962
rect 1917 939 1922 956
rect 1939 939 1944 956
rect 1917 920 1944 939
rect 1917 903 1922 920
rect 1939 903 1944 920
rect 1917 885 1944 903
rect 1917 868 1922 885
rect 1939 868 1944 885
rect 1917 862 1944 868
rect 2044 956 2073 962
rect 2044 939 2050 956
rect 2067 939 2073 956
rect 2044 920 2073 939
rect 2044 903 2050 920
rect 2067 903 2073 920
rect 2044 885 2073 903
rect 2044 868 2050 885
rect 2067 868 2073 885
rect 2044 862 2073 868
rect 2125 956 2153 962
rect 2125 939 2129 956
rect 2146 939 2153 956
rect 2125 920 2153 939
rect 2125 903 2129 920
rect 2146 903 2153 920
rect 2125 885 2153 903
rect 2125 868 2129 885
rect 2146 868 2153 885
rect 2125 862 2153 868
rect 2253 956 2281 962
rect 2253 939 2258 956
rect 2275 939 2281 956
rect 2253 920 2281 939
rect 2253 903 2258 920
rect 2275 903 2281 920
rect 2253 885 2281 903
rect 2253 868 2258 885
rect 2275 868 2281 885
rect 2253 862 2281 868
rect -618 850 -589 856
rect -1389 463 -1355 482
rect -1389 446 -1383 463
rect -1366 446 -1355 463
rect -1389 428 -1355 446
rect -1389 411 -1383 428
rect -1366 411 -1355 428
rect -1389 393 -1355 411
rect -1389 376 -1383 393
rect -1366 376 -1355 393
rect -1389 370 -1355 376
rect -1340 476 -1310 482
rect -1340 459 -1333 476
rect -1316 459 -1310 476
rect -1340 434 -1310 459
rect -706 476 -678 482
rect -706 459 -701 476
rect -684 459 -678 476
rect -1340 417 -1333 434
rect -1316 417 -1310 434
rect -1340 393 -1310 417
rect -1340 376 -1333 393
rect -1316 376 -1310 393
rect -1340 370 -1310 376
rect -706 434 -678 459
rect -706 417 -701 434
rect -684 417 -678 434
rect -706 393 -678 417
rect -706 376 -701 393
rect -684 376 -678 393
rect -706 370 -678 376
rect -663 476 -633 482
rect -663 459 -656 476
rect -639 459 -633 476
rect -663 434 -633 459
rect -663 417 -656 434
rect -639 417 -633 434
rect -663 393 -633 417
rect -663 376 -656 393
rect -639 376 -633 393
rect -663 370 -633 376
rect -618 476 -589 482
rect -618 459 -611 476
rect -594 459 -589 476
rect -618 434 -589 459
rect -618 417 -611 434
rect -594 417 -589 434
rect -618 393 -589 417
rect -562 468 -533 482
rect -562 451 -556 468
rect -539 451 -533 468
rect -562 421 -533 451
rect -562 404 -556 421
rect -539 404 -533 421
rect -562 398 -533 404
rect -518 423 -479 482
rect -518 406 -503 423
rect -486 406 -479 423
rect -518 398 -479 406
rect -618 376 -611 393
rect -594 376 -589 393
rect -509 382 -479 398
rect -464 382 -383 482
rect -368 476 -329 482
rect -368 459 -361 476
rect -344 459 -329 476
rect -368 417 -329 459
rect -368 400 -361 417
rect -344 400 -329 417
rect -368 382 -329 400
rect -314 382 -272 482
rect -257 476 -210 482
rect -257 459 -238 476
rect -221 459 -210 476
rect -257 434 -210 459
rect -257 417 -238 434
rect -221 417 -210 434
rect -257 393 -210 417
rect -257 382 -238 393
rect -618 370 -589 376
rect -244 376 -238 382
rect -221 376 -210 393
rect -244 370 -210 376
rect -195 476 -165 482
rect -195 459 -188 476
rect -171 459 -165 476
rect -195 434 -165 459
rect -195 417 -188 434
rect -171 417 -165 434
rect -195 393 -165 417
rect -195 376 -188 393
rect -171 376 -165 393
rect -195 370 -165 376
rect -130 463 -102 482
rect -130 446 -125 463
rect -108 446 -102 463
rect -130 428 -102 446
rect -130 411 -125 428
rect -108 411 -102 428
rect -130 393 -102 411
rect -130 376 -125 393
rect -108 376 -102 393
rect -130 370 -102 376
rect -87 476 -57 482
rect -87 459 -80 476
rect -63 459 -57 476
rect -87 434 -57 459
rect -87 417 -80 434
rect -63 417 -57 434
rect -87 393 -57 417
rect -87 376 -80 393
rect -63 376 -57 393
rect -87 370 -57 376
rect -42 476 -13 482
rect -42 459 -35 476
rect -18 459 -13 476
rect -42 434 -13 459
rect -42 417 -35 434
rect -18 417 -13 434
rect -42 393 -13 417
rect -42 376 -35 393
rect -18 376 -13 393
rect -42 370 -13 376
rect 440 463 470 482
rect 440 446 446 463
rect 463 446 470 463
rect 109 427 139 434
rect 109 410 115 427
rect 132 410 139 427
rect 109 393 139 410
rect 109 376 115 393
rect 132 376 139 393
rect 109 370 139 376
rect 154 393 184 434
rect 154 376 160 393
rect 177 376 184 393
rect 154 370 184 376
rect 199 370 223 434
rect 238 423 268 434
rect 238 406 244 423
rect 261 406 268 423
rect 238 370 268 406
rect 283 428 312 434
rect 283 411 289 428
rect 306 411 312 428
rect 283 393 312 411
rect 283 376 289 393
rect 306 376 312 393
rect 283 370 312 376
rect 339 428 369 434
rect 339 411 345 428
rect 362 411 369 428
rect 339 393 369 411
rect 339 376 345 393
rect 362 376 369 393
rect 339 370 369 376
rect 384 428 413 434
rect 384 411 390 428
rect 407 411 413 428
rect 384 393 413 411
rect 384 376 390 393
rect 407 376 413 393
rect 384 370 413 376
rect 440 428 470 446
rect 440 411 446 428
rect 463 411 470 428
rect 440 393 470 411
rect 440 376 446 393
rect 463 376 470 393
rect 440 370 470 376
rect 485 432 515 482
rect 485 415 491 432
rect 508 415 515 432
rect 485 393 515 415
rect 485 376 491 393
rect 508 376 515 393
rect 485 370 515 376
rect 530 474 559 482
rect 530 457 536 474
rect 553 457 559 474
rect 530 433 559 457
rect 530 416 536 433
rect 553 416 559 433
rect 530 393 559 416
rect 530 376 536 393
rect 553 376 559 393
rect 586 419 616 434
rect 586 402 592 419
rect 609 402 616 419
rect 586 392 616 402
rect 631 392 658 434
rect 673 423 711 434
rect 673 406 688 423
rect 705 406 711 423
rect 673 392 711 406
rect 530 370 559 376
rect 682 370 711 392
rect 726 423 761 434
rect 726 406 738 423
rect 755 406 761 423
rect 726 370 761 406
rect 788 393 877 454
rect 788 376 794 393
rect 811 376 853 393
rect 870 376 877 393
rect 788 370 877 376
rect 892 370 919 454
rect 934 411 973 454
rect 934 394 940 411
rect 957 394 973 411
rect 934 370 973 394
rect 988 448 1017 454
rect 988 431 994 448
rect 1011 431 1017 448
rect 988 393 1017 431
rect 988 376 994 393
rect 1011 376 1017 393
rect 988 370 1017 376
rect 1044 429 1074 454
rect 1044 412 1050 429
rect 1067 412 1074 429
rect 1044 393 1074 412
rect 1044 376 1050 393
rect 1067 376 1074 393
rect 1044 370 1074 376
rect 1089 370 1113 454
rect 1128 448 1157 454
rect 1128 431 1134 448
rect 1151 431 1157 448
rect 1128 412 1157 431
rect 1278 432 1308 470
rect 1278 415 1284 432
rect 1301 415 1308 432
rect 1128 393 1166 412
rect 1128 376 1134 393
rect 1151 376 1166 393
rect 1128 370 1166 376
rect 1181 370 1205 412
rect 1220 395 1250 412
rect 1220 378 1227 395
rect 1244 378 1250 395
rect 1220 370 1250 378
rect 1278 393 1308 415
rect 1278 376 1284 393
rect 1301 376 1308 393
rect 1278 370 1308 376
rect 1323 395 1359 470
rect 1323 378 1334 395
rect 1351 378 1359 395
rect 1323 370 1359 378
rect 1374 370 1401 470
rect 1416 452 1445 470
rect 1593 466 1620 482
rect 1416 435 1422 452
rect 1439 435 1445 452
rect 1416 393 1445 435
rect 1472 457 1502 466
rect 1472 440 1478 457
rect 1495 440 1502 457
rect 1472 402 1502 440
rect 1517 459 1620 466
rect 1517 442 1588 459
rect 1605 442 1620 459
rect 1517 418 1620 442
rect 1517 402 1588 418
rect 1416 376 1422 393
rect 1439 376 1445 393
rect 1526 401 1588 402
rect 1605 401 1620 418
rect 1416 370 1445 376
rect 1526 373 1620 401
rect 1526 356 1532 373
rect 1549 356 1588 373
rect 1605 370 1620 373
rect 1635 476 1665 482
rect 1635 459 1641 476
rect 1658 459 1665 476
rect 1635 434 1665 459
rect 1635 417 1641 434
rect 1658 417 1665 434
rect 1635 393 1665 417
rect 1635 376 1641 393
rect 1658 376 1665 393
rect 1635 370 1665 376
rect 1680 463 1708 482
rect 1790 474 1817 482
rect 1680 446 1686 463
rect 1703 446 1708 463
rect 1680 428 1708 446
rect 1680 411 1686 428
rect 1703 411 1708 428
rect 1680 393 1708 411
rect 1680 376 1686 393
rect 1703 376 1708 393
rect 1680 370 1708 376
rect 1735 468 1764 474
rect 1735 451 1741 468
rect 1758 451 1764 468
rect 1735 432 1764 451
rect 1735 415 1741 432
rect 1758 415 1764 432
rect 1735 397 1764 415
rect 1735 380 1741 397
rect 1758 380 1764 397
rect 1735 374 1764 380
rect 1779 470 1817 474
rect 1779 453 1793 470
rect 1810 453 1817 470
rect 1779 434 1817 453
rect 1779 417 1793 434
rect 1810 417 1817 434
rect 1779 395 1817 417
rect 1779 378 1793 395
rect 1810 378 1817 395
rect 1779 374 1817 378
rect 1605 356 1611 370
rect 1788 370 1817 374
rect 1832 476 1862 482
rect 1832 459 1838 476
rect 1855 459 1862 476
rect 1832 434 1862 459
rect 1832 417 1838 434
rect 1855 417 1862 434
rect 1832 393 1862 417
rect 1832 376 1838 393
rect 1855 376 1862 393
rect 1832 370 1862 376
rect 1877 476 1906 482
rect 1877 459 1883 476
rect 1900 459 1906 476
rect 1877 434 1906 459
rect 1877 417 1883 434
rect 1900 417 1906 434
rect 1877 393 1906 417
rect 1877 376 1883 393
rect 1900 376 1906 393
rect 1877 370 1906 376
rect 1933 391 2002 482
rect 1933 374 1941 391
rect 1958 374 1977 391
rect 1994 374 2002 391
rect 1933 370 2002 374
rect 2029 473 2059 482
rect 2029 456 2035 473
rect 2052 456 2059 473
rect 2029 433 2059 456
rect 2029 416 2035 433
rect 2052 416 2059 433
rect 2029 393 2059 416
rect 2029 376 2035 393
rect 2052 376 2059 393
rect 2029 370 2059 376
rect 2074 463 2185 482
rect 2074 446 2081 463
rect 2098 446 2121 463
rect 2138 446 2162 463
rect 2179 446 2185 463
rect 2074 427 2185 446
rect 2074 410 2081 427
rect 2098 410 2121 427
rect 2138 410 2162 427
rect 2179 410 2185 427
rect 2074 393 2185 410
rect 2074 376 2081 393
rect 2098 376 2121 393
rect 2138 376 2162 393
rect 2179 376 2185 393
rect 2074 370 2185 376
rect 2200 432 2235 482
rect 2200 415 2207 432
rect 2224 415 2235 432
rect 2200 393 2235 415
rect 2200 376 2207 393
rect 2224 376 2235 393
rect 2200 370 2235 376
rect 2250 463 2385 482
rect 2250 446 2257 463
rect 2274 446 2291 463
rect 2308 446 2327 463
rect 2344 446 2361 463
rect 2378 446 2385 463
rect 2250 427 2385 446
rect 2250 410 2257 427
rect 2274 410 2291 427
rect 2308 410 2327 427
rect 2344 410 2361 427
rect 2378 410 2385 427
rect 2250 393 2385 410
rect 2250 376 2257 393
rect 2274 376 2291 393
rect 2308 376 2327 393
rect 2344 376 2361 393
rect 2378 376 2385 393
rect 2250 370 2385 376
rect 2400 432 2434 482
rect 2400 415 2411 432
rect 2428 415 2434 432
rect 2400 393 2434 415
rect 2400 376 2411 393
rect 2428 376 2434 393
rect 2400 370 2434 376
rect 1526 350 1611 356
rect 1526 309 1611 315
rect -813 290 -779 296
rect -813 273 -807 290
rect -790 273 -779 290
rect -813 255 -779 273
rect -813 238 -807 255
rect -790 238 -779 255
rect -813 220 -779 238
rect -813 203 -807 220
rect -790 203 -779 220
rect -813 184 -779 203
rect -764 290 -734 296
rect -764 273 -757 290
rect -740 273 -734 290
rect -764 248 -734 273
rect -764 231 -757 248
rect -740 231 -734 248
rect -764 207 -734 231
rect -130 290 -102 296
rect -130 273 -125 290
rect -108 273 -102 290
rect -130 248 -102 273
rect -130 231 -125 248
rect -108 231 -102 248
rect -764 190 -757 207
rect -740 190 -734 207
rect -764 184 -734 190
rect -130 207 -102 231
rect -130 190 -125 207
rect -108 190 -102 207
rect -130 184 -102 190
rect -87 290 -57 296
rect -87 273 -80 290
rect -63 273 -57 290
rect -87 248 -57 273
rect -87 231 -80 248
rect -63 231 -57 248
rect -87 207 -57 231
rect -87 190 -80 207
rect -63 190 -57 207
rect -87 184 -57 190
rect -42 290 -13 296
rect -42 273 -35 290
rect -18 273 -13 290
rect -42 248 -13 273
rect -42 231 -35 248
rect -18 231 -13 248
rect -42 207 -13 231
rect 109 290 139 296
rect 109 273 115 290
rect 132 273 139 290
rect 109 255 139 273
rect 109 238 115 255
rect 132 238 139 255
rect 109 232 139 238
rect 154 289 184 296
rect 154 272 160 289
rect 177 272 184 289
rect 154 232 184 272
rect 199 232 223 296
rect 238 260 268 296
rect 238 243 244 260
rect 261 243 268 260
rect 238 232 268 243
rect 283 290 312 296
rect 283 273 289 290
rect 306 273 312 290
rect 283 255 312 273
rect 283 238 289 255
rect 306 238 312 255
rect 283 232 312 238
rect 339 290 369 296
rect 339 273 345 290
rect 362 273 369 290
rect 339 255 369 273
rect 339 238 345 255
rect 362 238 369 255
rect 339 232 369 238
rect 384 290 413 296
rect 384 273 390 290
rect 407 273 413 290
rect 384 255 413 273
rect 384 238 390 255
rect 407 238 413 255
rect 384 232 413 238
rect 440 290 470 296
rect 440 273 446 290
rect 463 273 470 290
rect 440 255 470 273
rect 440 238 446 255
rect 463 238 470 255
rect -42 190 -35 207
rect -18 190 -13 207
rect -42 184 -13 190
rect 440 220 470 238
rect 440 203 446 220
rect 463 203 470 220
rect 440 184 470 203
rect 485 290 515 296
rect 485 273 491 290
rect 508 273 515 290
rect 485 251 515 273
rect 485 234 491 251
rect 508 234 515 251
rect 485 184 515 234
rect 530 290 559 296
rect 530 273 536 290
rect 553 273 559 290
rect 682 274 711 296
rect 530 249 559 273
rect 530 232 536 249
rect 553 232 559 249
rect 586 264 616 274
rect 586 247 592 264
rect 609 247 616 264
rect 586 232 616 247
rect 631 232 658 274
rect 673 260 711 274
rect 673 243 688 260
rect 705 243 711 260
rect 673 232 711 243
rect 726 260 761 296
rect 726 243 738 260
rect 755 243 761 260
rect 726 232 761 243
rect 788 290 877 296
rect 788 273 794 290
rect 811 273 853 290
rect 870 273 877 290
rect 530 209 559 232
rect 530 192 536 209
rect 553 192 559 209
rect 530 184 559 192
rect 788 212 877 273
rect 892 212 919 296
rect 934 271 973 296
rect 934 254 940 271
rect 957 254 973 271
rect 934 212 973 254
rect 988 290 1017 296
rect 988 273 994 290
rect 1011 273 1017 290
rect 988 235 1017 273
rect 988 218 994 235
rect 1011 218 1017 235
rect 988 212 1017 218
rect 1044 290 1074 296
rect 1044 273 1050 290
rect 1067 273 1074 290
rect 1044 254 1074 273
rect 1044 237 1050 254
rect 1067 237 1074 254
rect 1044 212 1074 237
rect 1089 212 1113 296
rect 1128 290 1166 296
rect 1128 273 1134 290
rect 1151 273 1166 290
rect 1128 254 1166 273
rect 1181 254 1205 296
rect 1220 287 1250 296
rect 1220 270 1227 287
rect 1244 270 1250 287
rect 1220 254 1250 270
rect 1278 290 1308 296
rect 1278 273 1284 290
rect 1301 273 1308 290
rect 1128 235 1157 254
rect 1278 251 1308 273
rect 1128 218 1134 235
rect 1151 218 1157 235
rect 1128 212 1157 218
rect 1278 234 1284 251
rect 1301 234 1308 251
rect 1278 196 1308 234
rect 1323 287 1359 296
rect 1323 270 1334 287
rect 1351 270 1359 287
rect 1323 196 1359 270
rect 1374 196 1401 296
rect 1416 290 1445 296
rect 1416 273 1422 290
rect 1439 273 1445 290
rect 1526 292 1532 309
rect 1549 292 1588 309
rect 1605 296 1611 309
rect 1605 292 1620 296
rect 1416 231 1445 273
rect 1526 264 1620 292
rect 1526 263 1588 264
rect 1416 214 1422 231
rect 1439 214 1445 231
rect 1416 196 1445 214
rect 1472 225 1502 263
rect 1472 208 1478 225
rect 1495 208 1502 225
rect 1472 199 1502 208
rect 1517 247 1588 263
rect 1605 247 1620 264
rect 1517 223 1620 247
rect 1517 206 1588 223
rect 1605 206 1620 223
rect 1517 199 1620 206
rect 1593 184 1620 199
rect 1635 290 1665 296
rect 1635 273 1641 290
rect 1658 273 1665 290
rect 1635 248 1665 273
rect 1635 231 1641 248
rect 1658 231 1665 248
rect 1635 207 1665 231
rect 1635 190 1641 207
rect 1658 190 1665 207
rect 1635 184 1665 190
rect 1680 290 1708 296
rect 1788 292 1817 296
rect 1680 273 1686 290
rect 1703 273 1708 290
rect 1680 255 1708 273
rect 1680 238 1686 255
rect 1703 238 1708 255
rect 1680 220 1708 238
rect 1680 203 1686 220
rect 1703 203 1708 220
rect 1680 184 1708 203
rect 1735 286 1764 292
rect 1735 269 1741 286
rect 1758 269 1764 286
rect 1735 250 1764 269
rect 1735 233 1741 250
rect 1758 233 1764 250
rect 1735 215 1764 233
rect 1735 198 1741 215
rect 1758 198 1764 215
rect 1735 192 1764 198
rect 1779 288 1817 292
rect 1779 271 1793 288
rect 1810 271 1817 288
rect 1779 249 1817 271
rect 1779 232 1793 249
rect 1810 232 1817 249
rect 1779 213 1817 232
rect 1779 196 1793 213
rect 1810 196 1817 213
rect 1779 192 1817 196
rect 1790 184 1817 192
rect 1832 290 1862 296
rect 1832 273 1838 290
rect 1855 273 1862 290
rect 1832 248 1862 273
rect 1832 231 1838 248
rect 1855 231 1862 248
rect 1832 207 1862 231
rect 1832 190 1838 207
rect 1855 190 1862 207
rect 1832 184 1862 190
rect 1877 290 1906 296
rect 1877 273 1883 290
rect 1900 273 1906 290
rect 1877 248 1906 273
rect 1877 231 1883 248
rect 1900 231 1906 248
rect 1877 207 1906 231
rect 1877 190 1883 207
rect 1900 190 1906 207
rect 1877 184 1906 190
rect 1933 292 2002 296
rect 1933 275 1941 292
rect 1958 275 1977 292
rect 1994 275 2002 292
rect 2223 290 2253 296
rect 2223 288 2229 290
rect 1933 184 2002 275
rect 2030 282 2059 288
rect 2030 265 2036 282
rect 2053 265 2059 282
rect 2030 227 2059 265
rect 2030 210 2036 227
rect 2053 210 2059 227
rect 2030 204 2059 210
rect 2074 282 2104 288
rect 2074 265 2081 282
rect 2098 265 2104 282
rect 2074 227 2104 265
rect 2074 210 2081 227
rect 2098 210 2104 227
rect 2074 204 2104 210
rect 2119 284 2152 288
rect 2119 267 2126 284
rect 2143 267 2152 284
rect 2119 250 2152 267
rect 2119 233 2126 250
rect 2143 233 2152 250
rect 2119 204 2152 233
rect 2167 282 2199 288
rect 2167 265 2176 282
rect 2193 265 2199 282
rect 2167 227 2199 265
rect 2167 210 2176 227
rect 2193 210 2199 227
rect 2167 204 2199 210
rect 2214 273 2229 288
rect 2246 273 2253 290
rect 2214 254 2253 273
rect 2214 237 2229 254
rect 2246 237 2253 254
rect 2214 204 2253 237
rect 2226 184 2253 204
rect 2268 290 2300 296
rect 2268 273 2276 290
rect 2293 273 2300 290
rect 2268 249 2300 273
rect 2268 232 2276 249
rect 2293 232 2300 249
rect 2268 209 2300 232
rect 2268 192 2276 209
rect 2293 192 2300 209
rect 2268 184 2300 192
rect 2315 290 2345 296
rect 2315 273 2321 290
rect 2338 273 2345 290
rect 2315 243 2345 273
rect 2315 226 2321 243
rect 2338 226 2345 243
rect 2315 184 2345 226
rect 2360 290 2390 296
rect 2360 273 2366 290
rect 2383 273 2390 290
rect 2360 249 2390 273
rect 2360 232 2366 249
rect 2383 232 2390 249
rect 2360 209 2390 232
rect 2360 192 2366 209
rect 2383 192 2390 209
rect 2360 184 2390 192
rect 2405 290 2434 296
rect 2405 273 2411 290
rect 2428 273 2434 290
rect 2405 248 2434 273
rect 2405 231 2411 248
rect 2428 231 2434 248
rect 2405 207 2434 231
rect 2405 190 2411 207
rect 2428 190 2434 207
rect 2405 184 2434 190
<< ndiffc >>
rect -869 1542 -852 1730
rect -825 1542 -808 1730
rect -869 1185 -852 1373
rect -825 1185 -808 1373
rect -478 1542 -461 1730
rect -434 1542 -417 1730
rect -478 1185 -461 1373
rect -434 1185 -417 1373
rect -1383 754 -1366 771
rect -1383 709 -1366 726
rect -1333 754 -1316 771
rect -699 750 -682 767
rect -1333 709 -1316 726
rect -699 709 -682 726
rect -617 750 -600 767
rect -617 709 -600 726
rect -551 721 -534 738
rect -423 721 -406 738
rect -295 721 -278 738
rect 121 721 138 738
rect 249 721 266 738
rect 377 721 394 738
rect 457 721 474 738
rect 585 721 602 738
rect 713 721 730 738
rect 793 721 810 738
rect 921 721 938 738
rect 1049 721 1066 738
rect 1129 721 1146 738
rect 1257 721 1274 738
rect 1385 721 1402 738
rect 1465 721 1482 738
rect 1593 721 1610 738
rect 1721 721 1738 738
rect 1801 721 1818 738
rect 1929 721 1946 738
rect 2057 721 2074 738
rect 2137 721 2154 738
rect 2265 721 2282 738
rect -1383 606 -1366 623
rect -1383 561 -1366 578
rect -1333 606 -1316 623
rect -699 606 -682 623
rect -1333 561 -1316 578
rect -699 565 -682 582
rect -617 606 -600 623
rect -617 565 -600 582
rect -556 574 -539 591
rect -503 606 -486 623
rect -512 561 -495 578
rect -405 602 -388 619
rect -238 593 -221 610
rect -181 606 -164 623
rect -181 561 -164 578
rect -123 606 -106 623
rect -123 561 -106 578
rect -80 606 -63 623
rect -80 561 -63 578
rect -37 606 -20 623
rect -37 561 -20 578
rect 497 625 514 642
rect 118 581 135 598
rect 200 578 217 595
rect 240 578 257 595
rect 322 581 339 598
rect 390 576 407 593
rect 446 549 463 566
rect 573 581 590 598
rect 573 547 590 564
rect 642 607 659 624
rect 843 606 860 623
rect 732 574 749 591
rect 782 576 799 593
rect 899 571 916 588
rect 954 580 971 597
rect 1009 580 1026 597
rect 1100 589 1117 606
rect 1141 589 1158 606
rect 1182 589 1199 606
rect 1274 623 1291 640
rect 1332 606 1349 623
rect 1379 580 1396 597
rect 1430 616 1447 633
rect 1589 606 1606 623
rect 1486 540 1503 557
rect 1589 561 1606 578
rect 1632 606 1649 623
rect 1632 561 1649 578
rect 1675 606 1692 623
rect 1675 561 1692 578
rect 1738 593 1755 610
rect 1738 559 1755 576
rect 1791 606 1808 623
rect 1791 569 1808 586
rect 1841 606 1858 623
rect 1841 569 1858 586
rect 1884 606 1901 623
rect 1884 561 1901 578
rect 1941 608 1958 625
rect 1977 608 1994 625
rect 2035 606 2052 623
rect 2035 561 2052 578
rect 2078 595 2095 612
rect 2121 606 2138 623
rect 2121 561 2138 578
rect 2164 595 2181 612
rect 2207 606 2224 623
rect 2207 561 2224 578
rect 2257 579 2274 596
rect 2307 595 2324 612
rect 2359 579 2376 596
rect 2411 595 2428 612
rect -807 88 -790 105
rect -807 43 -790 60
rect -757 88 -740 105
rect -123 84 -106 101
rect -757 43 -740 60
rect -123 43 -106 60
rect -41 84 -24 101
rect -41 43 -24 60
rect 118 68 135 85
rect 200 70 217 87
rect 240 70 257 87
rect 322 67 339 84
rect 390 73 407 90
rect 446 100 463 117
rect 573 101 590 118
rect 573 67 590 84
rect 732 75 749 92
rect 782 72 799 89
rect 899 77 916 94
rect 954 68 971 85
rect 1009 68 1026 85
rect 497 24 514 41
rect 642 42 659 59
rect 843 42 860 59
rect 1100 60 1117 77
rect 1141 60 1158 77
rect 1182 60 1199 77
rect 1274 26 1291 43
rect 1332 43 1349 60
rect 1379 69 1396 86
rect 1486 108 1503 125
rect 1589 88 1606 105
rect 1430 32 1447 49
rect 1589 43 1606 60
rect 1632 88 1649 105
rect 1632 43 1649 60
rect 1675 88 1692 105
rect 1675 43 1692 60
rect 1738 90 1755 107
rect 1738 56 1755 73
rect 1791 80 1808 97
rect 1791 43 1808 60
rect 1841 80 1858 97
rect 1841 43 1858 60
rect 1884 88 1901 105
rect 1884 43 1901 60
rect 2035 100 2052 117
rect 2035 65 2052 82
rect 2080 67 2097 84
rect 2123 102 2140 119
rect 2123 63 2140 80
rect 2173 97 2190 114
rect 2173 63 2190 80
rect 2224 100 2241 117
rect 2224 61 2241 78
rect 1941 41 1958 58
rect 1977 41 1994 58
rect 2275 92 2292 109
rect 2275 55 2292 72
rect 2325 58 2342 75
rect 2368 100 2385 117
rect 2368 55 2385 72
rect 2411 100 2428 117
rect 2411 55 2428 72
rect -694 -343 -677 -155
rect -650 -343 -633 -155
rect -694 -700 -677 -512
rect -650 -700 -633 -512
<< pdiffc >>
rect -1383 939 -1366 956
rect -1383 904 -1366 921
rect -1383 869 -1366 886
rect -1333 939 -1316 956
rect -1333 897 -1316 914
rect -701 939 -684 956
rect -701 897 -684 914
rect -1333 856 -1316 873
rect -701 856 -684 873
rect -656 939 -639 956
rect -656 897 -639 914
rect -656 856 -639 873
rect -611 939 -594 956
rect -611 897 -594 914
rect -611 856 -594 873
rect -558 939 -541 956
rect -558 903 -541 920
rect -558 868 -541 885
rect -429 939 -412 956
rect -429 903 -412 920
rect -429 868 -412 885
rect -302 939 -285 956
rect -302 903 -285 920
rect -302 868 -285 885
rect 113 939 130 956
rect 113 903 130 920
rect 113 868 130 885
rect 242 939 259 956
rect 242 903 259 920
rect 242 868 259 885
rect 370 939 387 956
rect 370 903 387 920
rect 370 868 387 885
rect 449 939 466 956
rect 449 903 466 920
rect 449 868 466 885
rect 578 939 595 956
rect 578 903 595 920
rect 578 868 595 885
rect 706 939 723 956
rect 706 903 723 920
rect 706 868 723 885
rect 785 939 802 956
rect 785 903 802 920
rect 785 868 802 885
rect 914 939 931 956
rect 914 903 931 920
rect 914 868 931 885
rect 1042 939 1059 956
rect 1042 903 1059 920
rect 1042 868 1059 885
rect 1121 939 1138 956
rect 1121 903 1138 920
rect 1121 868 1138 885
rect 1250 939 1267 956
rect 1250 903 1267 920
rect 1250 868 1267 885
rect 1378 939 1395 956
rect 1378 903 1395 920
rect 1378 868 1395 885
rect 1457 939 1474 956
rect 1457 903 1474 920
rect 1457 868 1474 885
rect 1586 939 1603 956
rect 1586 903 1603 920
rect 1586 868 1603 885
rect 1714 939 1731 956
rect 1714 903 1731 920
rect 1714 868 1731 885
rect 1793 939 1810 956
rect 1793 903 1810 920
rect 1793 868 1810 885
rect 1922 939 1939 956
rect 1922 903 1939 920
rect 1922 868 1939 885
rect 2050 939 2067 956
rect 2050 903 2067 920
rect 2050 868 2067 885
rect 2129 939 2146 956
rect 2129 903 2146 920
rect 2129 868 2146 885
rect 2258 939 2275 956
rect 2258 903 2275 920
rect 2258 868 2275 885
rect -1383 446 -1366 463
rect -1383 411 -1366 428
rect -1383 376 -1366 393
rect -1333 459 -1316 476
rect -701 459 -684 476
rect -1333 417 -1316 434
rect -1333 376 -1316 393
rect -701 417 -684 434
rect -701 376 -684 393
rect -656 459 -639 476
rect -656 417 -639 434
rect -656 376 -639 393
rect -611 459 -594 476
rect -611 417 -594 434
rect -556 451 -539 468
rect -556 404 -539 421
rect -503 406 -486 423
rect -611 376 -594 393
rect -361 459 -344 476
rect -361 400 -344 417
rect -238 459 -221 476
rect -238 417 -221 434
rect -238 376 -221 393
rect -188 459 -171 476
rect -188 417 -171 434
rect -188 376 -171 393
rect -125 446 -108 463
rect -125 411 -108 428
rect -125 376 -108 393
rect -80 459 -63 476
rect -80 417 -63 434
rect -80 376 -63 393
rect -35 459 -18 476
rect -35 417 -18 434
rect -35 376 -18 393
rect 446 446 463 463
rect 115 410 132 427
rect 115 376 132 393
rect 160 376 177 393
rect 244 406 261 423
rect 289 411 306 428
rect 289 376 306 393
rect 345 411 362 428
rect 345 376 362 393
rect 390 411 407 428
rect 390 376 407 393
rect 446 411 463 428
rect 446 376 463 393
rect 491 415 508 432
rect 491 376 508 393
rect 536 457 553 474
rect 536 416 553 433
rect 536 376 553 393
rect 592 402 609 419
rect 688 406 705 423
rect 738 406 755 423
rect 794 376 811 393
rect 853 376 870 393
rect 940 394 957 411
rect 994 431 1011 448
rect 994 376 1011 393
rect 1050 412 1067 429
rect 1050 376 1067 393
rect 1134 431 1151 448
rect 1284 415 1301 432
rect 1134 376 1151 393
rect 1227 378 1244 395
rect 1284 376 1301 393
rect 1334 378 1351 395
rect 1422 435 1439 452
rect 1478 440 1495 457
rect 1588 442 1605 459
rect 1422 376 1439 393
rect 1588 401 1605 418
rect 1532 356 1549 373
rect 1588 356 1605 373
rect 1641 459 1658 476
rect 1641 417 1658 434
rect 1641 376 1658 393
rect 1686 446 1703 463
rect 1686 411 1703 428
rect 1686 376 1703 393
rect 1741 451 1758 468
rect 1741 415 1758 432
rect 1741 380 1758 397
rect 1793 453 1810 470
rect 1793 417 1810 434
rect 1793 378 1810 395
rect 1838 459 1855 476
rect 1838 417 1855 434
rect 1838 376 1855 393
rect 1883 459 1900 476
rect 1883 417 1900 434
rect 1883 376 1900 393
rect 1941 374 1958 391
rect 1977 374 1994 391
rect 2035 456 2052 473
rect 2035 416 2052 433
rect 2035 376 2052 393
rect 2081 446 2098 463
rect 2121 446 2138 463
rect 2162 446 2179 463
rect 2081 410 2098 427
rect 2121 410 2138 427
rect 2162 410 2179 427
rect 2081 376 2098 393
rect 2121 376 2138 393
rect 2162 376 2179 393
rect 2207 415 2224 432
rect 2207 376 2224 393
rect 2257 446 2274 463
rect 2291 446 2308 463
rect 2327 446 2344 463
rect 2361 446 2378 463
rect 2257 410 2274 427
rect 2291 410 2308 427
rect 2327 410 2344 427
rect 2361 410 2378 427
rect 2257 376 2274 393
rect 2291 376 2308 393
rect 2327 376 2344 393
rect 2361 376 2378 393
rect 2411 415 2428 432
rect 2411 376 2428 393
rect -807 273 -790 290
rect -807 238 -790 255
rect -807 203 -790 220
rect -757 273 -740 290
rect -757 231 -740 248
rect -125 273 -108 290
rect -125 231 -108 248
rect -757 190 -740 207
rect -125 190 -108 207
rect -80 273 -63 290
rect -80 231 -63 248
rect -80 190 -63 207
rect -35 273 -18 290
rect -35 231 -18 248
rect 115 273 132 290
rect 115 238 132 255
rect 160 272 177 289
rect 244 243 261 260
rect 289 273 306 290
rect 289 238 306 255
rect 345 273 362 290
rect 345 238 362 255
rect 390 273 407 290
rect 390 238 407 255
rect 446 273 463 290
rect 446 238 463 255
rect -35 190 -18 207
rect 446 203 463 220
rect 491 273 508 290
rect 491 234 508 251
rect 536 273 553 290
rect 536 232 553 249
rect 592 247 609 264
rect 688 243 705 260
rect 738 243 755 260
rect 794 273 811 290
rect 853 273 870 290
rect 536 192 553 209
rect 940 254 957 271
rect 994 273 1011 290
rect 994 218 1011 235
rect 1050 273 1067 290
rect 1050 237 1067 254
rect 1134 273 1151 290
rect 1227 270 1244 287
rect 1284 273 1301 290
rect 1134 218 1151 235
rect 1284 234 1301 251
rect 1334 270 1351 287
rect 1422 273 1439 290
rect 1532 292 1549 309
rect 1588 292 1605 309
rect 1422 214 1439 231
rect 1478 208 1495 225
rect 1588 247 1605 264
rect 1588 206 1605 223
rect 1641 273 1658 290
rect 1641 231 1658 248
rect 1641 190 1658 207
rect 1686 273 1703 290
rect 1686 238 1703 255
rect 1686 203 1703 220
rect 1741 269 1758 286
rect 1741 233 1758 250
rect 1741 198 1758 215
rect 1793 271 1810 288
rect 1793 232 1810 249
rect 1793 196 1810 213
rect 1838 273 1855 290
rect 1838 231 1855 248
rect 1838 190 1855 207
rect 1883 273 1900 290
rect 1883 231 1900 248
rect 1883 190 1900 207
rect 1941 275 1958 292
rect 1977 275 1994 292
rect 2036 265 2053 282
rect 2036 210 2053 227
rect 2081 265 2098 282
rect 2081 210 2098 227
rect 2126 267 2143 284
rect 2126 233 2143 250
rect 2176 265 2193 282
rect 2176 210 2193 227
rect 2229 273 2246 290
rect 2229 237 2246 254
rect 2276 273 2293 290
rect 2276 232 2293 249
rect 2276 192 2293 209
rect 2321 273 2338 290
rect 2321 226 2338 243
rect 2366 273 2383 290
rect 2366 232 2383 249
rect 2366 192 2383 209
rect 2411 273 2428 290
rect 2411 231 2428 248
rect 2411 190 2428 207
<< psubdiff >>
rect -926 1806 -878 1823
rect -799 1806 -751 1823
rect -926 1775 -909 1806
rect -768 1775 -751 1806
rect -926 1466 -909 1497
rect -768 1466 -751 1497
rect -926 1449 -878 1466
rect -799 1449 -751 1466
rect -926 1418 -909 1449
rect -768 1418 -751 1449
rect -926 1109 -909 1140
rect -768 1109 -751 1140
rect -926 1092 -878 1109
rect -799 1092 -751 1109
rect -535 1806 -487 1823
rect -408 1806 -360 1823
rect -535 1775 -518 1806
rect -377 1775 -360 1806
rect -535 1466 -518 1497
rect -377 1466 -360 1497
rect -535 1449 -487 1466
rect -408 1449 -360 1466
rect -535 1418 -518 1449
rect -377 1418 -360 1449
rect -535 1109 -518 1140
rect -377 1109 -360 1140
rect -535 1092 -487 1109
rect -408 1092 -360 1109
rect 15 768 80 780
rect 32 751 63 768
rect 15 727 80 751
rect 32 710 63 727
rect 15 698 80 710
rect 15 622 80 634
rect 32 605 63 622
rect 15 580 80 605
rect 32 563 63 580
rect 15 551 80 563
rect 15 102 80 114
rect 32 85 63 102
rect 15 61 80 85
rect 32 44 63 61
rect 15 32 80 44
rect -751 -79 -703 -62
rect -624 -79 -576 -62
rect -751 -110 -734 -79
rect -593 -110 -576 -79
rect -751 -419 -734 -388
rect -593 -419 -576 -388
rect -751 -436 -703 -419
rect -624 -436 -576 -419
rect -751 -467 -734 -436
rect -593 -467 -576 -436
rect -751 -776 -734 -745
rect -593 -776 -576 -745
rect -751 -793 -703 -776
rect -624 -793 -576 -776
<< nsubdiff >>
rect 15 955 80 967
rect 32 938 63 955
rect 15 912 80 938
rect 32 895 63 912
rect 15 883 80 895
rect 15 437 80 449
rect 32 420 63 437
rect 15 394 80 420
rect 32 377 63 394
rect 15 365 80 377
rect 15 289 80 301
rect 32 272 63 289
rect 15 246 80 272
rect 32 229 63 246
rect 15 217 80 229
<< psubdiffcont >>
rect -878 1806 -799 1823
rect -926 1497 -909 1775
rect -768 1497 -751 1775
rect -878 1449 -799 1466
rect -926 1140 -909 1418
rect -768 1140 -751 1418
rect -878 1092 -799 1109
rect -487 1806 -408 1823
rect -535 1497 -518 1775
rect -377 1497 -360 1775
rect -487 1449 -408 1466
rect -535 1140 -518 1418
rect -377 1140 -360 1418
rect -487 1092 -408 1109
rect 15 751 32 768
rect 63 751 80 768
rect 15 710 32 727
rect 63 710 80 727
rect 15 605 32 622
rect 63 605 80 622
rect 15 563 32 580
rect 63 563 80 580
rect 15 85 32 102
rect 63 85 80 102
rect 15 44 32 61
rect 63 44 80 61
rect -703 -79 -624 -62
rect -751 -388 -734 -110
rect -593 -388 -576 -110
rect -703 -436 -624 -419
rect -751 -745 -734 -467
rect -593 -745 -576 -467
rect -703 -793 -624 -776
<< nsubdiffcont >>
rect 15 938 32 955
rect 63 938 80 955
rect 15 895 32 912
rect 63 895 80 912
rect 15 420 32 437
rect 63 420 80 437
rect 15 377 32 394
rect 63 377 80 394
rect 15 272 32 289
rect 63 272 80 289
rect 15 229 32 246
rect 63 229 80 246
<< poly >>
rect -855 1747 -822 1780
rect -846 1736 -831 1747
rect -846 1525 -831 1536
rect -855 1517 -822 1525
rect -855 1500 -847 1517
rect -830 1500 -822 1517
rect -855 1492 -822 1500
rect -855 1390 -822 1423
rect -846 1379 -831 1390
rect -846 1168 -831 1179
rect -855 1160 -822 1168
rect -855 1143 -847 1160
rect -830 1143 -822 1160
rect -855 1135 -822 1143
rect -464 1747 -431 1780
rect -455 1736 -440 1747
rect -455 1525 -440 1536
rect -464 1517 -431 1525
rect -464 1500 -456 1517
rect -439 1500 -431 1517
rect -464 1492 -431 1500
rect -464 1390 -431 1423
rect -455 1379 -440 1390
rect -455 1168 -440 1179
rect -464 1160 -431 1168
rect -464 1143 -456 1160
rect -439 1143 -431 1160
rect -464 1135 -431 1143
rect -1355 962 -1340 975
rect -678 962 -663 975
rect -633 962 -618 975
rect -535 962 -435 975
rect -407 962 -307 975
rect -1355 842 -1340 850
rect -1356 829 -1338 842
rect -1425 825 -1338 829
rect -1426 821 -1338 825
rect -1426 804 -1417 821
rect -1400 804 -1383 821
rect -1366 804 -1338 821
rect -1426 799 -1338 804
rect -1425 796 -1338 799
rect -1354 777 -1339 796
rect 137 962 237 975
rect 264 962 364 975
rect 473 962 573 975
rect 600 962 700 975
rect 809 962 909 975
rect 936 962 1036 975
rect 1145 962 1245 975
rect 1272 962 1372 975
rect 1481 962 1581 975
rect 1608 962 1708 975
rect 1817 962 1917 975
rect 1944 962 2044 975
rect 2153 962 2253 975
rect -678 842 -663 850
rect -633 842 -618 850
rect -535 849 -435 862
rect -407 849 -307 862
rect -679 821 -661 842
rect -634 821 -616 842
rect -709 813 -661 821
rect -709 796 -701 813
rect -684 796 -661 813
rect -709 788 -661 796
rect -676 777 -661 788
rect -637 813 -586 821
rect -637 796 -611 813
rect -594 796 -586 813
rect -637 788 -586 796
rect -535 816 -502 849
rect -535 799 -527 816
rect -510 799 -502 816
rect -535 791 -502 799
rect -461 816 -368 824
rect -461 799 -453 816
rect -436 799 -393 816
rect -376 799 -368 816
rect -637 777 -622 788
rect -461 785 -368 799
rect -340 816 -307 849
rect -340 799 -332 816
rect -315 799 -307 816
rect -340 791 -307 799
rect 137 849 237 862
rect 264 849 364 862
rect 137 816 170 849
rect 137 799 145 816
rect 162 799 170 816
rect 137 791 170 799
rect 210 816 304 824
rect 210 799 218 816
rect 235 799 279 816
rect 296 799 304 816
rect -461 770 -428 785
rect -528 750 -428 770
rect -400 770 -368 785
rect 210 785 304 799
rect 331 816 364 849
rect 331 799 339 816
rect 356 799 364 816
rect 331 791 364 799
rect 473 849 573 862
rect 600 849 700 862
rect 473 816 506 849
rect 473 799 481 816
rect 498 799 506 816
rect 473 791 506 799
rect 546 816 640 824
rect 546 799 554 816
rect 571 799 615 816
rect 632 799 640 816
rect -400 750 -300 770
rect 210 770 243 785
rect 143 750 243 770
rect 271 770 304 785
rect 546 785 640 799
rect 667 816 700 849
rect 667 799 675 816
rect 692 799 700 816
rect 667 791 700 799
rect 809 849 909 862
rect 936 849 1036 862
rect 809 816 842 849
rect 809 799 817 816
rect 834 799 842 816
rect 809 791 842 799
rect 882 816 976 824
rect 882 799 890 816
rect 907 799 951 816
rect 968 799 976 816
rect 546 770 579 785
rect 271 750 371 770
rect 479 750 579 770
rect 607 770 640 785
rect 882 785 976 799
rect 1003 816 1036 849
rect 1003 799 1011 816
rect 1028 799 1036 816
rect 1003 791 1036 799
rect 1145 849 1245 862
rect 1272 849 1372 862
rect 1145 816 1178 849
rect 1145 799 1153 816
rect 1170 799 1178 816
rect 1145 791 1178 799
rect 1218 816 1312 824
rect 1218 799 1226 816
rect 1243 799 1287 816
rect 1304 799 1312 816
rect 882 770 915 785
rect 607 750 707 770
rect 815 750 915 770
rect 943 770 976 785
rect 1218 785 1312 799
rect 1339 816 1372 849
rect 1339 799 1347 816
rect 1364 799 1372 816
rect 1339 791 1372 799
rect 1481 849 1581 862
rect 1608 849 1708 862
rect 1481 816 1514 849
rect 1481 799 1489 816
rect 1506 799 1514 816
rect 1481 791 1514 799
rect 1554 816 1648 824
rect 1554 799 1562 816
rect 1579 799 1623 816
rect 1640 799 1648 816
rect 1218 770 1251 785
rect 943 750 1043 770
rect 1151 750 1251 770
rect 1279 770 1312 785
rect 1554 785 1648 799
rect 1675 816 1708 849
rect 1675 799 1683 816
rect 1700 799 1708 816
rect 1675 791 1708 799
rect 1817 849 1917 862
rect 1944 849 2044 862
rect 1817 816 1850 849
rect 1817 799 1825 816
rect 1842 799 1850 816
rect 1817 791 1850 799
rect 1890 816 1984 824
rect 1890 799 1898 816
rect 1915 799 1959 816
rect 1976 799 1984 816
rect 1554 770 1587 785
rect 1279 750 1379 770
rect 1487 750 1587 770
rect 1615 770 1648 785
rect 1890 785 1984 799
rect 2011 816 2044 849
rect 2011 799 2019 816
rect 2036 799 2044 816
rect 2011 791 2044 799
rect 2153 849 2253 862
rect 2153 816 2186 849
rect 2153 799 2161 816
rect 2178 799 2186 816
rect 2153 791 2186 799
rect 2226 816 2259 824
rect 2226 799 2234 816
rect 2251 799 2259 816
rect 1890 770 1923 785
rect 1615 750 1715 770
rect 1823 750 1923 770
rect 1951 770 1984 785
rect 2226 770 2259 799
rect 1951 750 2051 770
rect 2159 750 2259 770
rect -1354 690 -1339 703
rect -676 690 -661 703
rect -637 690 -622 703
rect -528 689 -428 708
rect -400 689 -300 708
rect 143 689 243 708
rect 271 689 371 708
rect 479 689 579 708
rect 607 689 707 708
rect 815 689 915 708
rect 943 689 1043 708
rect 1151 689 1251 708
rect 1279 689 1379 708
rect 1487 689 1587 708
rect 1615 689 1715 708
rect 1823 689 1923 708
rect 1951 689 2051 708
rect 2159 689 2259 708
rect -1354 629 -1339 642
rect -676 629 -661 642
rect -637 629 -622 642
rect -478 629 -463 642
rect -439 629 -424 642
rect -369 629 -354 642
rect -273 629 -258 642
rect -202 629 -187 642
rect -100 629 -85 642
rect -57 629 -42 642
rect 179 640 384 655
rect -1354 536 -1339 555
rect -1425 532 -1338 536
rect -1426 528 -1338 532
rect -1426 511 -1417 528
rect -1400 511 -1383 528
rect -1366 511 -1338 528
rect -1426 506 -1338 511
rect -1425 503 -1338 506
rect -1356 489 -1338 503
rect -1355 482 -1340 489
rect -534 610 -519 623
rect 140 606 155 619
rect 179 606 194 640
rect 262 606 277 619
rect 301 606 316 619
rect 369 606 384 640
rect 468 617 483 630
rect 552 640 1094 655
rect 552 617 567 640
rect -676 544 -661 555
rect -709 536 -661 544
rect -709 519 -701 536
rect -684 519 -661 536
rect -709 511 -661 519
rect -637 544 -622 555
rect -637 536 -586 544
rect -637 519 -611 536
rect -594 519 -586 536
rect -637 511 -586 519
rect -534 531 -519 555
rect -478 531 -463 555
rect -439 544 -424 555
rect -369 544 -354 555
rect -534 523 -463 531
rect -679 489 -661 511
rect -634 489 -616 511
rect -534 506 -517 523
rect -500 506 -463 523
rect -441 536 -408 544
rect -441 519 -433 536
rect -416 519 -408 536
rect -441 511 -408 519
rect -387 536 -354 544
rect -387 519 -379 536
rect -362 519 -354 536
rect -387 511 -354 519
rect -330 536 -297 544
rect -330 519 -322 536
rect -305 519 -297 536
rect -330 511 -297 519
rect -273 534 -258 555
rect -202 536 -187 555
rect -100 536 -85 555
rect -57 536 -42 555
rect 140 553 155 564
rect 179 553 194 564
rect 118 545 155 553
rect -273 526 -240 534
rect -534 498 -463 506
rect -534 489 -516 498
rect -481 489 -463 498
rect -384 489 -366 511
rect -330 489 -312 511
rect -273 509 -265 526
rect -248 509 -240 526
rect -273 501 -240 509
rect -219 528 -186 536
rect -219 511 -211 528
rect -194 511 -186 528
rect -219 503 -186 511
rect -133 528 -40 536
rect -133 511 -125 528
rect -108 521 -40 528
rect -108 511 -85 521
rect -133 503 -85 511
rect -273 489 -255 501
rect -211 489 -193 503
rect -103 489 -85 503
rect -58 489 -40 521
rect 118 528 126 545
rect 143 528 155 545
rect 118 511 155 528
rect 118 494 126 511
rect 143 494 155 511
rect -678 482 -663 489
rect -633 482 -618 489
rect -533 482 -518 489
rect -479 482 -464 489
rect -383 482 -368 489
rect -329 482 -314 489
rect -272 482 -257 489
rect -210 482 -195 489
rect -102 482 -87 489
rect -57 482 -42 489
rect -533 385 -518 398
rect -1355 357 -1340 370
rect -678 357 -663 370
rect -633 357 -618 370
rect -479 369 -464 382
rect -383 369 -368 382
rect -329 369 -314 382
rect -272 369 -257 382
rect 118 477 155 494
rect 176 545 209 553
rect 176 528 184 545
rect 201 528 209 545
rect 176 511 209 528
rect 262 520 277 564
rect 176 494 184 511
rect 201 494 209 511
rect 176 486 209 494
rect 230 512 277 520
rect 230 495 252 512
rect 269 495 277 512
rect 230 487 277 495
rect 301 500 316 564
rect 369 557 384 564
rect 369 542 428 557
rect 673 603 688 616
rect 709 603 724 640
rect 1079 625 1094 640
rect 1204 625 1219 638
rect 1243 625 1258 638
rect 755 603 770 616
rect 878 603 893 616
rect 921 603 936 616
rect 982 603 997 616
rect 1032 603 1047 616
rect 673 554 688 561
rect 356 510 389 518
rect 356 500 364 510
rect 301 493 364 500
rect 381 493 389 510
rect 118 460 126 477
rect 143 460 155 477
rect 118 452 155 460
rect 137 441 155 452
rect 182 441 200 486
rect 230 462 245 487
rect 221 447 245 462
rect 301 485 389 493
rect 301 461 316 485
rect 413 461 428 542
rect 468 531 483 543
rect 552 532 567 543
rect 452 523 486 531
rect 452 506 460 523
rect 477 506 486 523
rect 452 498 486 506
rect 507 524 567 532
rect 507 507 515 524
rect 532 507 567 524
rect 507 499 567 507
rect 616 539 688 554
rect 468 489 486 498
rect 513 489 531 499
rect 470 482 485 489
rect 515 482 530 489
rect 616 483 631 539
rect 655 507 688 515
rect 655 490 663 507
rect 680 490 688 507
rect 221 441 239 447
rect 266 446 316 461
rect 367 446 428 461
rect 266 441 284 446
rect 367 441 385 446
rect 139 434 154 441
rect 184 434 199 441
rect 223 434 238 441
rect 268 434 283 441
rect 369 434 384 441
rect -210 357 -195 370
rect -102 357 -87 370
rect -57 357 -42 370
rect 599 475 632 483
rect 655 482 688 490
rect 599 458 607 475
rect 624 458 632 475
rect 599 450 632 458
rect 614 441 632 450
rect 656 441 674 482
rect 709 456 724 561
rect 755 513 770 561
rect 1307 629 1322 642
rect 1359 629 1374 642
rect 1402 629 1417 642
rect 1079 562 1094 570
rect 878 537 893 548
rect 921 537 936 548
rect 799 529 893 537
rect 745 505 778 513
rect 745 488 753 505
rect 770 488 778 505
rect 745 480 778 488
rect 799 512 807 529
rect 824 522 893 529
rect 824 512 832 522
rect 799 495 832 512
rect 799 478 807 495
rect 824 478 832 495
rect 799 470 832 478
rect 875 461 893 522
rect 917 529 950 537
rect 917 512 925 529
rect 942 512 950 529
rect 982 521 997 548
rect 917 495 950 512
rect 917 478 925 495
rect 942 478 950 495
rect 917 470 950 478
rect 971 513 1008 521
rect 971 496 983 513
rect 1000 496 1008 513
rect 971 488 1008 496
rect 1032 508 1047 548
rect 1079 547 1180 562
rect 1111 515 1144 523
rect 1032 500 1090 508
rect 917 461 935 470
rect 971 461 989 488
rect 1032 483 1065 500
rect 1082 483 1090 500
rect 1032 475 1090 483
rect 1072 461 1090 475
rect 1111 498 1119 515
rect 1136 498 1144 515
rect 1111 490 1144 498
rect 1111 461 1129 490
rect 1165 466 1180 547
rect 1204 539 1219 583
rect 1243 575 1258 583
rect 1243 560 1270 575
rect 1201 531 1234 539
rect 1201 514 1209 531
rect 1226 514 1234 531
rect 1201 506 1234 514
rect 709 441 728 456
rect 877 454 892 461
rect 919 454 934 461
rect 973 454 988 461
rect 1074 454 1089 461
rect 1113 454 1128 461
rect 616 434 631 441
rect 658 434 673 441
rect 711 434 726 441
rect 616 379 631 392
rect 658 379 673 392
rect 1165 419 1183 466
rect 1255 461 1270 560
rect 1611 629 1626 642
rect 1654 629 1669 642
rect 1508 576 1523 589
rect 1307 544 1322 555
rect 1359 544 1374 555
rect 1291 536 1324 544
rect 1291 519 1299 536
rect 1316 519 1324 536
rect 1291 511 1324 519
rect 1345 536 1378 544
rect 1345 519 1353 536
rect 1370 519 1378 536
rect 1402 519 1417 555
rect 1760 619 1775 632
rect 1820 629 1835 642
rect 1863 629 1878 642
rect 2058 629 2073 642
rect 2101 629 2116 642
rect 2144 629 2159 642
rect 2187 629 2202 642
rect 2234 629 2249 642
rect 2280 629 2295 642
rect 2330 629 2345 642
rect 2386 629 2401 642
rect 1345 511 1378 519
rect 1399 511 1432 519
rect 1508 515 1523 534
rect 1611 531 1626 555
rect 1654 531 1669 555
rect 1760 531 1775 555
rect 1820 544 1835 555
rect 1863 544 1878 555
rect 1799 536 1878 544
rect 1611 523 1778 531
rect 1306 477 1324 511
rect 1357 477 1375 511
rect 1399 494 1407 511
rect 1424 494 1432 511
rect 1399 486 1432 494
rect 1490 507 1523 515
rect 1490 490 1498 507
rect 1515 490 1523 507
rect 1544 515 1778 523
rect 1544 498 1552 515
rect 1569 501 1778 515
rect 1799 519 1807 536
rect 1824 519 1878 536
rect 1799 511 1878 519
rect 1569 498 1577 501
rect 1544 490 1577 498
rect 1399 477 1417 486
rect 1490 482 1523 490
rect 1618 489 1636 501
rect 1663 489 1681 501
rect 1620 482 1635 489
rect 1665 482 1680 489
rect 1308 470 1323 477
rect 1359 470 1374 477
rect 1401 470 1416 477
rect 1500 474 1518 482
rect 1204 453 1270 461
rect 1204 436 1212 453
rect 1229 446 1270 453
rect 1229 436 1237 446
rect 1204 428 1237 436
rect 1204 419 1222 428
rect 1166 412 1181 419
rect 1205 412 1220 419
rect 1502 466 1517 474
rect 1502 389 1517 402
rect 139 357 154 370
rect 184 357 199 370
rect 223 357 238 370
rect 268 357 283 370
rect 369 357 384 370
rect 470 357 485 370
rect 515 357 530 370
rect 711 357 726 370
rect 877 357 892 370
rect 919 357 934 370
rect 973 357 988 370
rect 1074 357 1089 370
rect 1113 357 1128 370
rect 1166 357 1181 370
rect 1205 357 1220 370
rect 1308 357 1323 370
rect 1359 357 1374 370
rect 1401 357 1416 370
rect 1763 481 1781 501
rect 1815 489 1833 511
rect 1860 489 1878 511
rect 2058 531 2073 555
rect 2101 531 2116 555
rect 2144 531 2159 555
rect 2187 531 2202 555
rect 2058 523 2202 531
rect 2058 506 2075 523
rect 2092 506 2109 523
rect 2126 506 2143 523
rect 2160 506 2177 523
rect 2194 506 2202 523
rect 2058 498 2202 506
rect 2058 489 2076 498
rect 2184 489 2202 498
rect 2234 531 2249 555
rect 2280 531 2295 555
rect 2330 531 2345 555
rect 2386 531 2401 555
rect 2234 523 2401 531
rect 2234 506 2268 523
rect 2285 506 2302 523
rect 2319 506 2336 523
rect 2353 506 2370 523
rect 2387 506 2401 523
rect 2234 498 2401 506
rect 2234 489 2252 498
rect 2383 489 2401 498
rect 1817 482 1832 489
rect 1862 482 1877 489
rect 2059 482 2074 489
rect 2185 482 2200 489
rect 2235 482 2250 489
rect 2385 482 2400 489
rect 1764 474 1779 481
rect 1620 357 1635 370
rect 1665 357 1680 370
rect 1764 361 1779 374
rect 1817 357 1832 370
rect 1862 357 1877 370
rect 2059 357 2074 370
rect 2185 357 2200 370
rect 2235 357 2250 370
rect 2385 357 2400 370
rect -779 296 -764 309
rect -102 296 -87 309
rect -57 296 -42 309
rect -779 176 -764 184
rect -780 163 -762 176
rect -849 159 -762 163
rect -850 155 -762 159
rect -850 138 -841 155
rect -824 138 -807 155
rect -790 138 -762 155
rect -850 133 -762 138
rect -849 130 -762 133
rect -778 111 -763 130
rect 139 296 154 309
rect 184 296 199 309
rect 223 296 238 309
rect 268 296 283 309
rect 369 296 384 309
rect 470 296 485 309
rect 515 296 530 309
rect 711 296 726 309
rect 877 296 892 309
rect 919 296 934 309
rect 973 296 988 309
rect 1074 296 1089 309
rect 1113 296 1128 309
rect 1166 296 1181 309
rect 1205 296 1220 309
rect 1308 296 1323 309
rect 1359 296 1374 309
rect 1401 296 1416 309
rect 139 224 154 232
rect 184 224 199 232
rect 223 224 238 232
rect 268 224 283 232
rect 369 224 384 232
rect 137 213 155 224
rect 118 205 155 213
rect 118 188 126 205
rect 143 188 155 205
rect -102 176 -87 184
rect -57 176 -42 184
rect -103 155 -85 176
rect -58 155 -40 176
rect 118 171 155 188
rect 182 179 200 224
rect 221 218 239 224
rect 266 220 284 224
rect 367 220 385 224
rect 221 203 245 218
rect 266 205 316 220
rect 367 205 428 220
rect 230 179 245 203
rect 301 181 316 205
rect -133 147 -85 155
rect -133 130 -125 147
rect -108 130 -85 147
rect -133 122 -85 130
rect -100 111 -85 122
rect -61 147 -10 155
rect -61 130 -35 147
rect -18 130 -10 147
rect -61 122 -10 130
rect 118 154 126 171
rect 143 154 155 171
rect 118 137 155 154
rect -61 111 -46 122
rect 118 120 126 137
rect 143 120 155 137
rect 118 112 155 120
rect 176 171 209 179
rect 176 154 184 171
rect 201 154 209 171
rect 176 137 209 154
rect 230 171 277 179
rect 230 154 252 171
rect 269 154 277 171
rect 230 146 277 154
rect 176 120 184 137
rect 201 120 209 137
rect 176 112 209 120
rect 140 101 155 112
rect 179 101 194 112
rect 262 101 277 146
rect 301 173 389 181
rect 301 166 364 173
rect 301 101 316 166
rect 356 156 364 166
rect 381 156 389 173
rect 356 148 389 156
rect 413 124 428 205
rect 616 274 631 287
rect 658 274 673 287
rect 616 224 631 232
rect 658 224 673 232
rect 711 224 726 232
rect 614 216 632 224
rect 599 208 632 216
rect 599 191 607 208
rect 624 191 632 208
rect 470 176 485 184
rect 515 176 530 184
rect 599 183 632 191
rect 656 184 674 224
rect 709 209 728 224
rect 1166 246 1181 254
rect 1205 246 1220 254
rect 468 168 486 176
rect 452 160 486 168
rect 513 167 531 176
rect 452 143 460 160
rect 477 143 486 160
rect 452 135 486 143
rect 507 159 567 167
rect 507 142 515 159
rect 532 142 567 159
rect 369 109 428 124
rect 468 123 483 135
rect 507 134 567 142
rect 552 123 567 134
rect 616 127 631 183
rect 655 176 688 184
rect 655 159 663 176
rect 680 159 688 176
rect 655 151 688 159
rect 369 101 384 109
rect 140 46 155 59
rect -778 24 -763 37
rect -100 24 -85 37
rect -61 24 -46 37
rect 179 25 194 59
rect 262 46 277 59
rect 301 46 316 59
rect 369 25 384 59
rect 616 112 688 127
rect 673 104 688 112
rect 709 104 724 209
rect 877 204 892 212
rect 919 204 934 212
rect 973 204 988 212
rect 1074 204 1089 212
rect 1113 204 1128 212
rect 799 187 832 195
rect 745 177 778 185
rect 745 160 753 177
rect 770 160 778 177
rect 745 152 778 160
rect 799 170 807 187
rect 824 170 832 187
rect 799 153 832 170
rect 755 104 770 152
rect 799 136 807 153
rect 824 143 832 153
rect 875 143 893 204
rect 824 136 893 143
rect 799 128 893 136
rect 917 195 935 204
rect 917 187 950 195
rect 917 170 925 187
rect 942 170 950 187
rect 917 153 950 170
rect 917 136 925 153
rect 942 136 950 153
rect 971 178 989 204
rect 1072 191 1090 204
rect 1032 183 1090 191
rect 971 170 1008 178
rect 971 153 983 170
rect 1000 153 1008 170
rect 971 145 1008 153
rect 1032 166 1065 183
rect 1082 166 1090 183
rect 1032 158 1090 166
rect 1111 175 1129 204
rect 1165 199 1183 246
rect 1204 238 1222 246
rect 1204 230 1237 238
rect 1204 213 1212 230
rect 1229 220 1237 230
rect 1229 213 1270 220
rect 1204 205 1270 213
rect 1111 167 1144 175
rect 917 128 950 136
rect 878 117 893 128
rect 921 117 936 128
rect 982 117 997 145
rect 1032 117 1047 158
rect 1111 150 1119 167
rect 1136 150 1144 167
rect 1111 142 1144 150
rect 1165 118 1180 199
rect 1201 151 1234 159
rect 1201 134 1209 151
rect 1226 134 1234 151
rect 1201 126 1234 134
rect 1079 103 1180 118
rect 1079 96 1094 103
rect 468 36 483 49
rect 179 10 384 25
rect 552 25 567 49
rect 673 49 688 62
rect 709 25 724 62
rect 755 49 770 62
rect 878 49 893 62
rect 921 49 936 62
rect 982 49 997 62
rect 1032 49 1047 62
rect 1204 83 1219 126
rect 1255 105 1270 205
rect 1620 296 1635 309
rect 1665 296 1680 309
rect 1502 263 1517 276
rect 1308 188 1323 196
rect 1359 188 1374 196
rect 1401 188 1416 196
rect 1502 192 1517 199
rect 1306 155 1324 188
rect 1357 155 1375 188
rect 1399 180 1417 188
rect 1500 183 1518 192
rect 1764 292 1779 305
rect 1817 296 1832 309
rect 1862 296 1877 309
rect 1764 184 1779 192
rect 2059 288 2074 301
rect 2104 288 2119 301
rect 2152 288 2167 301
rect 2199 288 2214 301
rect 2253 296 2268 309
rect 2300 296 2315 309
rect 2345 296 2360 309
rect 2390 296 2405 309
rect 2059 197 2074 204
rect 2104 197 2119 204
rect 2152 197 2167 204
rect 2199 197 2214 204
rect 1399 172 1432 180
rect 1399 155 1407 172
rect 1424 155 1432 172
rect 1291 147 1324 155
rect 1291 130 1299 147
rect 1316 130 1324 147
rect 1291 122 1324 130
rect 1345 147 1378 155
rect 1399 147 1432 155
rect 1490 175 1523 183
rect 1620 176 1635 184
rect 1665 176 1680 184
rect 1490 158 1498 175
rect 1515 158 1523 175
rect 1490 150 1523 158
rect 1345 130 1353 147
rect 1370 130 1378 147
rect 1345 122 1378 130
rect 1307 111 1322 122
rect 1359 111 1374 122
rect 1402 111 1417 147
rect 1508 132 1523 150
rect 1544 168 1577 176
rect 1544 151 1552 168
rect 1569 164 1577 168
rect 1618 164 1636 176
rect 1663 164 1681 176
rect 1763 165 1781 184
rect 1817 176 1832 184
rect 1862 176 1877 184
rect 1763 164 1778 165
rect 1569 151 1778 164
rect 1815 155 1833 176
rect 1860 155 1878 176
rect 1544 143 1778 151
rect 1611 135 1778 143
rect 1799 147 1878 155
rect 1243 90 1270 105
rect 1243 83 1258 90
rect 1079 25 1094 41
rect 1204 28 1219 41
rect 1243 28 1258 41
rect 552 10 1094 25
rect 1611 111 1626 135
rect 1654 111 1669 135
rect 1760 111 1775 135
rect 1799 130 1807 147
rect 1824 130 1878 147
rect 1799 122 1878 130
rect 2058 131 2076 197
rect 2103 191 2121 197
rect 2150 191 2168 197
rect 2103 170 2168 191
rect 2103 153 2130 170
rect 2147 153 2168 170
rect 2198 167 2216 197
rect 2253 176 2268 184
rect 2300 176 2315 184
rect 2345 176 2360 184
rect 2390 176 2405 184
rect 2251 167 2269 176
rect 2298 167 2316 176
rect 2343 167 2361 176
rect 2388 167 2406 176
rect 2103 145 2168 153
rect 2189 159 2222 167
rect 2058 123 2073 131
rect 2103 123 2118 145
rect 2150 123 2165 145
rect 2189 142 2197 159
rect 2214 142 2222 159
rect 2189 134 2222 142
rect 2246 159 2406 167
rect 2246 142 2254 159
rect 2271 142 2288 159
rect 2305 142 2322 159
rect 2339 142 2406 159
rect 2246 134 2406 142
rect 2196 123 2211 134
rect 2247 123 2262 134
rect 2305 123 2320 134
rect 2348 123 2363 134
rect 2391 123 2406 134
rect 1820 111 1835 122
rect 1863 111 1878 122
rect 1508 77 1523 90
rect 1307 24 1322 37
rect 1359 24 1374 37
rect 1402 24 1417 37
rect 1611 24 1626 37
rect 1654 24 1669 37
rect 1760 34 1775 47
rect 1820 24 1835 37
rect 1863 24 1878 37
rect 2058 25 2073 59
rect 2103 46 2118 59
rect 2150 46 2165 59
rect 2196 25 2211 59
rect 2247 36 2262 49
rect 2305 36 2320 49
rect 2348 36 2363 49
rect 2391 36 2406 49
rect 2058 10 2211 25
rect -680 -138 -647 -105
rect -671 -149 -656 -138
rect -671 -360 -656 -349
rect -680 -368 -647 -360
rect -680 -385 -672 -368
rect -655 -385 -647 -368
rect -680 -393 -647 -385
rect -680 -495 -647 -462
rect -671 -506 -656 -495
rect -671 -717 -656 -706
rect -680 -725 -647 -717
rect -680 -742 -672 -725
rect -655 -742 -647 -725
rect -680 -750 -647 -742
<< polycont >>
rect -847 1500 -830 1517
rect -847 1143 -830 1160
rect -456 1500 -439 1517
rect -456 1143 -439 1160
rect -1417 804 -1400 821
rect -1383 804 -1366 821
rect -701 796 -684 813
rect -611 796 -594 813
rect -527 799 -510 816
rect -453 799 -436 816
rect -393 799 -376 816
rect -332 799 -315 816
rect 145 799 162 816
rect 218 799 235 816
rect 279 799 296 816
rect 339 799 356 816
rect 481 799 498 816
rect 554 799 571 816
rect 615 799 632 816
rect 675 799 692 816
rect 817 799 834 816
rect 890 799 907 816
rect 951 799 968 816
rect 1011 799 1028 816
rect 1153 799 1170 816
rect 1226 799 1243 816
rect 1287 799 1304 816
rect 1347 799 1364 816
rect 1489 799 1506 816
rect 1562 799 1579 816
rect 1623 799 1640 816
rect 1683 799 1700 816
rect 1825 799 1842 816
rect 1898 799 1915 816
rect 1959 799 1976 816
rect 2019 799 2036 816
rect 2161 799 2178 816
rect 2234 799 2251 816
rect -1417 511 -1400 528
rect -1383 511 -1366 528
rect -701 519 -684 536
rect -611 519 -594 536
rect -517 506 -500 523
rect -433 519 -416 536
rect -379 519 -362 536
rect -322 519 -305 536
rect -265 509 -248 526
rect -211 511 -194 528
rect -125 511 -108 528
rect 126 528 143 545
rect 126 494 143 511
rect 184 528 201 545
rect 184 494 201 511
rect 252 495 269 512
rect 364 493 381 510
rect 126 460 143 477
rect 460 506 477 523
rect 515 507 532 524
rect 663 490 680 507
rect 607 458 624 475
rect 753 488 770 505
rect 807 512 824 529
rect 807 478 824 495
rect 925 512 942 529
rect 925 478 942 495
rect 983 496 1000 513
rect 1065 483 1082 500
rect 1119 498 1136 515
rect 1209 514 1226 531
rect 1299 519 1316 536
rect 1353 519 1370 536
rect 1407 494 1424 511
rect 1498 490 1515 507
rect 1552 498 1569 515
rect 1807 519 1824 536
rect 1212 436 1229 453
rect 2075 506 2092 523
rect 2109 506 2126 523
rect 2143 506 2160 523
rect 2177 506 2194 523
rect 2268 506 2285 523
rect 2302 506 2319 523
rect 2336 506 2353 523
rect 2370 506 2387 523
rect -841 138 -824 155
rect -807 138 -790 155
rect 126 188 143 205
rect -125 130 -108 147
rect -35 130 -18 147
rect 126 154 143 171
rect 126 120 143 137
rect 184 154 201 171
rect 252 154 269 171
rect 184 120 201 137
rect 364 156 381 173
rect 607 191 624 208
rect 460 143 477 160
rect 515 142 532 159
rect 663 159 680 176
rect 753 160 770 177
rect 807 170 824 187
rect 807 136 824 153
rect 925 170 942 187
rect 925 136 942 153
rect 983 153 1000 170
rect 1065 166 1082 183
rect 1212 213 1229 230
rect 1119 150 1136 167
rect 1209 134 1226 151
rect 1407 155 1424 172
rect 1299 130 1316 147
rect 1498 158 1515 175
rect 1353 130 1370 147
rect 1552 151 1569 168
rect 1807 130 1824 147
rect 2130 153 2147 170
rect 2197 142 2214 159
rect 2254 142 2271 159
rect 2288 142 2305 159
rect 2322 142 2339 159
rect -672 -385 -655 -368
rect -672 -742 -655 -725
<< xpolycontact >>
rect -1258 733 -1042 874
rect -992 733 -776 874
rect -1258 457 -1042 598
rect -992 457 -776 598
rect -682 67 -466 208
rect -416 67 -200 208
<< xpolyres >>
rect -1042 733 -992 874
rect -1042 457 -992 598
rect -466 67 -416 208
<< locali >>
rect -926 1806 -878 1823
rect -799 1806 -734 1823
rect -926 1775 -909 1806
rect -768 1775 -734 1806
rect -869 1730 -852 1738
rect -869 1534 -852 1542
rect -825 1730 -808 1738
rect -825 1534 -808 1542
rect -855 1500 -847 1517
rect -830 1500 -822 1517
rect -926 1466 -909 1497
rect -751 1497 -734 1775
rect -768 1466 -734 1497
rect -926 1449 -878 1466
rect -799 1449 -734 1466
rect -926 1418 -909 1449
rect -768 1418 -734 1449
rect -869 1373 -852 1381
rect -869 1177 -852 1185
rect -825 1373 -808 1381
rect -825 1177 -808 1185
rect -855 1143 -847 1160
rect -830 1143 -822 1160
rect -926 1109 -909 1140
rect -751 1140 -734 1418
rect -768 1109 -734 1140
rect -926 1092 -878 1109
rect -799 1092 -734 1109
rect -552 1806 -487 1823
rect -408 1806 -360 1823
rect -552 1775 -518 1806
rect -552 1497 -535 1775
rect -377 1775 -360 1806
rect -478 1730 -461 1738
rect -478 1534 -461 1542
rect -434 1730 -417 1738
rect -434 1534 -417 1542
rect -464 1500 -456 1517
rect -439 1500 -431 1517
rect -552 1466 -518 1497
rect -377 1466 -360 1497
rect -552 1449 -487 1466
rect -408 1449 -360 1466
rect -552 1418 -518 1449
rect -552 1140 -535 1418
rect -377 1418 -360 1449
rect -478 1373 -461 1381
rect -478 1177 -461 1185
rect -434 1373 -417 1381
rect -434 1177 -417 1185
rect -464 1143 -456 1160
rect -439 1143 -431 1160
rect -552 1109 -518 1140
rect -377 1109 -360 1140
rect -552 1092 -487 1109
rect -408 1092 -360 1109
rect -1440 990 -1424 1007
rect -1407 990 -1376 1007
rect -1359 990 -1328 1007
rect -1311 990 -1280 1007
rect -1263 990 -1232 1007
rect -1215 990 -1184 1007
rect -1167 990 -1136 1007
rect -1119 990 -1088 1007
rect -1071 990 -1040 1007
rect -1023 990 -992 1007
rect -975 990 -944 1007
rect -927 990 -896 1007
rect -879 990 -848 1007
rect -831 990 -800 1007
rect -783 990 -752 1007
rect -735 990 -704 1007
rect -687 990 -656 1007
rect -639 990 -608 1007
rect -591 990 -560 1007
rect -543 990 -512 1007
rect -495 990 -464 1007
rect -447 990 -416 1007
rect -399 990 -368 1007
rect -351 990 -320 1007
rect -303 990 -272 1007
rect -255 990 -224 1007
rect -207 990 -176 1007
rect -159 990 -128 1007
rect -111 990 -80 1007
rect -63 990 -32 1007
rect -15 990 15 1007
rect 32 990 63 1007
rect 80 990 111 1007
rect 128 990 159 1007
rect 176 990 207 1007
rect 224 990 255 1007
rect 272 990 303 1007
rect 320 990 351 1007
rect 368 990 399 1007
rect 416 990 447 1007
rect 464 990 495 1007
rect 512 990 543 1007
rect 560 990 591 1007
rect 608 990 639 1007
rect 656 990 687 1007
rect 704 990 735 1007
rect 752 990 783 1007
rect 800 990 831 1007
rect 848 990 879 1007
rect 896 990 927 1007
rect 944 990 975 1007
rect 992 990 1023 1007
rect 1040 990 1071 1007
rect 1088 990 1119 1007
rect 1136 990 1167 1007
rect 1184 990 1215 1007
rect 1232 990 1263 1007
rect 1280 990 1311 1007
rect 1328 990 1359 1007
rect 1376 990 1407 1007
rect 1424 990 1455 1007
rect 1472 990 1503 1007
rect 1520 990 1551 1007
rect 1568 990 1599 1007
rect 1616 990 1647 1007
rect 1664 990 1695 1007
rect 1712 990 1743 1007
rect 1760 990 1791 1007
rect 1808 990 1839 1007
rect 1856 990 1887 1007
rect 1904 990 1935 1007
rect 1952 990 1983 1007
rect 2000 990 2031 1007
rect 2048 990 2079 1007
rect 2096 990 2127 1007
rect 2144 990 2175 1007
rect 2192 990 2223 1007
rect 2240 990 2271 1007
rect 2288 990 2319 1007
rect 2336 990 2367 1007
rect 2384 990 2415 1007
rect 2432 990 2448 1007
rect -1391 956 -1358 990
rect -1391 939 -1383 956
rect -1366 939 -1358 956
rect -1391 921 -1358 939
rect -1391 904 -1383 921
rect -1366 904 -1358 921
rect -1391 886 -1358 904
rect -1391 869 -1383 886
rect -1366 869 -1358 886
rect -1391 861 -1358 869
rect -1341 956 -1308 964
rect -1341 939 -1333 956
rect -1316 939 -1308 956
rect -1341 914 -1308 939
rect -1341 897 -1333 914
rect -1316 897 -1308 914
rect -1341 873 -1308 897
rect -709 956 -676 990
rect -709 939 -701 956
rect -684 939 -676 956
rect -709 914 -676 939
rect -709 897 -701 914
rect -684 897 -676 914
rect -1341 856 -1333 873
rect -1316 856 -1308 873
rect -1427 821 -1358 844
rect -1427 804 -1419 821
rect -1400 804 -1383 821
rect -1366 804 -1358 821
rect -1427 796 -1358 804
rect -1341 829 -1308 856
rect -1341 800 -1258 829
rect -1391 771 -1358 779
rect -1391 754 -1383 771
rect -1366 754 -1358 771
rect -1391 726 -1358 754
rect -1391 709 -1383 726
rect -1366 709 -1358 726
rect -1391 674 -1358 709
rect -1341 771 -1308 800
rect -1341 754 -1333 771
rect -1316 754 -1308 771
rect -1341 726 -1308 754
rect -709 873 -676 897
rect -709 856 -701 873
rect -684 856 -676 873
rect -709 848 -676 856
rect -659 956 -636 964
rect -659 939 -656 956
rect -639 939 -636 956
rect -659 914 -636 939
rect -659 897 -656 914
rect -639 897 -636 914
rect -659 873 -636 897
rect -659 856 -656 873
rect -639 856 -636 873
rect -776 813 -676 821
rect -776 796 -701 813
rect -684 796 -676 813
rect -776 788 -676 796
rect -709 784 -676 788
rect -659 784 -636 856
rect -619 956 -586 990
rect -619 939 -611 956
rect -594 939 -586 956
rect -619 914 -586 939
rect -619 897 -611 914
rect -594 897 -586 914
rect -619 873 -586 897
rect -619 856 -611 873
rect -594 856 -586 873
rect -566 956 -533 990
rect -566 939 -558 956
rect -541 939 -533 956
rect -566 920 -533 939
rect -566 903 -558 920
rect -541 903 -533 920
rect -566 885 -533 903
rect -566 868 -558 885
rect -541 868 -533 885
rect -566 859 -533 868
rect -461 956 -368 990
rect -461 939 -429 956
rect -412 939 -368 956
rect -461 920 -368 939
rect -461 903 -429 920
rect -412 903 -368 920
rect -461 885 -368 903
rect -461 868 -429 885
rect -412 868 -368 885
rect -619 848 -586 856
rect -619 813 -586 821
rect -619 796 -611 813
rect -594 796 -586 813
rect -619 784 -586 796
rect -559 816 -502 824
rect -559 799 -527 816
rect -510 799 -502 816
rect -653 767 -636 784
rect -707 750 -699 767
rect -682 750 -674 767
rect -653 750 -617 767
rect -600 750 -592 767
rect -1341 709 -1333 726
rect -1316 709 -1308 726
rect -1341 701 -1308 709
rect -707 726 -674 750
rect -707 709 -699 726
rect -682 709 -674 726
rect -707 674 -674 709
rect -625 729 -592 750
rect -625 726 -616 729
rect -625 709 -617 726
rect -599 712 -592 729
rect -600 709 -592 712
rect -625 701 -592 709
rect -559 738 -502 799
rect -461 816 -368 868
rect -310 956 -277 990
rect -310 939 -302 956
rect -285 939 -277 956
rect -310 920 -277 939
rect -310 903 -302 920
rect -285 903 -277 920
rect -310 885 -277 903
rect 9 955 87 972
rect 9 938 15 955
rect 32 938 63 955
rect 9 935 63 938
rect 80 935 87 955
rect 9 912 87 935
rect 9 895 15 912
rect 32 895 63 912
rect 80 895 87 912
rect 9 887 87 895
rect 105 956 138 990
rect 105 939 113 956
rect 130 939 138 956
rect 105 920 138 939
rect 105 903 113 920
rect 130 903 138 920
rect -310 868 -302 885
rect -285 868 -277 885
rect -310 860 -277 868
rect 105 885 138 903
rect 105 868 113 885
rect 130 868 138 885
rect 105 859 138 868
rect 210 956 304 990
rect 210 939 242 956
rect 259 939 304 956
rect 210 920 304 939
rect 210 903 242 920
rect 259 903 304 920
rect 210 885 304 903
rect 210 868 242 885
rect 259 868 304 885
rect -461 799 -453 816
rect -436 799 -393 816
rect -376 799 -368 816
rect -461 791 -368 799
rect -340 816 -270 824
rect -340 799 -332 816
rect -315 799 -270 816
rect -559 721 -551 738
rect -534 721 -502 738
rect -559 674 -502 721
rect -431 738 -398 746
rect -431 721 -423 738
rect -406 721 -398 738
rect -431 674 -398 721
rect -340 738 -270 799
rect 113 816 170 824
rect 113 799 145 816
rect 162 799 170 816
rect -340 721 -295 738
rect -278 721 -270 738
rect -340 674 -270 721
rect 9 768 87 776
rect 9 751 15 768
rect 32 751 63 768
rect 80 751 87 768
rect 9 730 87 751
rect 9 710 15 730
rect 32 727 87 730
rect 32 710 63 727
rect 80 710 87 727
rect 9 692 87 710
rect 113 738 170 799
rect 210 816 304 868
rect 362 956 395 990
rect 362 939 370 956
rect 387 939 395 956
rect 362 920 395 939
rect 362 903 370 920
rect 387 903 395 920
rect 362 885 395 903
rect 362 868 370 885
rect 387 868 395 885
rect 362 860 395 868
rect 441 956 474 990
rect 441 939 449 956
rect 466 939 474 956
rect 441 920 474 939
rect 441 903 449 920
rect 466 903 474 920
rect 441 885 474 903
rect 441 868 449 885
rect 466 868 474 885
rect 441 859 474 868
rect 546 956 640 990
rect 546 939 578 956
rect 595 939 640 956
rect 546 920 640 939
rect 546 903 578 920
rect 595 903 640 920
rect 546 885 640 903
rect 546 868 578 885
rect 595 868 640 885
rect 210 799 218 816
rect 235 799 279 816
rect 296 799 304 816
rect 210 791 304 799
rect 331 816 401 824
rect 331 799 339 816
rect 356 799 401 816
rect 113 721 121 738
rect 138 721 170 738
rect 113 674 170 721
rect 241 738 274 746
rect 241 721 249 738
rect 266 721 274 738
rect 241 674 274 721
rect 331 738 401 799
rect 331 721 377 738
rect 394 721 401 738
rect 331 674 401 721
rect 449 816 506 824
rect 449 799 481 816
rect 498 799 506 816
rect 449 738 506 799
rect 546 816 640 868
rect 698 956 731 990
rect 698 939 706 956
rect 723 939 731 956
rect 698 920 731 939
rect 698 903 706 920
rect 723 903 731 920
rect 698 885 731 903
rect 698 868 706 885
rect 723 868 731 885
rect 698 860 731 868
rect 777 956 810 990
rect 777 939 785 956
rect 802 939 810 956
rect 777 920 810 939
rect 777 903 785 920
rect 802 903 810 920
rect 777 885 810 903
rect 777 868 785 885
rect 802 868 810 885
rect 777 859 810 868
rect 882 956 976 990
rect 882 939 914 956
rect 931 939 976 956
rect 882 920 976 939
rect 882 903 914 920
rect 931 903 976 920
rect 882 885 976 903
rect 882 868 914 885
rect 931 868 976 885
rect 546 799 554 816
rect 571 799 615 816
rect 632 799 640 816
rect 546 791 640 799
rect 667 816 737 824
rect 667 799 675 816
rect 692 799 737 816
rect 449 721 457 738
rect 474 721 506 738
rect 449 674 506 721
rect 577 738 610 746
rect 577 721 585 738
rect 602 721 610 738
rect 577 674 610 721
rect 667 738 737 799
rect 667 721 713 738
rect 730 721 737 738
rect 667 674 737 721
rect 785 816 842 824
rect 785 799 817 816
rect 834 799 842 816
rect 785 738 842 799
rect 882 816 976 868
rect 1034 956 1067 990
rect 1034 939 1042 956
rect 1059 939 1067 956
rect 1034 920 1067 939
rect 1034 903 1042 920
rect 1059 903 1067 920
rect 1034 885 1067 903
rect 1034 868 1042 885
rect 1059 868 1067 885
rect 1034 860 1067 868
rect 1113 956 1146 990
rect 1113 939 1121 956
rect 1138 939 1146 956
rect 1113 920 1146 939
rect 1113 903 1121 920
rect 1138 903 1146 920
rect 1113 885 1146 903
rect 1113 868 1121 885
rect 1138 868 1146 885
rect 1113 859 1146 868
rect 1218 956 1312 990
rect 1218 939 1250 956
rect 1267 939 1312 956
rect 1218 920 1312 939
rect 1218 903 1250 920
rect 1267 903 1312 920
rect 1218 885 1312 903
rect 1218 868 1250 885
rect 1267 868 1312 885
rect 882 799 890 816
rect 907 799 951 816
rect 968 799 976 816
rect 882 791 976 799
rect 1003 816 1073 824
rect 1003 799 1011 816
rect 1028 799 1073 816
rect 785 721 793 738
rect 810 721 842 738
rect 785 674 842 721
rect 913 738 946 746
rect 913 721 921 738
rect 938 721 946 738
rect 913 674 946 721
rect 1003 738 1073 799
rect 1003 721 1049 738
rect 1066 721 1073 738
rect 1003 674 1073 721
rect 1121 816 1178 824
rect 1121 799 1153 816
rect 1170 799 1178 816
rect 1121 738 1178 799
rect 1218 816 1312 868
rect 1370 956 1403 990
rect 1370 939 1378 956
rect 1395 939 1403 956
rect 1370 920 1403 939
rect 1370 903 1378 920
rect 1395 903 1403 920
rect 1370 885 1403 903
rect 1370 868 1378 885
rect 1395 868 1403 885
rect 1370 860 1403 868
rect 1449 956 1482 990
rect 1449 939 1457 956
rect 1474 939 1482 956
rect 1449 920 1482 939
rect 1449 903 1457 920
rect 1474 903 1482 920
rect 1449 885 1482 903
rect 1449 868 1457 885
rect 1474 868 1482 885
rect 1449 859 1482 868
rect 1554 956 1648 990
rect 1554 939 1586 956
rect 1603 939 1648 956
rect 1554 920 1648 939
rect 1554 903 1586 920
rect 1603 903 1648 920
rect 1554 885 1648 903
rect 1554 868 1586 885
rect 1603 868 1648 885
rect 1218 799 1226 816
rect 1243 799 1287 816
rect 1304 799 1312 816
rect 1218 791 1312 799
rect 1339 816 1409 824
rect 1339 799 1347 816
rect 1364 799 1409 816
rect 1121 721 1129 738
rect 1146 721 1178 738
rect 1121 674 1178 721
rect 1249 738 1282 746
rect 1249 721 1257 738
rect 1274 721 1282 738
rect 1249 674 1282 721
rect 1339 738 1409 799
rect 1339 721 1385 738
rect 1402 721 1409 738
rect 1339 674 1409 721
rect 1457 816 1514 824
rect 1457 799 1489 816
rect 1506 799 1514 816
rect 1457 738 1514 799
rect 1554 816 1648 868
rect 1706 956 1739 990
rect 1706 939 1714 956
rect 1731 939 1739 956
rect 1706 920 1739 939
rect 1706 903 1714 920
rect 1731 903 1739 920
rect 1706 885 1739 903
rect 1706 868 1714 885
rect 1731 868 1739 885
rect 1706 860 1739 868
rect 1785 956 1818 990
rect 1785 939 1793 956
rect 1810 939 1818 956
rect 1785 920 1818 939
rect 1785 903 1793 920
rect 1810 903 1818 920
rect 1785 885 1818 903
rect 1785 868 1793 885
rect 1810 868 1818 885
rect 1785 859 1818 868
rect 1890 956 1984 990
rect 1890 939 1922 956
rect 1939 939 1984 956
rect 1890 920 1984 939
rect 1890 903 1922 920
rect 1939 903 1984 920
rect 1890 885 1984 903
rect 1890 868 1922 885
rect 1939 868 1984 885
rect 1554 799 1562 816
rect 1579 799 1623 816
rect 1640 799 1648 816
rect 1554 791 1648 799
rect 1675 816 1745 824
rect 1675 799 1683 816
rect 1700 799 1745 816
rect 1457 721 1465 738
rect 1482 721 1514 738
rect 1457 674 1514 721
rect 1585 738 1618 746
rect 1585 721 1593 738
rect 1610 721 1618 738
rect 1585 674 1618 721
rect 1675 738 1745 799
rect 1675 721 1721 738
rect 1738 721 1745 738
rect 1675 674 1745 721
rect 1793 816 1850 824
rect 1793 799 1825 816
rect 1842 799 1850 816
rect 1793 738 1850 799
rect 1890 816 1984 868
rect 2042 956 2075 990
rect 2042 939 2050 956
rect 2067 939 2075 956
rect 2042 920 2075 939
rect 2042 903 2050 920
rect 2067 903 2075 920
rect 2042 885 2075 903
rect 2042 868 2050 885
rect 2067 868 2075 885
rect 2042 860 2075 868
rect 2121 956 2154 990
rect 2121 939 2129 956
rect 2146 939 2154 956
rect 2121 920 2154 939
rect 2121 903 2129 920
rect 2146 903 2154 920
rect 2121 885 2154 903
rect 2121 868 2129 885
rect 2146 868 2154 885
rect 2121 859 2154 868
rect 2226 956 2283 990
rect 2226 939 2258 956
rect 2275 939 2283 956
rect 2226 920 2283 939
rect 2226 903 2258 920
rect 2275 903 2283 920
rect 2226 885 2283 903
rect 2226 868 2258 885
rect 2275 868 2283 885
rect 1890 799 1898 816
rect 1915 799 1959 816
rect 1976 799 1984 816
rect 1890 791 1984 799
rect 2011 816 2081 824
rect 2011 799 2019 816
rect 2036 799 2081 816
rect 1793 721 1801 738
rect 1818 721 1850 738
rect 1793 674 1850 721
rect 1921 738 1954 746
rect 1921 721 1929 738
rect 1946 721 1954 738
rect 1921 674 1954 721
rect 2011 738 2081 799
rect 2011 721 2057 738
rect 2074 721 2081 738
rect 2011 674 2081 721
rect 2129 816 2186 824
rect 2129 799 2161 816
rect 2178 799 2186 816
rect 2129 738 2186 799
rect 2226 816 2283 868
rect 2226 799 2234 816
rect 2251 799 2283 816
rect 2226 791 2283 799
rect 2129 721 2137 738
rect 2154 721 2186 738
rect 2129 674 2186 721
rect 2257 738 2290 746
rect 2257 721 2265 738
rect 2282 721 2290 738
rect 2257 674 2290 721
rect -1440 657 -1424 674
rect -1407 657 -1376 674
rect -1359 657 -1328 674
rect -1311 657 -1280 674
rect -1263 657 -1232 674
rect -1215 657 -1184 674
rect -1167 657 -1136 674
rect -1119 657 -1088 674
rect -1071 657 -1040 674
rect -1023 657 -992 674
rect -975 657 -944 674
rect -927 657 -896 674
rect -879 657 -848 674
rect -831 657 -800 674
rect -783 657 -752 674
rect -735 657 -704 674
rect -687 657 -656 674
rect -639 657 -608 674
rect -591 657 -560 674
rect -543 657 -512 674
rect -495 657 -464 674
rect -447 657 -416 674
rect -399 657 -368 674
rect -351 657 -320 674
rect -303 657 -272 674
rect -255 657 -224 674
rect -207 657 -176 674
rect -159 657 -128 674
rect -111 657 -80 674
rect -63 657 -32 674
rect -15 657 15 674
rect 32 657 63 674
rect 80 657 111 674
rect 128 657 159 674
rect 176 657 207 674
rect 224 657 255 674
rect 272 657 303 674
rect 320 657 351 674
rect 368 657 399 674
rect 416 657 447 674
rect 464 657 495 674
rect 512 657 543 674
rect 560 657 591 674
rect 608 657 639 674
rect 656 657 687 674
rect 704 657 735 674
rect 752 657 783 674
rect 800 657 831 674
rect 848 657 879 674
rect 896 657 927 674
rect 944 657 975 674
rect 992 657 1023 674
rect 1040 657 1071 674
rect 1088 657 1119 674
rect 1136 657 1167 674
rect 1184 657 1215 674
rect 1232 657 1263 674
rect 1280 657 1311 674
rect 1328 657 1359 674
rect 1376 657 1407 674
rect 1424 657 1455 674
rect 1472 657 1503 674
rect 1520 657 1551 674
rect 1568 657 1599 674
rect 1616 657 1647 674
rect 1664 657 1695 674
rect 1712 657 1743 674
rect 1760 657 1791 674
rect 1808 657 1839 674
rect 1856 657 1887 674
rect 1904 657 1935 674
rect 1952 657 1983 674
rect 2000 657 2031 674
rect 2048 657 2079 674
rect 2096 657 2127 674
rect 2144 657 2175 674
rect 2192 657 2223 674
rect 2240 657 2271 674
rect 2288 657 2319 674
rect 2336 657 2367 674
rect 2384 657 2415 674
rect 2432 657 2448 674
rect -1391 623 -1358 657
rect -1391 606 -1383 623
rect -1366 606 -1358 623
rect -1391 578 -1358 606
rect -1391 561 -1383 578
rect -1366 561 -1358 578
rect -1391 553 -1358 561
rect -1341 623 -1308 631
rect -1341 606 -1333 623
rect -1316 606 -1308 623
rect -1341 578 -1308 606
rect -707 623 -674 657
rect -707 606 -699 623
rect -682 606 -674 623
rect -1341 561 -1333 578
rect -1316 561 -1308 578
rect -1427 528 -1358 536
rect -1427 511 -1419 528
rect -1400 511 -1383 528
rect -1366 511 -1358 528
rect -1427 488 -1358 511
rect -1341 532 -1308 561
rect -1341 502 -1258 532
rect -1341 476 -1308 502
rect -1391 463 -1358 471
rect -1391 446 -1383 463
rect -1366 446 -1358 463
rect -1391 428 -1358 446
rect -1391 411 -1383 428
rect -1366 411 -1358 428
rect -1391 393 -1358 411
rect -1391 376 -1383 393
rect -1366 376 -1358 393
rect -1391 341 -1358 376
rect -1341 459 -1333 476
rect -1316 459 -1308 476
rect -1341 434 -1308 459
rect -707 582 -674 606
rect -625 623 -592 631
rect -625 606 -617 623
rect -600 620 -592 623
rect -625 603 -616 606
rect -599 603 -592 620
rect -513 623 -475 657
rect -625 582 -592 603
rect -707 565 -699 582
rect -682 565 -674 582
rect -653 565 -617 582
rect -600 565 -592 582
rect -564 591 -531 612
rect -564 574 -556 591
rect -539 574 -531 591
rect -653 548 -636 565
rect -564 553 -531 574
rect -513 606 -503 623
rect -486 606 -475 623
rect -513 598 -475 606
rect -458 619 -263 627
rect -458 602 -405 619
rect -388 602 -263 619
rect -513 578 -492 598
rect -458 581 -441 602
rect -513 561 -512 578
rect -495 561 -492 578
rect -513 553 -492 561
rect -475 564 -441 581
rect -424 568 -297 585
rect -709 544 -676 548
rect -776 536 -676 544
rect -776 519 -701 536
rect -684 519 -676 536
rect -776 511 -676 519
rect -709 476 -676 484
rect -709 459 -701 476
rect -684 459 -676 476
rect -1341 417 -1333 434
rect -1316 417 -1308 434
rect -1341 393 -1308 417
rect -1341 376 -1333 393
rect -1316 376 -1308 393
rect -1341 368 -1308 376
rect -709 434 -676 459
rect -709 417 -701 434
rect -684 417 -676 434
rect -709 393 -676 417
rect -709 376 -701 393
rect -684 376 -676 393
rect -709 341 -676 376
rect -659 476 -636 548
rect -619 536 -586 548
rect -619 519 -611 536
rect -594 519 -586 536
rect -619 511 -586 519
rect -659 459 -656 476
rect -639 459 -636 476
rect -659 434 -636 459
rect -659 417 -656 434
rect -639 417 -636 434
rect -659 393 -636 417
rect -659 376 -656 393
rect -639 376 -636 393
rect -659 368 -636 376
rect -619 476 -586 484
rect -619 459 -611 476
rect -594 459 -586 476
rect -619 434 -586 459
rect -619 417 -611 434
rect -594 417 -586 434
rect -619 393 -586 417
rect -564 471 -547 553
rect -525 524 -492 531
rect -525 507 -518 524
rect -501 523 -492 524
rect -525 506 -517 507
rect -500 506 -492 523
rect -525 488 -492 506
rect -475 494 -458 564
rect -424 544 -407 568
rect -441 536 -407 544
rect -441 519 -433 536
rect -416 519 -407 536
rect -441 511 -407 519
rect -387 536 -348 548
rect -387 519 -379 536
rect -362 519 -348 536
rect -387 511 -348 519
rect -330 537 -297 568
rect -280 568 -263 602
rect -246 610 -213 657
rect -246 593 -238 610
rect -221 593 -213 610
rect -246 585 -213 593
rect -189 623 -152 631
rect -189 606 -181 623
rect -164 606 -152 623
rect -189 578 -152 606
rect -280 551 -206 568
rect -189 561 -181 578
rect -164 561 -152 578
rect -189 553 -152 561
rect -131 623 -106 657
rect -131 606 -123 623
rect -131 578 -106 606
rect -131 561 -123 578
rect -131 553 -106 561
rect -88 623 -55 631
rect -88 606 -80 623
rect -63 606 -55 623
rect -88 578 -55 606
rect -88 561 -80 578
rect -63 561 -55 578
rect -88 553 -55 561
rect -37 623 -12 657
rect -20 606 -12 623
rect -37 578 -12 606
rect -20 561 -12 578
rect -37 553 -12 561
rect 9 622 87 639
rect 9 602 15 622
rect 32 605 63 622
rect 80 605 87 622
rect 32 602 87 605
rect 9 580 87 602
rect 9 563 15 580
rect 32 563 63 580
rect 80 563 87 580
rect 9 555 87 563
rect 110 598 143 657
rect 110 581 118 598
rect 135 581 143 598
rect 110 570 143 581
rect 192 595 265 603
rect 192 578 200 595
rect 217 578 240 595
rect 257 578 265 595
rect 192 570 265 578
rect 314 598 339 657
rect 489 642 514 657
rect 314 581 322 598
rect 314 571 339 581
rect 356 623 449 640
rect 110 553 142 570
rect 244 554 265 570
rect 356 554 373 623
rect -330 519 -322 537
rect -305 519 -297 537
rect -223 536 -206 551
rect -330 511 -297 519
rect -280 526 -240 534
rect -280 509 -265 526
rect -248 509 -240 526
rect -280 501 -240 509
rect -223 528 -186 536
rect -223 511 -211 528
rect -194 511 -186 528
rect -223 503 -186 511
rect -475 477 -336 494
rect -369 476 -336 477
rect -564 468 -531 471
rect -564 451 -556 468
rect -539 460 -531 468
rect -539 451 -444 460
rect -564 443 -444 451
rect -564 421 -531 443
rect -564 404 -556 421
rect -539 404 -531 421
rect -564 396 -531 404
rect -511 423 -478 426
rect -511 406 -503 423
rect -486 406 -478 423
rect -619 376 -611 393
rect -594 376 -586 393
rect -619 341 -586 376
rect -511 341 -478 406
rect -461 375 -444 443
rect -369 459 -361 476
rect -344 459 -336 476
rect -369 417 -336 459
rect -369 400 -361 417
rect -344 400 -336 417
rect -369 392 -336 400
rect -280 375 -263 501
rect -169 484 -152 553
rect -133 530 -100 536
rect -133 513 -126 530
rect -109 528 -100 530
rect -133 511 -125 513
rect -108 511 -100 528
rect -133 488 -100 511
rect -461 358 -263 375
rect -246 476 -213 484
rect -246 459 -238 476
rect -221 459 -213 476
rect -246 434 -213 459
rect -246 417 -238 434
rect -221 417 -213 434
rect -246 393 -213 417
rect -246 376 -238 393
rect -221 376 -213 393
rect -246 341 -213 376
rect -196 476 -152 484
rect -196 459 -188 476
rect -171 459 -152 476
rect -83 476 -55 553
rect 108 545 227 553
rect 108 528 126 545
rect 143 528 184 545
rect 201 528 227 545
rect 244 537 373 554
rect 390 593 415 606
rect 407 576 415 593
rect 432 600 449 623
rect 489 625 497 642
rect 489 617 514 625
rect 531 623 624 640
rect 531 600 548 623
rect 432 583 548 600
rect 565 598 590 606
rect 108 520 227 528
rect 108 511 151 520
rect 108 494 126 511
rect 143 494 151 511
rect -196 443 -152 459
rect -196 434 -180 443
rect -196 417 -188 434
rect -163 426 -152 443
rect -171 417 -152 426
rect -196 393 -152 417
rect -196 376 -188 393
rect -171 376 -152 393
rect -196 368 -152 376
rect -133 463 -100 471
rect -133 446 -125 463
rect -108 446 -100 463
rect -133 428 -100 446
rect -133 411 -125 428
rect -108 411 -100 428
rect -133 393 -100 411
rect -133 376 -125 393
rect -108 376 -100 393
rect -133 341 -100 376
rect -83 459 -80 476
rect -63 459 -55 476
rect -83 434 -55 459
rect -83 417 -80 434
rect -63 417 -55 434
rect -83 407 -55 417
rect -83 393 -79 407
rect -83 376 -80 393
rect -62 390 -55 407
rect -63 376 -55 390
rect -83 368 -55 376
rect -35 476 -10 484
rect -18 459 -10 476
rect -35 434 -10 459
rect 108 477 151 494
rect 176 511 227 520
rect 176 494 184 511
rect 201 494 227 511
rect 176 486 227 494
rect 244 512 277 520
rect 244 495 252 512
rect 271 495 277 512
rect 244 487 277 495
rect 108 460 126 477
rect 143 460 151 477
rect 294 470 311 537
rect 390 518 415 576
rect 565 581 573 598
rect 438 549 446 566
rect 463 549 519 566
rect 502 532 519 549
rect 565 564 590 581
rect 607 582 624 623
rect 641 624 668 657
rect 641 607 642 624
rect 659 607 668 624
rect 641 599 668 607
rect 690 622 807 639
rect 690 582 707 622
rect 607 565 707 582
rect 724 591 757 605
rect 724 574 732 591
rect 749 574 757 591
rect 565 548 573 564
rect 557 547 573 548
rect 590 547 707 548
rect 557 545 707 547
rect 356 510 415 518
rect 356 493 364 510
rect 381 493 415 510
rect 356 485 415 493
rect 444 523 485 531
rect 444 506 458 523
rect 477 506 485 523
rect 444 488 485 506
rect 502 524 540 532
rect 502 507 515 524
rect 532 507 540 524
rect 502 499 540 507
rect 557 531 687 545
rect 108 452 151 460
rect 244 453 311 470
rect -18 417 -10 434
rect -35 393 -10 417
rect -18 376 -10 393
rect -35 341 -10 376
rect 9 437 87 445
rect 9 420 15 437
rect 32 420 63 437
rect 80 420 87 437
rect 244 436 261 453
rect 9 397 87 420
rect 9 394 63 397
rect 9 377 15 394
rect 32 377 63 394
rect 80 377 87 397
rect 9 359 87 377
rect 107 427 219 435
rect 107 410 115 427
rect 132 418 219 427
rect 107 393 132 410
rect 107 376 115 393
rect 107 368 132 376
rect 152 393 185 401
rect 152 376 160 393
rect 177 376 185 393
rect 152 341 185 376
rect 202 375 219 418
rect 236 423 261 436
rect 236 406 244 423
rect 236 392 261 406
rect 281 428 314 436
rect 281 411 289 428
rect 306 411 314 428
rect 281 393 314 411
rect 281 376 289 393
rect 306 376 314 393
rect 281 375 314 376
rect 202 358 314 375
rect 337 428 370 436
rect 337 411 345 428
rect 362 411 370 428
rect 337 393 370 411
rect 337 376 345 393
rect 362 376 370 393
rect 337 341 370 376
rect 390 428 415 485
rect 502 471 519 499
rect 557 482 574 531
rect 655 528 687 531
rect 704 528 707 545
rect 724 547 757 574
rect 774 593 807 622
rect 830 623 958 639
rect 830 606 843 623
rect 860 622 958 623
rect 860 606 873 622
rect 830 598 873 606
rect 941 605 958 622
rect 774 576 782 593
rect 799 581 807 593
rect 891 588 924 605
rect 799 576 866 581
rect 774 564 866 576
rect 891 571 899 588
rect 916 571 924 588
rect 941 597 984 605
rect 941 580 954 597
rect 971 580 984 597
rect 941 572 984 580
rect 1001 597 1034 657
rect 1264 640 1301 657
rect 1001 580 1009 597
rect 1026 580 1034 597
rect 1001 572 1034 580
rect 1051 623 1247 640
rect 1264 623 1274 640
rect 1291 623 1301 640
rect 1319 633 1455 640
rect 1319 623 1430 633
rect 724 530 832 547
rect 655 513 707 528
rect 799 529 832 530
rect 655 507 778 513
rect 655 490 663 507
rect 680 505 778 507
rect 680 490 753 505
rect 655 488 753 490
rect 770 488 778 505
rect 407 411 415 428
rect 390 393 415 411
rect 407 376 415 393
rect 390 368 415 376
rect 438 463 519 471
rect 438 446 446 463
rect 463 454 519 463
rect 536 474 574 482
rect 553 457 574 474
rect 438 428 463 446
rect 438 411 446 428
rect 438 393 463 411
rect 438 376 446 393
rect 438 368 463 376
rect 483 432 516 437
rect 483 415 491 432
rect 508 415 516 432
rect 483 393 516 415
rect 483 376 491 393
rect 508 376 516 393
rect 483 341 516 376
rect 536 433 574 457
rect 599 475 632 483
rect 655 482 778 488
rect 745 480 778 482
rect 799 512 807 529
rect 824 512 832 529
rect 799 495 832 512
rect 599 458 607 475
rect 624 465 632 475
rect 799 478 807 495
rect 824 478 832 495
rect 624 458 651 465
rect 799 462 832 478
rect 599 448 651 458
rect 553 416 574 433
rect 536 393 574 416
rect 553 376 574 393
rect 536 368 574 376
rect 592 419 617 431
rect 609 402 617 419
rect 592 341 617 402
rect 634 375 651 448
rect 680 445 832 462
rect 680 423 713 445
rect 849 428 866 564
rect 680 406 688 423
rect 705 406 713 423
rect 680 392 713 406
rect 730 423 866 428
rect 730 406 738 423
rect 755 411 866 423
rect 883 554 924 571
rect 1051 555 1068 623
rect 1230 606 1247 623
rect 1319 606 1332 623
rect 1349 606 1361 623
rect 1422 616 1430 623
rect 1447 616 1455 633
rect 1578 623 1607 657
rect 1578 606 1589 623
rect 1606 606 1607 623
rect 1092 589 1100 606
rect 1117 589 1141 606
rect 1158 589 1182 606
rect 1199 589 1207 606
rect 1230 589 1302 606
rect 1379 599 1404 606
rect 1379 597 1545 599
rect 1092 581 1207 589
rect 1190 572 1207 581
rect 1285 572 1362 589
rect 1190 555 1268 572
rect 883 453 900 554
rect 941 538 1068 555
rect 1111 545 1144 548
rect 941 537 958 538
rect 917 529 958 537
rect 917 512 925 529
rect 942 512 958 529
rect 1111 528 1119 545
rect 1136 538 1144 545
rect 1136 531 1234 538
rect 1136 528 1209 531
rect 917 495 958 512
rect 917 478 925 495
rect 942 478 958 495
rect 975 513 1040 521
rect 975 496 983 513
rect 1000 508 1040 513
rect 1111 515 1209 528
rect 1000 496 1023 508
rect 975 491 1023 496
rect 975 488 1040 491
rect 1057 500 1090 508
rect 917 470 958 478
rect 1057 483 1065 500
rect 1082 483 1090 500
rect 1111 498 1119 515
rect 1136 514 1209 515
rect 1226 514 1234 531
rect 1136 508 1234 514
rect 1136 498 1144 508
rect 1111 490 1144 498
rect 1251 491 1268 555
rect 1345 553 1362 572
rect 1396 582 1545 597
rect 1396 580 1404 582
rect 1379 570 1404 580
rect 1528 565 1561 582
rect 1456 557 1511 565
rect 1456 553 1486 557
rect 1291 536 1328 548
rect 1291 519 1299 536
rect 1316 519 1328 536
rect 1291 508 1328 519
rect 1345 540 1486 553
rect 1503 540 1511 557
rect 1345 536 1511 540
rect 1345 519 1353 536
rect 1370 519 1378 536
rect 1456 532 1511 536
rect 1345 511 1378 519
rect 1399 511 1432 519
rect 1291 491 1311 508
rect 1399 494 1407 511
rect 1424 494 1432 511
rect 1057 471 1090 483
rect 986 454 1090 471
rect 1170 474 1271 491
rect 1345 477 1432 494
rect 1345 474 1362 477
rect 1170 456 1187 474
rect 1254 457 1362 474
rect 1456 465 1473 532
rect 1544 523 1561 565
rect 1578 578 1607 606
rect 1578 561 1589 578
rect 1606 561 1607 578
rect 1578 553 1607 561
rect 1624 623 1657 631
rect 1624 606 1632 623
rect 1649 606 1657 623
rect 1624 578 1657 606
rect 1624 561 1632 578
rect 1649 561 1657 578
rect 1624 544 1657 561
rect 1674 623 1707 657
rect 1674 606 1675 623
rect 1692 606 1707 623
rect 1783 623 1816 657
rect 1674 578 1707 606
rect 1674 561 1675 578
rect 1692 561 1707 578
rect 1674 553 1707 561
rect 1730 610 1763 612
rect 1730 593 1738 610
rect 1755 593 1763 610
rect 1730 576 1763 593
rect 1730 559 1738 576
rect 1755 559 1763 576
rect 1783 606 1791 623
rect 1808 606 1816 623
rect 1783 586 1816 606
rect 1783 569 1791 586
rect 1808 569 1816 586
rect 1783 561 1816 569
rect 1833 623 1866 631
rect 1833 606 1841 623
rect 1858 606 1866 623
rect 1833 586 1866 606
rect 1833 569 1841 586
rect 1858 569 1866 586
rect 1833 561 1866 569
rect 1544 515 1577 523
rect 1490 507 1523 515
rect 1490 490 1498 507
rect 1515 490 1523 507
rect 1490 482 1523 490
rect 1544 498 1552 515
rect 1569 498 1577 515
rect 1544 490 1577 498
rect 1633 511 1657 544
rect 1730 544 1763 559
rect 1730 536 1832 544
rect 1730 519 1807 536
rect 1824 519 1832 536
rect 1730 511 1832 519
rect 986 453 1019 454
rect 883 448 1019 453
rect 883 436 994 448
rect 755 406 763 411
rect 730 392 763 406
rect 883 393 900 436
rect 986 431 994 436
rect 1011 431 1019 448
rect 1126 448 1187 456
rect 786 376 794 393
rect 811 376 853 393
rect 870 376 900 393
rect 932 411 965 419
rect 932 394 940 411
rect 957 394 965 411
rect 786 375 878 376
rect 634 358 878 375
rect 932 341 965 394
rect 986 393 1019 431
rect 986 376 994 393
rect 1011 376 1019 393
rect 986 368 1019 376
rect 1042 429 1075 437
rect 1042 412 1050 429
rect 1067 412 1075 429
rect 1042 393 1075 412
rect 1042 376 1050 393
rect 1067 376 1075 393
rect 1042 341 1075 376
rect 1126 431 1134 448
rect 1151 439 1187 448
rect 1204 453 1237 457
rect 1151 431 1159 439
rect 1126 393 1159 431
rect 1204 436 1212 453
rect 1229 440 1237 453
rect 1414 452 1439 460
rect 1414 440 1422 452
rect 1229 436 1422 440
rect 1204 435 1422 436
rect 1204 432 1439 435
rect 1456 457 1503 465
rect 1456 440 1478 457
rect 1495 440 1503 457
rect 1456 432 1503 440
rect 1204 423 1284 432
rect 1276 415 1284 423
rect 1301 423 1439 432
rect 1301 415 1309 423
rect 1126 376 1134 393
rect 1151 376 1159 393
rect 1126 368 1159 376
rect 1219 395 1252 406
rect 1219 378 1227 395
rect 1244 378 1252 395
rect 1219 341 1252 378
rect 1276 393 1309 415
rect 1414 415 1439 423
rect 1544 415 1561 490
rect 1633 488 1667 511
rect 1633 476 1658 488
rect 1276 376 1284 393
rect 1301 376 1309 393
rect 1276 368 1309 376
rect 1326 395 1359 406
rect 1326 378 1334 395
rect 1351 378 1359 395
rect 1326 341 1359 378
rect 1414 398 1561 415
rect 1578 459 1613 471
rect 1578 442 1588 459
rect 1605 442 1613 459
rect 1578 418 1613 442
rect 1578 401 1588 418
rect 1605 401 1613 418
rect 1414 393 1439 398
rect 1414 376 1422 393
rect 1578 381 1613 401
rect 1414 368 1439 376
rect 1524 373 1613 381
rect 1524 356 1532 373
rect 1549 356 1588 373
rect 1605 356 1613 373
rect 1633 459 1641 476
rect 1633 434 1658 459
rect 1633 417 1641 434
rect 1633 393 1658 417
rect 1633 376 1641 393
rect 1633 368 1658 376
rect 1678 463 1711 471
rect 1678 446 1686 463
rect 1703 446 1711 463
rect 1678 428 1711 446
rect 1678 411 1686 428
rect 1703 411 1711 428
rect 1678 393 1711 411
rect 1678 376 1686 393
rect 1703 376 1711 393
rect 1524 341 1613 356
rect 1678 341 1711 376
rect 1730 468 1766 511
rect 1849 484 1866 561
rect 1884 623 1909 657
rect 1901 606 1909 623
rect 1933 625 2002 657
rect 1933 608 1941 625
rect 1958 608 1977 625
rect 1994 608 2002 625
rect 2027 623 2052 631
rect 1884 578 1909 606
rect 1901 561 1909 578
rect 1884 553 1909 561
rect 2027 606 2035 623
rect 2027 578 2052 606
rect 2070 612 2103 657
rect 2070 595 2078 612
rect 2095 595 2103 612
rect 2070 585 2103 595
rect 2121 623 2138 631
rect 2027 561 2035 578
rect 2121 578 2138 606
rect 2156 612 2189 657
rect 2156 595 2164 612
rect 2181 595 2189 612
rect 2156 585 2189 595
rect 2207 623 2436 640
rect 2224 606 2232 623
rect 2052 561 2121 565
rect 2207 578 2232 606
rect 2299 612 2332 623
rect 2138 561 2207 565
rect 2224 561 2232 578
rect 2027 548 2232 561
rect 2249 596 2282 605
rect 2249 579 2257 596
rect 2274 579 2282 596
rect 2299 595 2307 612
rect 2324 595 2332 612
rect 2403 612 2436 623
rect 2299 585 2332 595
rect 2349 596 2386 605
rect 2249 565 2282 579
rect 2349 579 2359 596
rect 2376 579 2386 596
rect 2403 595 2411 612
rect 2428 595 2436 612
rect 2403 585 2436 595
rect 2349 565 2386 579
rect 2249 548 2435 565
rect 2412 540 2435 548
rect 2067 523 2243 531
rect 2067 506 2075 523
rect 2092 506 2109 523
rect 2126 506 2141 523
rect 2160 506 2177 523
rect 2194 506 2243 523
rect 2067 498 2243 506
rect 2124 488 2243 498
rect 2260 523 2395 531
rect 2260 506 2268 523
rect 2285 506 2302 523
rect 2319 506 2334 523
rect 2353 506 2370 523
rect 2387 506 2395 523
rect 2260 488 2395 506
rect 2412 500 2470 540
rect 1730 451 1741 468
rect 1758 451 1766 468
rect 1730 432 1766 451
rect 1730 415 1741 432
rect 1758 415 1766 432
rect 1730 397 1766 415
rect 1730 380 1741 397
rect 1758 380 1766 397
rect 1730 372 1766 380
rect 1785 470 1818 484
rect 1785 453 1793 470
rect 1810 453 1818 470
rect 1785 434 1818 453
rect 1785 417 1793 434
rect 1810 417 1818 434
rect 1785 395 1818 417
rect 1785 378 1793 395
rect 1810 378 1818 395
rect 1785 341 1818 378
rect 1835 476 1866 484
rect 1835 459 1838 476
rect 1855 471 1866 476
rect 1835 454 1840 459
rect 1857 454 1866 471
rect 1835 435 1866 454
rect 1835 434 1840 435
rect 1835 417 1838 434
rect 1857 418 1866 435
rect 1855 417 1866 418
rect 1835 393 1866 417
rect 1835 376 1838 393
rect 1855 376 1866 393
rect 1835 368 1866 376
rect 1883 476 1908 484
rect 1900 459 1908 476
rect 1883 434 1908 459
rect 1900 417 1908 434
rect 1883 393 1908 417
rect 1900 376 1908 393
rect 2027 473 2060 481
rect 2027 456 2035 473
rect 2052 456 2060 473
rect 2412 471 2435 500
rect 2027 433 2060 456
rect 2027 416 2035 433
rect 2052 416 2060 433
rect 2027 393 2060 416
rect 1883 341 1908 376
rect 1933 374 1941 391
rect 1958 374 1977 391
rect 1994 374 2002 391
rect 1933 341 2002 374
rect 2027 376 2035 393
rect 2052 376 2060 393
rect 2027 341 2060 376
rect 2077 463 2435 471
rect 2077 446 2081 463
rect 2098 446 2121 463
rect 2138 446 2162 463
rect 2179 454 2257 463
rect 2179 446 2182 454
rect 2077 427 2182 446
rect 2249 446 2257 454
rect 2274 446 2291 463
rect 2308 446 2327 463
rect 2344 446 2361 463
rect 2378 454 2435 463
rect 2378 446 2386 454
rect 2077 410 2081 427
rect 2098 410 2121 427
rect 2138 410 2162 427
rect 2179 410 2182 427
rect 2077 393 2182 410
rect 2077 376 2081 393
rect 2098 376 2121 393
rect 2138 376 2162 393
rect 2179 376 2182 393
rect 2077 368 2182 376
rect 2199 432 2232 437
rect 2199 415 2207 432
rect 2224 415 2232 432
rect 2199 393 2232 415
rect 2199 376 2207 393
rect 2224 376 2232 393
rect 2199 341 2232 376
rect 2249 427 2386 446
rect 2249 410 2257 427
rect 2274 410 2291 427
rect 2308 410 2327 427
rect 2344 410 2361 427
rect 2378 410 2386 427
rect 2249 393 2386 410
rect 2249 376 2257 393
rect 2274 376 2291 393
rect 2308 376 2327 393
rect 2344 376 2361 393
rect 2378 376 2386 393
rect 2249 368 2386 376
rect 2403 432 2436 437
rect 2403 415 2411 432
rect 2428 415 2436 432
rect 2403 393 2436 415
rect 2403 376 2411 393
rect 2428 376 2436 393
rect 2403 341 2436 376
rect -1440 324 -1424 341
rect -1407 324 -1376 341
rect -1359 324 -1328 341
rect -1311 324 -1280 341
rect -1263 324 -1232 341
rect -1215 324 -1184 341
rect -1167 324 -1136 341
rect -1119 324 -1088 341
rect -1071 324 -1040 341
rect -1023 324 -992 341
rect -975 324 -944 341
rect -927 324 -896 341
rect -879 324 -848 341
rect -831 324 -800 341
rect -783 324 -752 341
rect -735 324 -704 341
rect -687 324 -656 341
rect -639 324 -608 341
rect -591 324 -560 341
rect -543 324 -512 341
rect -495 324 -464 341
rect -447 324 -416 341
rect -399 324 -368 341
rect -351 324 -320 341
rect -303 324 -272 341
rect -255 324 -224 341
rect -207 324 -176 341
rect -159 324 -128 341
rect -111 324 -80 341
rect -63 324 -32 341
rect -15 324 15 341
rect 32 324 63 341
rect 80 324 111 341
rect 128 324 159 341
rect 176 324 207 341
rect 224 324 255 341
rect 272 324 303 341
rect 320 324 351 341
rect 368 324 399 341
rect 416 324 447 341
rect 464 324 495 341
rect 512 324 543 341
rect 560 324 591 341
rect 608 324 639 341
rect 656 324 687 341
rect 704 324 735 341
rect 752 324 783 341
rect 800 324 831 341
rect 848 324 879 341
rect 896 324 927 341
rect 944 324 975 341
rect 992 324 1023 341
rect 1040 324 1071 341
rect 1088 324 1119 341
rect 1136 324 1167 341
rect 1184 324 1215 341
rect 1232 324 1263 341
rect 1280 324 1311 341
rect 1328 324 1359 341
rect 1376 324 1407 341
rect 1424 324 1455 341
rect 1472 324 1503 341
rect 1520 324 1551 341
rect 1568 324 1599 341
rect 1616 324 1647 341
rect 1664 324 1695 341
rect 1712 324 1743 341
rect 1760 324 1791 341
rect 1808 324 1839 341
rect 1856 324 1887 341
rect 1904 324 1935 341
rect 1952 324 1983 341
rect 2000 324 2031 341
rect 2048 324 2079 341
rect 2096 324 2127 341
rect 2144 324 2175 341
rect 2192 324 2223 341
rect 2240 324 2271 341
rect 2288 324 2319 341
rect 2336 324 2367 341
rect 2384 324 2415 341
rect 2432 324 2448 341
rect -815 290 -782 324
rect -815 273 -807 290
rect -790 273 -782 290
rect -815 255 -782 273
rect -815 238 -807 255
rect -790 238 -782 255
rect -815 220 -782 238
rect -815 203 -807 220
rect -790 203 -782 220
rect -815 195 -782 203
rect -765 290 -732 298
rect -765 273 -757 290
rect -740 273 -732 290
rect -765 248 -732 273
rect -765 231 -757 248
rect -740 231 -732 248
rect -765 207 -732 231
rect -133 290 -100 324
rect -133 273 -125 290
rect -108 273 -100 290
rect -133 248 -100 273
rect -133 231 -125 248
rect -108 231 -100 248
rect -765 190 -757 207
rect -740 190 -732 207
rect -851 155 -782 178
rect -851 138 -843 155
rect -824 138 -807 155
rect -790 138 -782 155
rect -851 130 -782 138
rect -765 163 -732 190
rect -765 134 -682 163
rect -815 105 -782 113
rect -815 88 -807 105
rect -790 88 -782 105
rect -815 60 -782 88
rect -815 43 -807 60
rect -790 43 -782 60
rect -815 8 -782 43
rect -765 105 -732 134
rect -765 88 -757 105
rect -740 88 -732 105
rect -765 60 -732 88
rect -133 207 -100 231
rect -133 190 -125 207
rect -108 190 -100 207
rect -133 182 -100 190
rect -83 290 -60 298
rect -83 273 -80 290
rect -63 273 -60 290
rect -83 248 -60 273
rect -83 231 -80 248
rect -63 231 -60 248
rect -83 207 -60 231
rect -83 190 -80 207
rect -63 190 -60 207
rect -200 147 -100 155
rect -200 130 -125 147
rect -108 130 -100 147
rect -200 122 -100 130
rect -133 118 -100 122
rect -83 118 -60 190
rect -43 290 -10 324
rect -43 273 -35 290
rect -18 273 -10 290
rect -43 248 -10 273
rect -43 231 -35 248
rect -18 231 -10 248
rect -43 207 -10 231
rect 9 289 87 306
rect 9 272 15 289
rect 32 272 63 289
rect 9 269 63 272
rect 80 269 87 289
rect 9 246 87 269
rect 9 229 15 246
rect 32 229 63 246
rect 80 229 87 246
rect 107 290 132 298
rect 107 273 115 290
rect 107 255 132 273
rect 152 289 185 324
rect 152 272 160 289
rect 177 272 185 289
rect 152 264 185 272
rect 202 290 314 307
rect 107 238 115 255
rect 202 247 219 290
rect 281 273 289 290
rect 306 273 314 290
rect 132 238 219 247
rect 107 230 219 238
rect 236 260 261 273
rect 236 243 244 260
rect 236 230 261 243
rect 281 255 314 273
rect 281 238 289 255
rect 306 238 314 255
rect 281 230 314 238
rect 337 290 370 324
rect 337 273 345 290
rect 362 273 370 290
rect 337 255 370 273
rect 337 238 345 255
rect 362 238 370 255
rect 337 230 370 238
rect 390 290 415 298
rect 407 273 415 290
rect 390 255 415 273
rect 407 238 415 255
rect 9 221 87 229
rect 244 213 261 230
rect -43 190 -35 207
rect -18 190 -10 207
rect -43 182 -10 190
rect 108 205 151 213
rect 108 188 126 205
rect 143 188 151 205
rect 244 196 311 213
rect 108 171 151 188
rect -43 147 -10 155
rect -43 130 -35 147
rect -18 130 -10 147
rect -43 118 -10 130
rect 108 154 126 171
rect 143 154 151 171
rect 108 146 151 154
rect 176 171 227 179
rect 176 154 184 171
rect 201 154 227 171
rect 176 146 227 154
rect 244 171 277 179
rect 244 154 252 171
rect 269 154 277 171
rect 244 146 277 154
rect 108 137 227 146
rect 108 120 126 137
rect 143 120 184 137
rect 201 120 227 137
rect 294 129 311 196
rect 390 181 415 238
rect 438 290 463 298
rect 438 273 446 290
rect 438 255 463 273
rect 438 238 446 255
rect 438 220 463 238
rect 483 290 516 324
rect 483 273 491 290
rect 508 273 516 290
rect 483 251 516 273
rect 483 234 491 251
rect 508 234 516 251
rect 483 229 516 234
rect 536 290 574 298
rect 553 273 574 290
rect 536 249 574 273
rect 553 232 574 249
rect 592 264 617 324
rect 609 247 617 264
rect 592 235 617 247
rect 634 290 878 307
rect 438 203 446 220
rect 463 203 519 212
rect 438 195 519 203
rect 356 173 415 181
rect 356 156 364 173
rect 381 156 415 173
rect 356 148 415 156
rect -77 101 -60 118
rect 108 112 227 120
rect 244 112 373 129
rect 9 102 87 110
rect -131 84 -123 101
rect -106 84 -98 101
rect -77 84 -41 101
rect -24 84 -16 101
rect -765 43 -757 60
rect -740 43 -732 60
rect -765 35 -732 43
rect -131 60 -98 84
rect -131 43 -123 60
rect -106 43 -98 60
rect -131 8 -98 43
rect -49 63 -16 84
rect -49 60 -40 63
rect -49 43 -41 60
rect -23 46 -16 63
rect -24 43 -16 46
rect -49 35 -16 43
rect 9 85 15 102
rect 32 85 63 102
rect 80 85 87 102
rect 9 64 87 85
rect 9 44 15 64
rect 32 61 87 64
rect 32 44 63 61
rect 80 44 87 61
rect 9 26 87 44
rect 110 85 143 112
rect 244 95 265 112
rect 110 68 118 85
rect 135 68 143 85
rect 110 8 143 68
rect 192 87 265 95
rect 192 70 200 87
rect 217 70 240 87
rect 257 70 265 87
rect 192 62 265 70
rect 314 84 339 95
rect 314 67 322 84
rect 314 8 339 67
rect 356 42 373 112
rect 390 90 415 148
rect 444 160 485 178
rect 444 143 460 160
rect 477 143 485 160
rect 444 135 485 143
rect 502 167 519 195
rect 536 209 574 232
rect 634 218 651 290
rect 786 273 794 290
rect 811 273 853 290
rect 870 273 900 290
rect 553 192 574 209
rect 536 184 574 192
rect 502 159 540 167
rect 502 142 515 159
rect 532 142 540 159
rect 502 134 540 142
rect 557 135 574 184
rect 599 208 651 218
rect 599 191 607 208
rect 624 201 651 208
rect 680 260 713 273
rect 680 243 688 260
rect 705 243 713 260
rect 680 221 713 243
rect 730 260 763 273
rect 730 243 738 260
rect 755 255 763 260
rect 755 243 866 255
rect 730 238 866 243
rect 680 204 832 221
rect 624 191 632 201
rect 599 183 632 191
rect 799 187 832 204
rect 745 184 778 185
rect 655 177 778 184
rect 655 176 753 177
rect 655 159 663 176
rect 680 160 753 176
rect 770 160 778 177
rect 680 159 778 160
rect 655 152 778 159
rect 799 170 807 187
rect 824 170 832 187
rect 799 153 832 170
rect 655 138 707 152
rect 655 135 687 138
rect 502 117 519 134
rect 557 121 687 135
rect 704 121 707 138
rect 799 136 807 153
rect 824 136 832 153
rect 799 135 832 136
rect 557 118 707 121
rect 724 118 832 135
rect 438 100 446 117
rect 463 100 519 117
rect 565 101 573 118
rect 407 73 415 90
rect 565 84 590 101
rect 390 59 415 73
rect 432 66 548 83
rect 432 42 449 66
rect 356 25 449 42
rect 489 41 514 49
rect 489 24 497 41
rect 531 42 548 66
rect 565 67 573 84
rect 565 59 590 67
rect 607 84 707 101
rect 607 42 624 84
rect 531 25 624 42
rect 641 59 668 67
rect 641 42 642 59
rect 659 42 668 59
rect 489 8 514 24
rect 641 8 668 42
rect 690 43 707 84
rect 724 92 757 118
rect 849 101 866 238
rect 724 75 732 92
rect 749 75 757 92
rect 724 60 757 75
rect 774 89 866 101
rect 883 229 900 273
rect 932 271 965 324
rect 932 254 940 271
rect 957 254 965 271
rect 932 246 965 254
rect 986 290 1019 298
rect 986 273 994 290
rect 1011 273 1019 290
rect 986 235 1019 273
rect 986 229 994 235
rect 883 218 994 229
rect 1011 218 1019 235
rect 1042 290 1075 324
rect 1042 273 1050 290
rect 1067 273 1075 290
rect 1042 254 1075 273
rect 1042 237 1050 254
rect 1067 237 1075 254
rect 1042 229 1075 237
rect 1126 290 1159 298
rect 1126 273 1134 290
rect 1151 273 1159 290
rect 1126 235 1159 273
rect 1219 287 1252 324
rect 1219 270 1227 287
rect 1244 270 1252 287
rect 1219 260 1252 270
rect 1276 290 1309 298
rect 1276 273 1284 290
rect 1301 273 1309 290
rect 1276 251 1309 273
rect 1326 287 1359 324
rect 1524 309 1613 324
rect 1326 270 1334 287
rect 1351 270 1359 287
rect 1326 260 1359 270
rect 1414 290 1439 298
rect 1414 273 1422 290
rect 1524 292 1532 309
rect 1549 292 1588 309
rect 1605 292 1613 309
rect 1524 284 1613 292
rect 1414 267 1439 273
rect 1276 243 1284 251
rect 883 212 1019 218
rect 1126 218 1134 235
rect 1151 227 1159 235
rect 1204 234 1284 243
rect 1301 243 1309 251
rect 1414 250 1561 267
rect 1414 243 1439 250
rect 1301 234 1439 243
rect 1204 231 1439 234
rect 1204 230 1422 231
rect 1151 218 1187 227
rect 883 111 900 212
rect 986 195 1090 212
rect 1126 210 1187 218
rect 917 187 958 195
rect 917 170 925 187
rect 942 170 958 187
rect 1057 183 1090 195
rect 917 153 958 170
rect 917 136 925 153
rect 942 136 958 153
rect 975 175 1040 178
rect 975 170 1023 175
rect 975 153 983 170
rect 1000 158 1023 170
rect 1057 166 1065 183
rect 1082 166 1090 183
rect 1170 192 1187 210
rect 1204 213 1212 230
rect 1229 226 1422 230
rect 1229 213 1237 226
rect 1204 209 1237 213
rect 1414 214 1422 226
rect 1254 192 1362 209
rect 1414 206 1439 214
rect 1456 225 1503 233
rect 1456 208 1478 225
rect 1495 208 1503 225
rect 1170 175 1271 192
rect 1345 189 1362 192
rect 1456 200 1503 208
rect 1057 158 1090 166
rect 1111 167 1144 175
rect 1000 153 1040 158
rect 975 145 1040 153
rect 1111 150 1119 167
rect 1136 158 1144 167
rect 1136 151 1234 158
rect 1136 150 1209 151
rect 917 128 958 136
rect 1111 138 1209 150
rect 941 111 1068 128
rect 1111 121 1119 138
rect 1136 134 1209 138
rect 1226 134 1234 151
rect 1136 128 1234 134
rect 1136 121 1144 128
rect 1111 118 1144 121
rect 1251 111 1268 175
rect 1291 158 1311 175
rect 1345 172 1432 189
rect 1291 147 1328 158
rect 1399 155 1407 172
rect 1424 155 1432 172
rect 1291 130 1299 147
rect 1316 130 1328 147
rect 1291 118 1328 130
rect 1345 147 1378 155
rect 1399 147 1432 155
rect 1345 130 1353 147
rect 1370 130 1378 147
rect 1456 133 1473 200
rect 1490 176 1523 183
rect 1490 175 1499 176
rect 1490 158 1498 175
rect 1516 159 1523 176
rect 1515 158 1523 159
rect 1490 150 1523 158
rect 1544 176 1561 250
rect 1578 264 1613 284
rect 1578 247 1588 264
rect 1605 247 1613 264
rect 1633 290 1658 298
rect 1633 273 1641 290
rect 1633 252 1658 273
rect 1578 223 1613 247
rect 1578 206 1588 223
rect 1605 206 1613 223
rect 1578 195 1613 206
rect 1632 248 1658 252
rect 1632 245 1641 248
rect 1632 228 1637 245
rect 1654 228 1658 231
rect 1632 209 1658 228
rect 1632 192 1637 209
rect 1654 207 1658 209
rect 1678 290 1711 324
rect 1678 273 1686 290
rect 1703 273 1711 290
rect 1678 255 1711 273
rect 1678 238 1686 255
rect 1703 238 1711 255
rect 1678 220 1711 238
rect 1678 203 1686 220
rect 1703 203 1711 220
rect 1678 195 1711 203
rect 1730 286 1766 294
rect 1730 269 1741 286
rect 1758 269 1766 286
rect 1730 250 1766 269
rect 1730 233 1741 250
rect 1758 233 1766 250
rect 1730 215 1766 233
rect 1730 198 1741 215
rect 1758 198 1766 215
rect 1632 190 1641 192
rect 1632 184 1658 190
rect 1633 178 1658 184
rect 1544 168 1577 176
rect 1544 151 1552 168
rect 1569 151 1577 168
rect 1544 143 1577 151
rect 1633 155 1667 178
rect 1730 155 1766 198
rect 1785 288 1818 324
rect 1785 271 1793 288
rect 1810 271 1818 288
rect 1785 249 1818 271
rect 1785 232 1793 249
rect 1810 232 1818 249
rect 1785 213 1818 232
rect 1785 196 1793 213
rect 1810 196 1818 213
rect 1785 182 1818 196
rect 1835 290 1866 298
rect 1835 273 1838 290
rect 1855 273 1866 290
rect 1835 248 1866 273
rect 1835 231 1838 248
rect 1855 243 1866 248
rect 1835 226 1841 231
rect 1858 226 1866 243
rect 1835 207 1866 226
rect 1835 190 1838 207
rect 1858 190 1866 207
rect 1835 182 1866 190
rect 1883 290 1908 324
rect 1900 273 1908 290
rect 1933 292 2002 324
rect 1933 275 1941 292
rect 1958 275 1977 292
rect 1994 275 2002 292
rect 2028 282 2061 324
rect 1883 248 1908 273
rect 1900 231 1908 248
rect 1883 207 1908 231
rect 1900 190 1908 207
rect 2028 265 2036 282
rect 2053 265 2061 282
rect 2028 227 2061 265
rect 2028 210 2036 227
rect 2053 210 2061 227
rect 2028 202 2061 210
rect 2081 282 2098 290
rect 2081 227 2098 265
rect 2118 284 2151 324
rect 2221 290 2254 324
rect 2118 267 2126 284
rect 2143 267 2151 284
rect 2118 250 2151 267
rect 2118 233 2126 250
rect 2143 233 2151 250
rect 2118 229 2151 233
rect 2168 282 2201 290
rect 2168 265 2176 282
rect 2193 265 2201 282
rect 2168 227 2201 265
rect 2221 273 2229 290
rect 2246 273 2254 290
rect 2221 254 2254 273
rect 2221 237 2229 254
rect 2246 237 2254 254
rect 2221 229 2254 237
rect 2276 290 2301 298
rect 2293 273 2301 290
rect 2276 249 2301 273
rect 2293 232 2301 249
rect 2168 212 2176 227
rect 2098 210 2176 212
rect 2193 212 2201 227
rect 2193 210 2259 212
rect 1883 182 1908 190
rect 2081 195 2259 210
rect 1456 130 1511 133
rect 1345 125 1511 130
rect 883 94 924 111
rect 774 72 782 89
rect 799 84 866 89
rect 799 72 807 84
rect 774 43 807 72
rect 891 77 899 94
rect 916 77 924 94
rect 690 26 807 43
rect 830 59 873 67
rect 891 60 924 77
rect 941 85 984 93
rect 941 68 954 85
rect 971 68 984 85
rect 941 60 984 68
rect 1001 85 1034 94
rect 1001 68 1009 85
rect 1026 68 1034 85
rect 830 42 843 59
rect 860 43 873 59
rect 941 43 958 60
rect 860 42 958 43
rect 830 26 958 42
rect 1001 8 1034 68
rect 1051 43 1068 111
rect 1190 94 1268 111
rect 1345 113 1486 125
rect 1345 94 1362 113
rect 1456 108 1486 113
rect 1503 108 1511 125
rect 1456 100 1511 108
rect 1544 100 1561 143
rect 1633 122 1657 155
rect 1190 85 1207 94
rect 1092 77 1207 85
rect 1285 77 1362 94
rect 1379 86 1404 96
rect 1092 60 1100 77
rect 1117 60 1141 77
rect 1158 60 1182 77
rect 1199 60 1207 77
rect 1230 60 1302 77
rect 1396 83 1404 86
rect 1528 83 1561 100
rect 1578 105 1607 113
rect 1578 88 1589 105
rect 1606 88 1607 105
rect 1396 69 1545 83
rect 1379 66 1545 69
rect 1230 43 1247 60
rect 1319 43 1332 60
rect 1349 43 1361 60
rect 1379 59 1404 66
rect 1578 60 1607 88
rect 1051 26 1247 43
rect 1264 26 1274 43
rect 1291 26 1301 43
rect 1264 8 1301 26
rect 1319 42 1361 43
rect 1422 42 1430 49
rect 1319 32 1430 42
rect 1447 32 1455 49
rect 1319 25 1455 32
rect 1578 43 1589 60
rect 1606 43 1607 60
rect 1578 8 1607 43
rect 1624 105 1657 122
rect 1730 147 1832 155
rect 1730 130 1807 147
rect 1824 130 1832 147
rect 1730 122 1832 130
rect 1624 88 1632 105
rect 1649 88 1657 105
rect 1624 60 1657 88
rect 1624 43 1632 60
rect 1649 43 1657 60
rect 1624 35 1657 43
rect 1674 105 1707 113
rect 1674 88 1675 105
rect 1692 88 1707 105
rect 1674 60 1707 88
rect 1674 43 1675 60
rect 1692 43 1707 60
rect 1730 107 1763 122
rect 1730 90 1738 107
rect 1755 90 1763 107
rect 1849 105 1866 182
rect 2081 128 2098 195
rect 2122 170 2155 178
rect 2122 153 2130 170
rect 2148 153 2155 170
rect 2122 145 2155 153
rect 2172 171 2222 178
rect 2172 167 2225 171
rect 2172 150 2193 167
rect 2210 159 2225 167
rect 2172 142 2197 150
rect 2214 145 2225 159
rect 2242 167 2259 195
rect 2276 209 2301 232
rect 2321 290 2346 324
rect 2338 273 2346 290
rect 2321 243 2346 273
rect 2338 226 2346 243
rect 2321 218 2346 226
rect 2366 290 2393 298
rect 2383 273 2393 290
rect 2366 249 2393 273
rect 2383 232 2393 249
rect 2293 201 2301 209
rect 2366 209 2393 232
rect 2293 192 2366 201
rect 2383 192 2393 209
rect 2276 184 2393 192
rect 2242 159 2347 167
rect 2214 142 2222 145
rect 2172 134 2222 142
rect 2242 142 2254 159
rect 2271 142 2288 159
rect 2305 142 2322 159
rect 2339 142 2347 159
rect 2364 163 2393 184
rect 2411 290 2436 324
rect 2428 273 2436 290
rect 2411 248 2436 273
rect 2428 231 2436 248
rect 2411 207 2436 231
rect 2428 190 2436 207
rect 2411 182 2436 190
rect 2458 163 2487 172
rect 2364 155 2487 163
rect 2242 134 2347 142
rect 2368 143 2487 155
rect 2027 117 2060 125
rect 1730 73 1763 90
rect 1730 56 1738 73
rect 1755 56 1763 73
rect 1730 54 1763 56
rect 1783 97 1816 105
rect 1783 80 1791 97
rect 1808 80 1816 97
rect 1783 60 1816 80
rect 1674 8 1707 43
rect 1783 43 1791 60
rect 1808 43 1816 60
rect 1783 8 1816 43
rect 1833 97 1866 105
rect 1833 80 1841 97
rect 1858 80 1866 97
rect 1833 60 1866 80
rect 1833 43 1841 60
rect 1858 43 1866 60
rect 1833 35 1866 43
rect 1884 105 1909 113
rect 1901 88 1909 105
rect 1884 60 1909 88
rect 1901 43 1909 60
rect 2027 100 2035 117
rect 2052 100 2060 117
rect 2081 119 2148 128
rect 2081 111 2123 119
rect 2027 82 2060 100
rect 2115 102 2123 111
rect 2140 102 2148 119
rect 2368 117 2393 143
rect 2458 132 2487 143
rect 2027 65 2035 82
rect 2052 65 2060 82
rect 1884 8 1909 43
rect 1933 41 1941 58
rect 1958 41 1977 58
rect 1994 41 2002 58
rect 1933 8 2002 41
rect 2027 8 2060 65
rect 2080 84 2097 94
rect 2080 42 2097 67
rect 2115 80 2148 102
rect 2115 63 2123 80
rect 2140 63 2148 80
rect 2115 59 2148 63
rect 2165 114 2198 117
rect 2165 97 2173 114
rect 2190 97 2198 114
rect 2165 80 2198 97
rect 2165 63 2173 80
rect 2190 63 2198 80
rect 2165 42 2198 63
rect 2080 25 2198 42
rect 2216 100 2224 117
rect 2241 100 2249 117
rect 2216 78 2249 100
rect 2216 61 2224 78
rect 2241 61 2249 78
rect 2216 8 2249 61
rect 2275 109 2368 117
rect 2292 100 2368 109
rect 2385 100 2393 117
rect 2292 92 2300 100
rect 2275 72 2300 92
rect 2292 55 2300 72
rect 2275 47 2300 55
rect 2317 75 2350 83
rect 2317 58 2325 75
rect 2342 58 2350 75
rect 2317 8 2350 58
rect 2368 72 2393 100
rect 2385 55 2393 72
rect 2368 47 2393 55
rect 2411 117 2436 125
rect 2428 100 2436 117
rect 2411 72 2436 100
rect 2428 55 2436 72
rect 2411 8 2436 55
rect -864 -8 -848 8
rect -831 -8 -800 8
rect -783 -8 -752 8
rect -735 -8 -704 8
rect -687 -8 -656 8
rect -639 -8 -608 8
rect -591 -8 -560 8
rect -543 -8 -512 8
rect -495 -8 -464 8
rect -447 -8 -416 8
rect -399 -8 -368 8
rect -351 -8 -320 8
rect -303 -8 -272 8
rect -255 -8 -224 8
rect -207 -8 -176 8
rect -159 -8 -128 8
rect -111 -8 -80 8
rect -63 -8 -32 8
rect -15 -8 15 8
rect 32 -8 63 8
rect 80 -8 111 8
rect 128 -8 159 8
rect 176 -8 207 8
rect 224 -8 255 8
rect 272 -8 303 8
rect 320 -8 351 8
rect 368 -8 399 8
rect 416 -8 447 8
rect 464 -8 495 8
rect 512 -8 543 8
rect 560 -8 591 8
rect 608 -8 639 8
rect 656 -8 687 8
rect 704 -8 735 8
rect 752 -8 783 8
rect 800 -8 831 8
rect 848 -8 879 8
rect 896 -8 927 8
rect 944 -8 975 8
rect 992 -8 1023 8
rect 1040 -8 1071 8
rect 1088 -8 1119 8
rect 1136 -8 1167 8
rect 1184 -8 1215 8
rect 1232 -8 1263 8
rect 1280 -8 1311 8
rect 1328 -8 1359 8
rect 1376 -8 1407 8
rect 1424 -8 1455 8
rect 1472 -8 1503 8
rect 1520 -8 1551 8
rect 1568 -8 1599 8
rect 1616 -8 1647 8
rect 1664 -8 1695 8
rect 1712 -8 1743 8
rect 1760 -8 1791 8
rect 1808 -8 1839 8
rect 1856 -8 1887 8
rect 1904 -8 1935 8
rect 1952 -8 1983 8
rect 2000 -8 2031 8
rect 2048 -8 2079 8
rect 2096 -8 2127 8
rect 2144 -8 2175 8
rect 2192 -8 2223 8
rect 2240 -8 2271 8
rect 2288 -8 2319 8
rect 2336 -8 2367 8
rect 2384 -8 2415 8
rect 2432 -8 2448 8
rect -768 -79 -703 -62
rect -624 -79 -576 -62
rect -768 -110 -734 -79
rect -768 -388 -751 -110
rect -593 -110 -576 -79
rect -694 -155 -677 -147
rect -694 -351 -677 -343
rect -650 -155 -633 -147
rect -650 -351 -633 -343
rect -680 -385 -672 -368
rect -655 -385 -647 -368
rect -768 -419 -734 -388
rect -593 -419 -576 -388
rect -768 -436 -703 -419
rect -624 -436 -576 -419
rect -768 -467 -734 -436
rect -768 -745 -751 -467
rect -593 -467 -576 -436
rect -694 -512 -677 -504
rect -694 -708 -677 -700
rect -650 -512 -633 -504
rect -650 -708 -633 -700
rect -680 -742 -672 -725
rect -655 -742 -647 -725
rect -768 -776 -734 -745
rect -593 -776 -576 -745
rect -768 -793 -703 -776
rect -624 -793 -576 -776
<< viali >>
rect -869 1542 -852 1730
rect -825 1542 -808 1730
rect -768 1539 -751 1733
rect -847 1500 -830 1517
rect -869 1185 -852 1373
rect -825 1185 -808 1373
rect -768 1182 -751 1376
rect -847 1143 -830 1160
rect -535 1539 -518 1733
rect -478 1542 -461 1730
rect -434 1542 -417 1730
rect -456 1500 -439 1517
rect -535 1182 -518 1376
rect -478 1185 -461 1373
rect -434 1185 -417 1373
rect -456 1143 -439 1160
rect -1424 990 -1407 1007
rect -1376 990 -1359 1007
rect -1328 990 -1311 1007
rect -1280 990 -1263 1007
rect -1232 990 -1215 1007
rect -1184 990 -1167 1007
rect -1136 990 -1119 1007
rect -1088 990 -1071 1007
rect -1040 990 -1023 1007
rect -992 990 -975 1007
rect -944 990 -927 1007
rect -896 990 -879 1007
rect -848 990 -831 1007
rect -800 990 -783 1007
rect -752 990 -735 1007
rect -704 990 -687 1007
rect -656 990 -639 1007
rect -608 990 -591 1007
rect -560 990 -543 1007
rect -512 990 -495 1007
rect -464 990 -447 1007
rect -416 990 -399 1007
rect -368 990 -351 1007
rect -320 990 -303 1007
rect -272 990 -255 1007
rect -224 990 -207 1007
rect -176 990 -159 1007
rect -128 990 -111 1007
rect -80 990 -63 1007
rect -32 990 -15 1007
rect 15 990 32 1007
rect 63 990 80 1007
rect 111 990 128 1007
rect 159 990 176 1007
rect 207 990 224 1007
rect 255 990 272 1007
rect 303 990 320 1007
rect 351 990 368 1007
rect 399 990 416 1007
rect 447 990 464 1007
rect 495 990 512 1007
rect 543 990 560 1007
rect 591 990 608 1007
rect 639 990 656 1007
rect 687 990 704 1007
rect 735 990 752 1007
rect 783 990 800 1007
rect 831 990 848 1007
rect 879 990 896 1007
rect 927 990 944 1007
rect 975 990 992 1007
rect 1023 990 1040 1007
rect 1071 990 1088 1007
rect 1119 990 1136 1007
rect 1167 990 1184 1007
rect 1215 990 1232 1007
rect 1263 990 1280 1007
rect 1311 990 1328 1007
rect 1359 990 1376 1007
rect 1407 990 1424 1007
rect 1455 990 1472 1007
rect 1503 990 1520 1007
rect 1551 990 1568 1007
rect 1599 990 1616 1007
rect 1647 990 1664 1007
rect 1695 990 1712 1007
rect 1743 990 1760 1007
rect 1791 990 1808 1007
rect 1839 990 1856 1007
rect 1887 990 1904 1007
rect 1935 990 1952 1007
rect 1983 990 2000 1007
rect 2031 990 2048 1007
rect 2079 990 2096 1007
rect 2127 990 2144 1007
rect 2175 990 2192 1007
rect 2223 990 2240 1007
rect 2271 990 2288 1007
rect 2319 990 2336 1007
rect 2367 990 2384 1007
rect 2415 990 2432 1007
rect -1419 804 -1417 821
rect -1417 804 -1402 821
rect -1383 804 -1366 821
rect -1249 741 -1050 866
rect -983 741 -785 866
rect -611 796 -594 813
rect -616 726 -599 729
rect -616 712 -600 726
rect -600 712 -599 726
rect 63 938 80 952
rect 63 935 80 938
rect 15 727 32 730
rect 15 713 32 727
rect -1424 657 -1407 674
rect -1376 657 -1359 674
rect -1328 657 -1311 674
rect -1280 657 -1263 674
rect -1232 657 -1215 674
rect -1184 657 -1167 674
rect -1136 657 -1119 674
rect -1088 657 -1071 674
rect -1040 657 -1023 674
rect -992 657 -975 674
rect -944 657 -927 674
rect -896 657 -879 674
rect -848 657 -831 674
rect -800 657 -783 674
rect -752 657 -735 674
rect -704 657 -687 674
rect -656 657 -639 674
rect -608 657 -591 674
rect -560 657 -543 674
rect -512 657 -495 674
rect -464 657 -447 674
rect -416 657 -399 674
rect -368 657 -351 674
rect -320 657 -303 674
rect -272 657 -255 674
rect -224 657 -207 674
rect -176 657 -159 674
rect -128 657 -111 674
rect -80 657 -63 674
rect -32 657 -15 674
rect 15 657 32 674
rect 63 657 80 674
rect 111 657 128 674
rect 159 657 176 674
rect 207 657 224 674
rect 255 657 272 674
rect 303 657 320 674
rect 351 657 368 674
rect 399 657 416 674
rect 447 657 464 674
rect 495 657 512 674
rect 543 657 560 674
rect 591 657 608 674
rect 639 657 656 674
rect 687 657 704 674
rect 735 657 752 674
rect 783 657 800 674
rect 831 657 848 674
rect 879 657 896 674
rect 927 657 944 674
rect 975 657 992 674
rect 1023 657 1040 674
rect 1071 657 1088 674
rect 1119 657 1136 674
rect 1167 657 1184 674
rect 1215 657 1232 674
rect 1263 657 1280 674
rect 1311 657 1328 674
rect 1359 657 1376 674
rect 1407 657 1424 674
rect 1455 657 1472 674
rect 1503 657 1520 674
rect 1551 657 1568 674
rect 1599 657 1616 674
rect 1647 657 1664 674
rect 1695 657 1712 674
rect 1743 657 1760 674
rect 1791 657 1808 674
rect 1839 657 1856 674
rect 1887 657 1904 674
rect 1935 657 1952 674
rect 1983 657 2000 674
rect 2031 657 2048 674
rect 2079 657 2096 674
rect 2127 657 2144 674
rect 2175 657 2192 674
rect 2223 657 2240 674
rect 2271 657 2288 674
rect 2319 657 2336 674
rect 2367 657 2384 674
rect 2415 657 2432 674
rect -1419 511 -1417 528
rect -1417 511 -1402 528
rect -1383 511 -1366 528
rect -1249 465 -1050 590
rect -983 465 -785 590
rect -616 606 -600 620
rect -600 606 -599 620
rect -616 603 -599 606
rect -611 519 -594 536
rect -518 523 -501 524
rect -518 507 -517 523
rect -517 507 -501 523
rect -379 519 -362 536
rect 15 605 32 619
rect 15 602 32 605
rect -322 536 -305 537
rect -322 520 -305 536
rect -126 528 -109 530
rect -126 513 -125 528
rect -125 513 -109 528
rect -180 434 -163 443
rect -180 426 -171 434
rect -171 426 -163 434
rect -79 393 -62 407
rect -79 390 -63 393
rect -63 390 -62 393
rect 254 495 269 512
rect 269 495 271 512
rect 458 506 460 523
rect 460 506 475 523
rect 63 394 80 397
rect 63 380 80 394
rect 687 528 704 545
rect 1119 528 1136 545
rect 1023 491 1040 508
rect 1311 491 1328 508
rect 1498 490 1515 507
rect 2141 506 2143 523
rect 2143 506 2158 523
rect 2177 506 2194 523
rect 2334 506 2336 523
rect 2336 506 2351 523
rect 2370 506 2387 523
rect 1840 459 1855 471
rect 1855 459 1857 471
rect 1840 454 1857 459
rect 1840 434 1857 435
rect 1840 418 1855 434
rect 1855 418 1857 434
rect -1424 324 -1407 341
rect -1376 324 -1359 341
rect -1328 324 -1311 341
rect -1280 324 -1263 341
rect -1232 324 -1215 341
rect -1184 324 -1167 341
rect -1136 324 -1119 341
rect -1088 324 -1071 341
rect -1040 324 -1023 341
rect -992 324 -975 341
rect -944 324 -927 341
rect -896 324 -879 341
rect -848 324 -831 341
rect -800 324 -783 341
rect -752 324 -735 341
rect -704 324 -687 341
rect -656 324 -639 341
rect -608 324 -591 341
rect -560 324 -543 341
rect -512 324 -495 341
rect -464 324 -447 341
rect -416 324 -399 341
rect -368 324 -351 341
rect -320 324 -303 341
rect -272 324 -255 341
rect -224 324 -207 341
rect -176 324 -159 341
rect -128 324 -111 341
rect -80 324 -63 341
rect -32 324 -15 341
rect 15 324 32 341
rect 63 324 80 341
rect 111 324 128 341
rect 159 324 176 341
rect 207 324 224 341
rect 255 324 272 341
rect 303 324 320 341
rect 351 324 368 341
rect 399 324 416 341
rect 447 324 464 341
rect 495 324 512 341
rect 543 324 560 341
rect 591 324 608 341
rect 639 324 656 341
rect 687 324 704 341
rect 735 324 752 341
rect 783 324 800 341
rect 831 324 848 341
rect 879 324 896 341
rect 927 324 944 341
rect 975 324 992 341
rect 1023 324 1040 341
rect 1071 324 1088 341
rect 1119 324 1136 341
rect 1167 324 1184 341
rect 1215 324 1232 341
rect 1263 324 1280 341
rect 1311 324 1328 341
rect 1359 324 1376 341
rect 1407 324 1424 341
rect 1455 324 1472 341
rect 1503 324 1520 341
rect 1551 324 1568 341
rect 1599 324 1616 341
rect 1647 324 1664 341
rect 1695 324 1712 341
rect 1743 324 1760 341
rect 1791 324 1808 341
rect 1839 324 1856 341
rect 1887 324 1904 341
rect 1935 324 1952 341
rect 1983 324 2000 341
rect 2031 324 2048 341
rect 2079 324 2096 341
rect 2127 324 2144 341
rect 2175 324 2192 341
rect 2223 324 2240 341
rect 2271 324 2288 341
rect 2319 324 2336 341
rect 2367 324 2384 341
rect 2415 324 2432 341
rect -843 138 -841 155
rect -841 138 -826 155
rect -807 138 -790 155
rect -673 75 -474 200
rect -407 75 -209 200
rect 63 272 80 286
rect 63 269 80 272
rect -35 130 -18 147
rect 252 154 269 171
rect -40 60 -23 63
rect -40 46 -24 60
rect -24 46 -23 60
rect 15 61 32 64
rect 15 47 32 61
rect 460 143 477 160
rect 687 121 704 138
rect 1023 158 1040 175
rect 1119 121 1136 138
rect 1311 158 1328 175
rect 1499 175 1516 176
rect 1499 159 1515 175
rect 1515 159 1516 175
rect 1637 231 1641 245
rect 1641 231 1654 245
rect 1637 228 1654 231
rect 1637 207 1654 209
rect 1637 192 1641 207
rect 1641 192 1654 207
rect 1841 231 1855 243
rect 1855 231 1858 243
rect 1841 226 1858 231
rect 1841 190 1855 207
rect 1855 190 1858 207
rect 2131 153 2147 170
rect 2147 153 2148 170
rect 2193 159 2210 167
rect 2193 150 2197 159
rect 2197 150 2210 159
rect -848 -8 -831 8
rect -800 -8 -783 8
rect -752 -8 -735 8
rect -704 -8 -687 8
rect -656 -8 -639 8
rect -608 -8 -591 8
rect -560 -8 -543 8
rect -512 -8 -495 8
rect -464 -8 -447 8
rect -416 -8 -399 8
rect -368 -8 -351 8
rect -320 -8 -303 8
rect -272 -8 -255 8
rect -224 -8 -207 8
rect -176 -8 -159 8
rect -128 -8 -111 8
rect -80 -8 -63 8
rect -32 -8 -15 8
rect 15 -8 32 8
rect 63 -8 80 8
rect 111 -8 128 8
rect 159 -8 176 8
rect 207 -8 224 8
rect 255 -8 272 8
rect 303 -8 320 8
rect 351 -8 368 8
rect 399 -8 416 8
rect 447 -8 464 8
rect 495 -8 512 8
rect 543 -8 560 8
rect 591 -8 608 8
rect 639 -8 656 8
rect 687 -8 704 8
rect 735 -8 752 8
rect 783 -8 800 8
rect 831 -8 848 8
rect 879 -8 896 8
rect 927 -8 944 8
rect 975 -8 992 8
rect 1023 -8 1040 8
rect 1071 -8 1088 8
rect 1119 -8 1136 8
rect 1167 -8 1184 8
rect 1215 -8 1232 8
rect 1263 -8 1280 8
rect 1311 -8 1328 8
rect 1359 -8 1376 8
rect 1407 -8 1424 8
rect 1455 -8 1472 8
rect 1503 -8 1520 8
rect 1551 -8 1568 8
rect 1599 -8 1616 8
rect 1647 -8 1664 8
rect 1695 -8 1712 8
rect 1743 -8 1760 8
rect 1791 -8 1808 8
rect 1839 -8 1856 8
rect 1887 -8 1904 8
rect 1935 -8 1952 8
rect 1983 -8 2000 8
rect 2031 -8 2048 8
rect 2079 -8 2096 8
rect 2127 -8 2144 8
rect 2175 -8 2192 8
rect 2223 -8 2240 8
rect 2271 -8 2288 8
rect 2319 -8 2336 8
rect 2367 -8 2384 8
rect 2415 -8 2432 8
rect -751 -346 -734 -152
rect -694 -343 -677 -155
rect -650 -343 -633 -155
rect -672 -385 -655 -368
rect -751 -703 -734 -509
rect -694 -700 -677 -512
rect -650 -700 -633 -512
rect -672 -742 -655 -725
<< metal1 >>
rect -929 1736 -869 1737
rect -416 1736 -356 1737
rect -929 1732 -849 1736
rect -929 1547 -924 1732
rect -874 1730 -849 1732
rect -874 1547 -869 1730
rect -929 1542 -869 1547
rect -852 1542 -849 1730
rect -872 1536 -849 1542
rect -828 1733 -734 1736
rect -828 1730 -768 1733
rect -828 1542 -825 1730
rect -808 1726 -768 1730
rect -783 1546 -768 1726
rect -808 1542 -768 1546
rect -828 1539 -768 1542
rect -751 1539 -734 1733
rect -828 1536 -734 1539
rect -552 1733 -458 1736
rect -552 1539 -535 1733
rect -518 1730 -458 1733
rect -518 1726 -478 1730
rect -518 1546 -503 1726
rect -518 1542 -478 1546
rect -461 1542 -458 1730
rect -518 1539 -458 1542
rect -552 1536 -458 1539
rect -437 1732 -356 1736
rect -437 1730 -411 1732
rect -437 1542 -434 1730
rect -417 1547 -411 1730
rect -361 1547 -356 1732
rect -417 1542 -356 1547
rect -437 1536 -414 1542
rect -855 1517 -782 1520
rect -855 1500 -847 1517
rect -830 1513 -782 1517
rect -830 1500 -815 1513
rect -855 1492 -815 1500
rect -822 1487 -815 1492
rect -789 1487 -782 1513
rect -822 1480 -782 1487
rect -504 1517 -431 1520
rect -504 1513 -456 1517
rect -504 1487 -497 1513
rect -471 1500 -456 1513
rect -439 1500 -431 1517
rect -471 1492 -431 1500
rect -471 1487 -464 1492
rect -504 1480 -464 1487
rect -872 1375 -849 1379
rect -929 1373 -849 1375
rect -929 1370 -869 1373
rect -929 1185 -924 1370
rect -874 1185 -869 1370
rect -852 1185 -849 1373
rect -929 1180 -849 1185
rect -872 1179 -849 1180
rect -828 1376 -734 1379
rect -828 1373 -768 1376
rect -828 1185 -825 1373
rect -808 1367 -768 1373
rect -808 1185 -768 1192
rect -828 1182 -768 1185
rect -751 1182 -734 1376
rect -828 1179 -734 1182
rect -552 1376 -458 1379
rect -552 1182 -535 1376
rect -518 1373 -458 1376
rect -518 1367 -478 1373
rect -518 1185 -478 1192
rect -461 1185 -458 1373
rect -518 1182 -458 1185
rect -552 1179 -458 1182
rect -437 1375 -414 1379
rect -437 1373 -356 1375
rect -437 1185 -434 1373
rect -417 1370 -356 1373
rect -417 1185 -411 1370
rect -361 1185 -356 1370
rect -437 1180 -356 1185
rect -437 1179 -414 1180
rect -855 1160 -782 1163
rect -855 1143 -847 1160
rect -830 1156 -782 1160
rect -830 1143 -815 1156
rect -855 1135 -815 1143
rect -822 1130 -815 1135
rect -789 1130 -782 1156
rect -822 1123 -782 1130
rect -504 1160 -431 1163
rect -504 1156 -456 1160
rect -504 1130 -497 1156
rect -471 1143 -456 1156
rect -439 1143 -431 1160
rect -471 1135 -431 1143
rect -471 1130 -464 1135
rect -504 1123 -464 1130
rect -1440 1020 2448 1023
rect -1440 1007 120 1020
rect 330 1007 720 1020
rect 930 1007 1320 1020
rect 1530 1007 1920 1020
rect 2130 1007 2448 1020
rect -1440 990 -1424 1007
rect -1407 990 -1376 1007
rect -1359 990 -1328 1007
rect -1311 990 -1280 1007
rect -1263 990 -1232 1007
rect -1215 990 -1184 1007
rect -1167 990 -1136 1007
rect -1119 990 -1088 1007
rect -1071 990 -1040 1007
rect -1023 990 -992 1007
rect -975 990 -944 1007
rect -927 990 -896 1007
rect -879 990 -848 1007
rect -831 990 -800 1007
rect -783 990 -752 1007
rect -735 990 -704 1007
rect -687 990 -656 1007
rect -639 990 -608 1007
rect -591 990 -560 1007
rect -543 990 -512 1007
rect -495 990 -464 1007
rect -447 990 -416 1007
rect -399 990 -368 1007
rect -351 990 -320 1007
rect -303 990 -272 1007
rect -255 990 -224 1007
rect -207 990 -176 1007
rect -159 990 -128 1007
rect -111 990 -80 1007
rect -63 990 -32 1007
rect -15 990 15 1007
rect 32 990 63 1007
rect 80 990 111 1007
rect 330 990 351 1007
rect 368 990 399 1007
rect 416 990 447 1007
rect 464 990 495 1007
rect 512 990 543 1007
rect 560 990 591 1007
rect 608 990 639 1007
rect 656 990 687 1007
rect 704 990 720 1007
rect 944 990 975 1007
rect 992 990 1023 1007
rect 1040 990 1071 1007
rect 1088 990 1119 1007
rect 1136 990 1167 1007
rect 1184 990 1215 1007
rect 1232 990 1263 1007
rect 1280 990 1311 1007
rect 1530 990 1551 1007
rect 1568 990 1599 1007
rect 1616 990 1647 1007
rect 1664 990 1695 1007
rect 1712 990 1743 1007
rect 1760 990 1791 1007
rect 1808 990 1839 1007
rect 1856 990 1887 1007
rect 1904 990 1920 1007
rect 2144 990 2175 1007
rect 2192 990 2223 1007
rect 2240 990 2271 1007
rect 2288 990 2319 1007
rect 2336 990 2367 1007
rect 2384 990 2415 1007
rect 2432 990 2448 1007
rect -1440 980 120 990
rect 330 980 720 990
rect 930 980 1320 990
rect 1530 980 1920 990
rect 2130 980 2448 990
rect -1440 974 2448 980
rect 56 952 88 956
rect 56 935 63 952
rect 80 935 88 952
rect 56 930 88 935
rect -1338 895 -586 928
rect -1338 836 -1305 895
rect -1390 825 -1305 836
rect -1427 799 -1424 825
rect -1398 799 -1388 825
rect -1362 803 -1305 825
rect -1255 866 -1044 869
rect -1362 799 -1359 803
rect -1255 741 -1249 866
rect -1050 741 -1044 866
rect -1255 738 -1044 741
rect -989 866 -779 869
rect -989 741 -983 866
rect -785 741 -779 866
rect -619 813 -586 895
rect -619 796 -611 813
rect -594 796 -586 813
rect -619 788 -586 796
rect -989 738 -779 741
rect -621 733 -595 739
rect 8 730 40 734
rect 8 713 15 730
rect 32 713 40 730
rect 8 708 40 713
rect -621 704 -595 707
rect -1440 674 -230 690
rect -20 680 2448 690
rect -20 674 420 680
rect 630 674 1020 680
rect 1230 674 1620 680
rect 1830 674 2220 680
rect 2430 674 2448 680
rect -1440 657 -1424 674
rect -1407 657 -1376 674
rect -1359 657 -1328 674
rect -1311 657 -1280 674
rect -1263 657 -1232 674
rect -1215 657 -1184 674
rect -1167 657 -1136 674
rect -1119 657 -1088 674
rect -1071 657 -1040 674
rect -1023 657 -992 674
rect -975 657 -944 674
rect -927 657 -896 674
rect -879 657 -848 674
rect -831 657 -800 674
rect -783 657 -752 674
rect -735 657 -704 674
rect -687 657 -656 674
rect -639 657 -608 674
rect -591 657 -560 674
rect -543 657 -512 674
rect -495 657 -464 674
rect -447 657 -416 674
rect -399 657 -368 674
rect -351 657 -320 674
rect -303 657 -272 674
rect -255 657 -230 674
rect -15 657 15 674
rect 32 657 63 674
rect 80 657 111 674
rect 128 657 159 674
rect 176 657 207 674
rect 224 657 255 674
rect 272 657 303 674
rect 320 657 351 674
rect 368 657 399 674
rect 416 657 420 674
rect 630 657 639 674
rect 656 657 687 674
rect 704 657 735 674
rect 752 657 783 674
rect 800 657 831 674
rect 848 657 879 674
rect 896 657 927 674
rect 944 657 975 674
rect 992 657 1020 674
rect 1232 657 1263 674
rect 1280 657 1311 674
rect 1328 657 1359 674
rect 1376 657 1407 674
rect 1424 657 1455 674
rect 1472 657 1503 674
rect 1520 657 1551 674
rect 1568 657 1599 674
rect 1616 657 1620 674
rect 1830 657 1839 674
rect 1856 657 1887 674
rect 1904 657 1935 674
rect 1952 657 1983 674
rect 2000 657 2031 674
rect 2048 657 2079 674
rect 2096 657 2127 674
rect 2144 657 2175 674
rect 2192 657 2220 674
rect 2432 657 2448 674
rect -1440 650 -230 657
rect -20 650 420 657
rect 630 650 1020 657
rect 1230 650 1620 657
rect 1830 650 2220 657
rect 2430 650 2448 657
rect -1440 641 2448 650
rect -621 624 -595 627
rect -621 593 -595 598
rect 8 619 40 623
rect 8 602 15 619
rect 32 602 40 619
rect 8 597 40 602
rect -1255 590 -1044 593
rect -1427 506 -1424 532
rect -1398 506 -1388 532
rect -1362 528 -1359 532
rect -1362 506 -1305 528
rect -1390 495 -1305 506
rect -1338 437 -1305 495
rect -1255 465 -1249 590
rect -1050 465 -1044 590
rect -1255 462 -1044 465
rect -989 590 -779 593
rect -989 465 -983 590
rect -785 465 -779 590
rect 681 545 710 548
rect -989 462 -779 465
rect -619 536 -586 544
rect -619 519 -611 536
rect -594 519 -586 536
rect -619 437 -586 519
rect -525 503 -522 529
rect -496 503 -493 529
rect -387 514 -384 540
rect -358 514 -355 540
rect -330 515 -327 541
rect -301 515 -298 541
rect -133 509 -130 535
rect -104 509 -101 535
rect 681 528 687 545
rect 704 543 710 545
rect 1113 545 1142 548
rect 1113 543 1119 545
rect 704 529 1119 543
rect 704 528 710 529
rect 248 512 277 517
rect 248 495 254 512
rect 271 495 277 512
rect 451 501 454 527
rect 480 501 483 527
rect 681 525 710 528
rect 1113 528 1119 529
rect 1136 528 1142 545
rect 1113 525 1142 528
rect 1017 508 1046 511
rect 248 491 277 495
rect 1017 491 1023 508
rect 1040 506 1046 508
rect 1305 508 1334 511
rect 1305 506 1311 508
rect 1040 492 1311 506
rect 1040 491 1046 492
rect -1338 404 -586 437
rect -187 422 -184 448
rect -158 422 -155 448
rect -83 412 -57 415
rect -83 383 -57 386
rect 56 397 88 401
rect 56 380 63 397
rect 80 380 88 397
rect 56 375 88 380
rect 250 357 273 491
rect 1017 488 1046 491
rect 1305 491 1311 492
rect 1328 491 1334 508
rect 1305 488 1334 491
rect 1316 357 1330 488
rect 1490 485 1493 511
rect 1519 485 1522 511
rect 2133 501 2136 527
rect 2162 501 2172 527
rect 2198 501 2201 527
rect 2327 501 2330 527
rect 2356 501 2366 527
rect 2392 501 2395 527
rect 1835 476 1861 479
rect 1835 440 1861 450
rect 1835 411 1861 414
rect -1440 350 2448 357
rect -1440 341 120 350
rect 330 341 720 350
rect 930 341 1320 350
rect 1530 341 1920 350
rect 2130 341 2448 350
rect -1440 324 -1424 341
rect -1407 324 -1376 341
rect -1359 324 -1328 341
rect -1311 324 -1280 341
rect -1263 324 -1232 341
rect -1215 324 -1184 341
rect -1167 324 -1136 341
rect -1119 324 -1088 341
rect -1071 324 -1040 341
rect -1023 324 -992 341
rect -975 324 -944 341
rect -927 324 -896 341
rect -879 324 -848 341
rect -831 324 -800 341
rect -783 324 -752 341
rect -735 324 -704 341
rect -687 324 -656 341
rect -639 324 -608 341
rect -591 324 -560 341
rect -543 324 -512 341
rect -495 324 -464 341
rect -447 324 -416 341
rect -399 324 -368 341
rect -351 324 -320 341
rect -303 324 -272 341
rect -255 324 -224 341
rect -207 324 -176 341
rect -159 324 -128 341
rect -111 324 -80 341
rect -63 324 -32 341
rect -15 324 15 341
rect 32 324 63 341
rect 80 324 111 341
rect 330 324 351 341
rect 368 324 399 341
rect 416 324 447 341
rect 464 324 495 341
rect 512 324 543 341
rect 560 324 591 341
rect 608 324 639 341
rect 656 324 687 341
rect 704 324 720 341
rect 944 324 975 341
rect 992 324 1023 341
rect 1040 324 1071 341
rect 1088 324 1119 341
rect 1136 324 1167 341
rect 1184 324 1215 341
rect 1232 324 1263 341
rect 1280 324 1311 341
rect 1530 324 1551 341
rect 1568 324 1599 341
rect 1616 324 1647 341
rect 1664 324 1695 341
rect 1712 324 1743 341
rect 1760 324 1791 341
rect 1808 324 1839 341
rect 1856 324 1887 341
rect 1904 324 1920 341
rect 2144 324 2175 341
rect 2192 324 2223 341
rect 2240 324 2271 341
rect 2288 324 2319 341
rect 2336 324 2367 341
rect 2384 324 2415 341
rect 2432 324 2448 341
rect -1440 320 120 324
rect 330 320 720 324
rect 930 320 1320 324
rect 1530 320 1920 324
rect 2130 320 2448 324
rect -1440 308 2448 320
rect 56 286 88 290
rect 56 269 63 286
rect 80 269 88 286
rect 56 264 88 269
rect -762 229 -10 262
rect -762 170 -729 229
rect -814 159 -729 170
rect -851 133 -848 159
rect -822 133 -812 159
rect -786 137 -729 159
rect -679 200 -468 203
rect -786 133 -783 137
rect -679 75 -673 200
rect -474 75 -468 200
rect -679 72 -468 75
rect -413 200 -203 203
rect -413 75 -407 200
rect -209 75 -203 200
rect -43 147 -10 229
rect 1316 178 1330 308
rect 1632 249 1658 252
rect 1632 213 1658 223
rect 1632 184 1658 187
rect 1837 247 1863 250
rect 1837 211 1863 221
rect 1837 182 1863 185
rect 1017 175 1046 178
rect 245 149 248 175
rect 274 149 277 175
rect -43 130 -35 147
rect -18 130 -10 147
rect 453 138 456 164
rect 482 138 485 164
rect 1017 158 1023 175
rect 1040 173 1046 175
rect 1305 175 1334 178
rect 1305 173 1311 175
rect 1040 159 1311 173
rect 1040 158 1046 159
rect 1017 155 1046 158
rect 1305 158 1311 159
rect 1328 158 1334 175
rect 1305 155 1334 158
rect 1491 155 1494 181
rect 1520 155 1523 181
rect 2122 175 2155 178
rect 2122 149 2126 175
rect 2152 149 2155 175
rect 2122 145 2155 149
rect 2186 145 2189 171
rect 2215 145 2225 171
rect 681 138 710 141
rect -43 122 -10 130
rect 681 121 687 138
rect 704 136 710 138
rect 1113 138 1142 141
rect 1113 136 1119 138
rect 704 122 1119 136
rect 704 121 710 122
rect 681 118 710 121
rect 1113 121 1119 122
rect 1136 121 1142 138
rect 1113 118 1142 121
rect -413 72 -203 75
rect -45 67 -19 73
rect 8 64 40 68
rect 8 47 15 64
rect 32 47 40 64
rect 8 42 40 47
rect -45 38 -19 41
rect -864 10 2448 24
rect -864 8 420 10
rect 630 8 1020 10
rect 1230 8 1620 10
rect 1830 8 2220 10
rect 2430 8 2448 10
rect -864 -8 -848 8
rect -831 -8 -800 8
rect -783 -8 -752 8
rect -735 -8 -704 8
rect -687 -8 -656 8
rect -639 -8 -608 8
rect -591 -8 -560 8
rect -543 -8 -512 8
rect -495 -8 -464 8
rect -447 -8 -416 8
rect -399 -8 -368 8
rect -351 -8 -320 8
rect -303 -8 -272 8
rect -255 -8 -224 8
rect -207 -8 -176 8
rect -159 -8 -128 8
rect -111 -8 -80 8
rect -63 -8 -32 8
rect -15 -8 15 8
rect 32 -8 63 8
rect 80 -8 111 8
rect 128 -8 159 8
rect 176 -8 207 8
rect 224 -8 255 8
rect 272 -8 303 8
rect 320 -8 351 8
rect 368 -8 399 8
rect 416 -8 420 8
rect 630 -8 639 8
rect 656 -8 687 8
rect 704 -8 735 8
rect 752 -8 783 8
rect 800 -8 831 8
rect 848 -8 879 8
rect 896 -8 927 8
rect 944 -8 975 8
rect 992 -8 1020 8
rect 1232 -8 1263 8
rect 1280 -8 1311 8
rect 1328 -8 1359 8
rect 1376 -8 1407 8
rect 1424 -8 1455 8
rect 1472 -8 1503 8
rect 1520 -8 1551 8
rect 1568 -8 1599 8
rect 1616 -8 1620 8
rect 1830 -8 1839 8
rect 1856 -8 1887 8
rect 1904 -8 1935 8
rect 1952 -8 1983 8
rect 2000 -8 2031 8
rect 2048 -8 2079 8
rect 2096 -8 2127 8
rect 2144 -8 2175 8
rect 2192 -8 2220 8
rect 2432 -8 2448 8
rect -864 -20 420 -8
rect 630 -20 1020 -8
rect 1230 -20 1620 -8
rect 1830 -20 2220 -8
rect 2430 -20 2448 -8
rect -864 -24 2448 -20
rect -633 -149 -573 -147
rect -768 -152 -674 -149
rect -768 -346 -751 -152
rect -734 -155 -674 -152
rect -734 -159 -694 -155
rect -734 -339 -719 -159
rect -734 -343 -694 -339
rect -677 -343 -674 -155
rect -734 -346 -674 -343
rect -768 -349 -674 -346
rect -653 -152 -573 -149
rect -653 -155 -628 -152
rect -653 -343 -650 -155
rect -633 -337 -628 -155
rect -578 -337 -573 -152
rect -633 -342 -573 -337
rect -633 -343 -630 -342
rect -653 -349 -630 -343
rect -720 -368 -647 -365
rect -720 -372 -672 -368
rect -720 -398 -713 -372
rect -687 -385 -672 -372
rect -655 -385 -647 -368
rect -687 -393 -647 -385
rect -687 -398 -680 -393
rect -720 -405 -680 -398
rect -768 -509 -674 -506
rect -768 -703 -751 -509
rect -734 -512 -674 -509
rect -734 -518 -694 -512
rect -734 -700 -694 -693
rect -677 -700 -674 -512
rect -734 -703 -674 -700
rect -768 -706 -674 -703
rect -653 -509 -630 -506
rect -653 -512 -573 -509
rect -653 -700 -650 -512
rect -633 -514 -573 -512
rect -633 -699 -628 -514
rect -578 -699 -573 -514
rect -633 -700 -573 -699
rect -653 -704 -573 -700
rect -653 -706 -630 -704
rect -720 -725 -647 -722
rect -720 -729 -672 -725
rect -720 -755 -713 -729
rect -687 -742 -672 -729
rect -655 -742 -647 -725
rect -687 -750 -647 -742
rect -687 -755 -680 -750
rect -720 -762 -680 -755
<< via1 >>
rect -924 1547 -874 1732
rect -818 1546 -808 1726
rect -808 1546 -783 1726
rect -503 1546 -478 1726
rect -478 1546 -468 1726
rect -411 1547 -361 1732
rect -815 1487 -789 1513
rect -497 1487 -471 1513
rect -924 1185 -874 1370
rect -818 1192 -808 1367
rect -808 1192 -768 1367
rect -768 1192 -763 1367
rect -523 1192 -518 1367
rect -518 1192 -478 1367
rect -478 1192 -468 1367
rect -411 1185 -361 1370
rect -815 1130 -789 1156
rect -497 1130 -471 1156
rect 120 1007 330 1020
rect 720 1007 930 1020
rect 1320 1007 1530 1020
rect 1920 1007 2130 1020
rect 120 990 128 1007
rect 128 990 159 1007
rect 159 990 176 1007
rect 176 990 207 1007
rect 207 990 224 1007
rect 224 990 255 1007
rect 255 990 272 1007
rect 272 990 303 1007
rect 303 990 320 1007
rect 320 990 330 1007
rect 720 990 735 1007
rect 735 990 752 1007
rect 752 990 783 1007
rect 783 990 800 1007
rect 800 990 831 1007
rect 831 990 848 1007
rect 848 990 879 1007
rect 879 990 896 1007
rect 896 990 927 1007
rect 927 990 930 1007
rect 1320 990 1328 1007
rect 1328 990 1359 1007
rect 1359 990 1376 1007
rect 1376 990 1407 1007
rect 1407 990 1424 1007
rect 1424 990 1455 1007
rect 1455 990 1472 1007
rect 1472 990 1503 1007
rect 1503 990 1520 1007
rect 1520 990 1530 1007
rect 1920 990 1935 1007
rect 1935 990 1952 1007
rect 1952 990 1983 1007
rect 1983 990 2000 1007
rect 2000 990 2031 1007
rect 2031 990 2048 1007
rect 2048 990 2079 1007
rect 2079 990 2096 1007
rect 2096 990 2127 1007
rect 2127 990 2130 1007
rect 120 980 330 990
rect 720 980 930 990
rect 1320 980 1530 990
rect 1920 980 2130 990
rect -1424 821 -1398 825
rect -1424 804 -1419 821
rect -1419 804 -1402 821
rect -1402 804 -1398 821
rect -1424 799 -1398 804
rect -1388 821 -1362 825
rect -1388 804 -1383 821
rect -1383 804 -1366 821
rect -1366 804 -1362 821
rect -1388 799 -1362 804
rect -978 744 -788 864
rect -621 729 -595 733
rect -621 712 -616 729
rect -616 712 -599 729
rect -599 712 -595 729
rect -621 707 -595 712
rect -230 674 -20 690
rect 420 674 630 680
rect 1020 674 1230 680
rect 1620 674 1830 680
rect 2220 674 2430 680
rect -230 657 -224 674
rect -224 657 -207 674
rect -207 657 -176 674
rect -176 657 -159 674
rect -159 657 -128 674
rect -128 657 -111 674
rect -111 657 -80 674
rect -80 657 -63 674
rect -63 657 -32 674
rect -32 657 -20 674
rect 420 657 447 674
rect 447 657 464 674
rect 464 657 495 674
rect 495 657 512 674
rect 512 657 543 674
rect 543 657 560 674
rect 560 657 591 674
rect 591 657 608 674
rect 608 657 630 674
rect 1020 657 1023 674
rect 1023 657 1040 674
rect 1040 657 1071 674
rect 1071 657 1088 674
rect 1088 657 1119 674
rect 1119 657 1136 674
rect 1136 657 1167 674
rect 1167 657 1184 674
rect 1184 657 1215 674
rect 1215 657 1230 674
rect 1620 657 1647 674
rect 1647 657 1664 674
rect 1664 657 1695 674
rect 1695 657 1712 674
rect 1712 657 1743 674
rect 1743 657 1760 674
rect 1760 657 1791 674
rect 1791 657 1808 674
rect 1808 657 1830 674
rect 2220 657 2223 674
rect 2223 657 2240 674
rect 2240 657 2271 674
rect 2271 657 2288 674
rect 2288 657 2319 674
rect 2319 657 2336 674
rect 2336 657 2367 674
rect 2367 657 2384 674
rect 2384 657 2415 674
rect 2415 657 2430 674
rect -230 650 -20 657
rect 420 650 630 657
rect 1020 650 1230 657
rect 1620 650 1830 657
rect 2220 650 2430 657
rect -621 620 -595 624
rect -621 603 -616 620
rect -616 603 -599 620
rect -599 603 -595 620
rect -621 598 -595 603
rect -1424 528 -1398 532
rect -1424 511 -1419 528
rect -1419 511 -1402 528
rect -1402 511 -1398 528
rect -1424 506 -1398 511
rect -1388 528 -1362 532
rect -1388 511 -1383 528
rect -1383 511 -1366 528
rect -1366 511 -1362 528
rect -1388 506 -1362 511
rect -978 468 -788 588
rect -522 524 -496 529
rect -522 507 -518 524
rect -518 507 -501 524
rect -501 507 -496 524
rect -522 503 -496 507
rect -384 536 -358 540
rect -384 519 -379 536
rect -379 519 -362 536
rect -362 519 -358 536
rect -384 514 -358 519
rect -327 537 -301 541
rect -327 520 -322 537
rect -322 520 -305 537
rect -305 520 -301 537
rect -327 515 -301 520
rect -130 530 -104 535
rect -130 513 -126 530
rect -126 513 -109 530
rect -109 513 -104 530
rect -130 509 -104 513
rect 454 523 480 527
rect 454 506 458 523
rect 458 506 475 523
rect 475 506 480 523
rect 454 501 480 506
rect -184 443 -158 448
rect -184 426 -180 443
rect -180 426 -163 443
rect -163 426 -158 443
rect -184 422 -158 426
rect -83 407 -57 412
rect -83 390 -79 407
rect -79 390 -62 407
rect -62 390 -57 407
rect -83 386 -57 390
rect 1493 507 1519 511
rect 1493 490 1498 507
rect 1498 490 1515 507
rect 1515 490 1519 507
rect 1493 485 1519 490
rect 2136 523 2162 527
rect 2136 506 2141 523
rect 2141 506 2158 523
rect 2158 506 2162 523
rect 2136 501 2162 506
rect 2172 523 2198 527
rect 2172 506 2177 523
rect 2177 506 2194 523
rect 2194 506 2198 523
rect 2172 501 2198 506
rect 2330 523 2356 527
rect 2330 506 2334 523
rect 2334 506 2351 523
rect 2351 506 2356 523
rect 2330 501 2356 506
rect 2366 523 2392 527
rect 2366 506 2370 523
rect 2370 506 2387 523
rect 2387 506 2392 523
rect 2366 501 2392 506
rect 1835 471 1861 476
rect 1835 454 1840 471
rect 1840 454 1857 471
rect 1857 454 1861 471
rect 1835 450 1861 454
rect 1835 435 1861 440
rect 1835 418 1840 435
rect 1840 418 1857 435
rect 1857 418 1861 435
rect 1835 414 1861 418
rect 120 341 330 350
rect 720 341 930 350
rect 1320 341 1530 350
rect 1920 341 2130 350
rect 120 324 128 341
rect 128 324 159 341
rect 159 324 176 341
rect 176 324 207 341
rect 207 324 224 341
rect 224 324 255 341
rect 255 324 272 341
rect 272 324 303 341
rect 303 324 320 341
rect 320 324 330 341
rect 720 324 735 341
rect 735 324 752 341
rect 752 324 783 341
rect 783 324 800 341
rect 800 324 831 341
rect 831 324 848 341
rect 848 324 879 341
rect 879 324 896 341
rect 896 324 927 341
rect 927 324 930 341
rect 1320 324 1328 341
rect 1328 324 1359 341
rect 1359 324 1376 341
rect 1376 324 1407 341
rect 1407 324 1424 341
rect 1424 324 1455 341
rect 1455 324 1472 341
rect 1472 324 1503 341
rect 1503 324 1520 341
rect 1520 324 1530 341
rect 1920 324 1935 341
rect 1935 324 1952 341
rect 1952 324 1983 341
rect 1983 324 2000 341
rect 2000 324 2031 341
rect 2031 324 2048 341
rect 2048 324 2079 341
rect 2079 324 2096 341
rect 2096 324 2127 341
rect 2127 324 2130 341
rect 120 320 330 324
rect 720 320 930 324
rect 1320 320 1530 324
rect 1920 320 2130 324
rect -848 155 -822 159
rect -848 138 -843 155
rect -843 138 -826 155
rect -826 138 -822 155
rect -848 133 -822 138
rect -812 155 -786 159
rect -812 138 -807 155
rect -807 138 -790 155
rect -790 138 -786 155
rect -812 133 -786 138
rect -402 78 -212 198
rect 1632 245 1658 249
rect 1632 228 1637 245
rect 1637 228 1654 245
rect 1654 228 1658 245
rect 1632 223 1658 228
rect 1632 209 1658 213
rect 1632 192 1637 209
rect 1637 192 1654 209
rect 1654 192 1658 209
rect 1632 187 1658 192
rect 1837 243 1863 247
rect 1837 226 1841 243
rect 1841 226 1858 243
rect 1858 226 1863 243
rect 1837 221 1863 226
rect 1837 207 1863 211
rect 1837 190 1841 207
rect 1841 190 1858 207
rect 1858 190 1863 207
rect 1837 185 1863 190
rect 248 171 274 175
rect 248 154 252 171
rect 252 154 269 171
rect 269 154 274 171
rect 248 149 274 154
rect 456 160 482 164
rect 456 143 460 160
rect 460 143 477 160
rect 477 143 482 160
rect 456 138 482 143
rect 1494 176 1520 181
rect 1494 159 1499 176
rect 1499 159 1516 176
rect 1516 159 1520 176
rect 1494 155 1520 159
rect 2126 170 2152 175
rect 2126 153 2131 170
rect 2131 153 2148 170
rect 2148 153 2152 170
rect 2126 149 2152 153
rect 2189 167 2215 171
rect 2189 150 2193 167
rect 2193 150 2210 167
rect 2210 150 2215 167
rect 2189 145 2215 150
rect -45 63 -19 67
rect -45 46 -40 63
rect -40 46 -23 63
rect -23 46 -19 63
rect -45 41 -19 46
rect 420 8 630 10
rect 1020 8 1230 10
rect 1620 8 1830 10
rect 2220 8 2430 10
rect 420 -8 447 8
rect 447 -8 464 8
rect 464 -8 495 8
rect 495 -8 512 8
rect 512 -8 543 8
rect 543 -8 560 8
rect 560 -8 591 8
rect 591 -8 608 8
rect 608 -8 630 8
rect 1020 -8 1023 8
rect 1023 -8 1040 8
rect 1040 -8 1071 8
rect 1071 -8 1088 8
rect 1088 -8 1119 8
rect 1119 -8 1136 8
rect 1136 -8 1167 8
rect 1167 -8 1184 8
rect 1184 -8 1215 8
rect 1215 -8 1230 8
rect 1620 -8 1647 8
rect 1647 -8 1664 8
rect 1664 -8 1695 8
rect 1695 -8 1712 8
rect 1712 -8 1743 8
rect 1743 -8 1760 8
rect 1760 -8 1791 8
rect 1791 -8 1808 8
rect 1808 -8 1830 8
rect 2220 -8 2223 8
rect 2223 -8 2240 8
rect 2240 -8 2271 8
rect 2271 -8 2288 8
rect 2288 -8 2319 8
rect 2319 -8 2336 8
rect 2336 -8 2367 8
rect 2367 -8 2384 8
rect 2384 -8 2415 8
rect 2415 -8 2430 8
rect 420 -20 630 -8
rect 1020 -20 1230 -8
rect 1620 -20 1830 -8
rect 2220 -20 2430 -8
rect -719 -339 -694 -159
rect -694 -339 -684 -159
rect -628 -337 -578 -152
rect -713 -398 -687 -372
rect -739 -693 -734 -518
rect -734 -693 -694 -518
rect -694 -693 -684 -518
rect -628 -699 -578 -514
rect -713 -755 -687 -729
<< metal2 >>
rect -929 1732 -869 1737
rect -929 1547 -924 1732
rect -874 1547 -869 1732
rect -416 1732 -356 1737
rect -929 1542 -869 1547
rect -823 1726 -778 1731
rect -823 1546 -818 1726
rect -783 1546 -778 1726
rect -823 1541 -778 1546
rect -508 1726 -463 1731
rect -508 1546 -503 1726
rect -468 1546 -463 1726
rect -508 1541 -463 1546
rect -416 1547 -411 1732
rect -361 1547 -356 1732
rect -416 1542 -356 1547
rect -1140 1513 -464 1520
rect -1140 1487 -815 1513
rect -789 1487 -497 1513
rect -471 1487 -464 1513
rect -1140 1480 -464 1487
rect -1460 825 -1410 830
rect -1460 799 -1424 825
rect -1398 799 -1388 825
rect -1362 799 -1359 825
rect -1460 790 -1410 799
rect -1470 532 -1420 540
rect -1470 506 -1424 532
rect -1398 506 -1388 532
rect -1362 506 -1359 532
rect -1470 500 -1420 506
rect -1140 90 -1100 1480
rect -929 1370 -869 1375
rect -929 1185 -924 1370
rect -874 1185 -869 1370
rect -823 1367 -758 1372
rect -823 1192 -818 1367
rect -763 1192 -758 1367
rect -823 1187 -758 1192
rect -528 1367 -463 1372
rect -528 1192 -523 1367
rect -468 1192 -463 1367
rect -528 1187 -463 1192
rect -416 1370 -356 1375
rect -929 1180 -869 1185
rect -416 1185 -411 1370
rect -361 1185 -356 1370
rect -416 1180 -356 1185
rect -1160 80 -1100 90
rect -1160 40 -1150 80
rect -1110 40 -1100 80
rect -1160 30 -1100 40
rect -1140 -730 -1100 30
rect -1070 1156 -464 1163
rect -1070 1130 -815 1156
rect -789 1130 -497 1156
rect -471 1130 -464 1156
rect -1070 1123 -464 1130
rect -1070 0 -1030 1123
rect 110 1020 340 1030
rect 110 980 120 1020
rect 330 980 340 1020
rect 110 970 340 980
rect 710 1020 940 1030
rect 710 980 720 1020
rect 930 980 940 1020
rect 710 970 940 980
rect 1310 1020 1540 1030
rect 1310 980 1320 1020
rect 1530 980 1540 1020
rect 1310 970 1540 980
rect 1910 1020 2140 1030
rect 1910 980 1920 1020
rect 2130 980 2140 1020
rect 1910 970 2140 980
rect -983 864 -783 869
rect -983 860 -978 864
rect -983 750 -980 860
rect -983 744 -978 750
rect -788 744 -783 864
rect -983 739 -783 744
rect -621 733 -595 739
rect -595 719 -570 730
rect -595 707 -306 719
rect -621 704 -306 707
rect -621 624 -595 627
rect -595 619 -570 624
rect -595 604 -363 619
rect -595 598 -570 604
rect -621 593 -595 598
rect -983 588 -783 593
rect -983 580 -978 588
rect -983 470 -980 580
rect -983 468 -978 470
rect -788 468 -783 588
rect -983 463 -783 468
rect -572 564 -455 582
rect -746 275 -720 276
rect -572 275 -553 564
rect -525 503 -522 529
rect -496 503 -493 529
rect -522 485 -496 503
rect -473 488 -455 564
rect -378 540 -363 604
rect -321 541 -306 704
rect -240 690 -10 700
rect -240 650 -230 690
rect -20 650 -10 690
rect -240 640 -10 650
rect 410 680 640 690
rect 410 640 420 680
rect 630 640 640 680
rect 410 630 640 640
rect 1010 680 1240 690
rect 1010 640 1020 680
rect 1230 640 1240 680
rect 1010 630 1240 640
rect 1610 680 1840 690
rect 1610 640 1620 680
rect 1830 640 1840 680
rect 1610 630 1840 640
rect 2210 680 2440 690
rect 2210 640 2220 680
rect 2430 640 2440 680
rect 2210 630 2440 640
rect 383 550 1516 570
rect -387 514 -384 540
rect -358 514 -355 540
rect -330 515 -327 541
rect -301 515 -298 541
rect -133 509 -130 535
rect -104 509 -101 535
rect -129 488 -111 509
rect -519 290 -498 485
rect -473 470 -111 488
rect 383 454 403 550
rect 451 520 454 527
rect -187 448 403 454
rect -187 422 -184 448
rect -158 434 403 448
rect 428 501 454 520
rect 480 501 483 527
rect 1496 511 1516 550
rect 2024 553 2357 572
rect -158 422 -155 434
rect 428 415 447 501
rect 1490 485 1493 511
rect 1519 485 1522 511
rect -83 412 447 415
rect -57 396 447 412
rect 1835 476 1861 479
rect 1861 471 1870 476
rect 2024 471 2043 553
rect 2338 527 2357 553
rect 2133 501 2136 527
rect 2162 501 2172 527
rect 2198 501 2201 527
rect 2327 501 2330 527
rect 2356 501 2366 527
rect 2392 501 2395 527
rect 1861 453 2043 471
rect 1861 450 1870 453
rect 1835 440 1861 450
rect 1835 411 1861 414
rect -83 383 -57 386
rect 110 360 340 370
rect 110 320 120 360
rect 330 320 340 360
rect 110 310 340 320
rect 710 360 940 370
rect 710 320 720 360
rect 930 320 940 360
rect 710 310 940 320
rect 1310 360 1540 370
rect 1310 320 1320 360
rect 1530 320 1540 360
rect 1310 310 1540 320
rect 1910 360 2140 370
rect 1910 320 1920 360
rect 2130 320 2140 360
rect 1910 310 2140 320
rect -746 249 -550 275
rect -519 270 1685 290
rect -990 170 -930 180
rect -990 130 -980 170
rect -940 159 -820 170
rect -746 159 -720 249
rect -940 133 -848 159
rect -822 133 -812 159
rect -786 133 -720 159
rect -410 200 -200 210
rect -410 198 -400 200
rect -940 130 -820 133
rect -990 120 -930 130
rect -410 78 -402 198
rect -210 80 -200 200
rect 251 175 271 270
rect 1632 249 1685 270
rect 1658 223 1685 249
rect 1632 213 1685 223
rect 1658 208 1685 213
rect 1837 247 1863 250
rect 1837 211 1863 221
rect 2165 211 2181 501
rect 1658 187 1797 208
rect 1632 184 1658 187
rect 245 149 248 175
rect 274 149 277 175
rect 453 162 456 164
rect -212 78 -200 80
rect -410 70 -200 78
rect 392 138 456 162
rect 482 138 485 164
rect 1491 155 1494 181
rect 1520 155 1523 181
rect -45 67 -19 73
rect 392 65 416 138
rect 1491 137 1523 155
rect 1774 163 1795 187
rect 1863 195 2181 211
rect 1863 185 1879 195
rect 1837 182 1863 185
rect 2102 175 2155 178
rect 2102 163 2126 175
rect 1774 149 2126 163
rect 2152 149 2155 175
rect 2350 171 2366 501
rect 1774 145 2155 149
rect 2186 145 2189 171
rect 2215 145 2366 171
rect 1774 143 2102 145
rect -19 41 416 65
rect -45 38 -19 41
rect 410 10 640 20
rect -1070 -10 -1010 0
rect -1070 -50 -1060 -10
rect -1020 -50 -1010 -10
rect 410 -30 420 10
rect 630 -30 640 10
rect 410 -40 640 -30
rect 1010 10 1240 20
rect 1010 -30 1020 10
rect 1230 -30 1240 10
rect 1010 -40 1240 -30
rect 1610 10 1840 20
rect 1610 -30 1620 10
rect 1830 -30 1840 10
rect 1610 -40 1840 -30
rect 2210 10 2440 20
rect 2210 -30 2220 10
rect 2430 -30 2440 10
rect 2210 -40 2440 -30
rect -1070 -60 -1010 -50
rect -1070 -370 -1030 -60
rect -633 -152 -573 -147
rect -724 -159 -679 -154
rect -724 -339 -719 -159
rect -684 -339 -679 -159
rect -724 -344 -679 -339
rect -633 -337 -628 -152
rect -578 -337 -573 -152
rect -633 -342 -573 -337
rect -720 -367 -680 -365
rect -723 -370 -680 -367
rect -1070 -372 -680 -370
rect -1070 -398 -713 -372
rect -687 -398 -680 -372
rect -1070 -405 -680 -398
rect -1070 -410 -720 -405
rect -744 -518 -679 -513
rect -744 -693 -739 -518
rect -684 -693 -679 -518
rect -744 -698 -679 -693
rect -633 -514 -573 -509
rect -633 -699 -628 -514
rect -578 -699 -573 -514
rect -633 -704 -573 -699
rect -720 -724 -680 -722
rect -723 -729 -680 -724
rect -723 -730 -713 -729
rect -1140 -755 -713 -730
rect -687 -755 -680 -729
rect -1140 -762 -680 -755
rect -1140 -770 -690 -762
<< via2 >>
rect -924 1547 -874 1732
rect -813 1546 -783 1726
rect -503 1546 -473 1726
rect -411 1547 -361 1732
rect -924 1185 -874 1370
rect -813 1192 -763 1367
rect -523 1192 -473 1367
rect -411 1185 -361 1370
rect -1150 40 -1110 80
rect 120 980 330 1020
rect 720 980 930 1020
rect 1320 980 1530 1020
rect 1920 980 2130 1020
rect -980 750 -978 860
rect -978 750 -790 860
rect -980 470 -978 580
rect -978 470 -790 580
rect -230 650 -20 690
rect 420 650 630 680
rect 420 640 630 650
rect 1020 650 1230 680
rect 1020 640 1230 650
rect 1620 650 1830 680
rect 1620 640 1830 650
rect 2220 650 2430 680
rect 2220 640 2430 650
rect 120 350 330 360
rect 120 320 330 350
rect 720 350 930 360
rect 720 320 930 350
rect 1320 350 1530 360
rect 1320 320 1530 350
rect 1920 350 2130 360
rect 1920 320 2130 350
rect -980 130 -940 170
rect -400 198 -210 200
rect -400 80 -212 198
rect -212 80 -210 198
rect -1060 -50 -1020 -10
rect 420 -20 630 10
rect 420 -30 630 -20
rect 1020 -20 1230 10
rect 1020 -30 1230 -20
rect 1620 -20 1830 10
rect 1620 -30 1830 -20
rect 2220 -20 2430 10
rect 2220 -30 2430 -20
rect -719 -339 -689 -159
rect -628 -337 -578 -152
rect -739 -693 -689 -518
rect -628 -699 -578 -514
<< metal3 >>
rect -1864 1732 -849 1737
rect -1864 1717 -924 1732
rect -874 1717 -849 1732
rect -1864 1557 -989 1717
rect -869 1557 -849 1717
rect -1864 1547 -924 1557
rect -874 1547 -849 1557
rect -1864 1540 -849 1547
rect -818 1726 -468 1736
rect -818 1546 -813 1726
rect -783 1666 -503 1726
rect -783 1616 -778 1666
rect -710 1616 -630 1666
rect -508 1616 -503 1666
rect -783 1546 -503 1616
rect -473 1546 -468 1726
rect -818 1541 -778 1546
rect -2649 1370 -849 1380
rect -710 1377 -630 1546
rect -508 1541 -468 1546
rect -436 1732 578 1737
rect -436 1717 -411 1732
rect -361 1717 578 1732
rect -436 1557 -416 1717
rect -296 1557 578 1717
rect -436 1547 -411 1557
rect -361 1547 578 1557
rect -436 1540 578 1547
rect -2649 1360 -924 1370
rect -874 1360 -849 1370
rect -2649 1200 -989 1360
rect -869 1200 -849 1360
rect -2649 1185 -924 1200
rect -874 1185 -849 1200
rect -818 1367 -468 1377
rect -818 1192 -813 1367
rect -763 1307 -523 1367
rect -763 1257 -758 1307
rect -710 1257 -630 1307
rect -528 1257 -523 1307
rect -763 1192 -523 1257
rect -473 1192 -468 1367
rect -818 1187 -468 1192
rect -436 1370 1363 1380
rect -436 1360 -411 1370
rect -361 1360 1363 1370
rect -436 1200 -416 1360
rect -296 1200 1363 1360
rect -2649 1183 -849 1185
rect -929 1180 -869 1183
rect -990 860 -780 870
rect -990 750 -980 860
rect -790 750 -780 860
rect -990 740 -780 750
rect -710 710 -630 1187
rect -436 1185 -411 1200
rect -361 1185 1363 1200
rect -436 1183 1363 1185
rect -416 1180 -356 1183
rect 110 1020 2140 1030
rect 110 980 120 1020
rect 330 980 720 1020
rect 930 980 1320 1020
rect 1530 980 1920 1020
rect 2130 980 2140 1020
rect 110 970 2140 980
rect -710 690 20 710
rect -710 650 -230 690
rect -20 650 20 690
rect -710 630 20 650
rect -990 580 -780 590
rect -990 470 -980 580
rect -790 470 -780 580
rect -990 460 -780 470
rect -710 410 -630 630
rect -890 330 -630 410
rect 110 370 170 970
rect 280 370 340 970
rect 110 360 340 370
rect -1240 170 -930 180
rect -1240 130 -980 170
rect -940 130 -930 170
rect -1240 120 -930 130
rect -1240 80 -1100 90
rect -1240 40 -1150 80
rect -1110 40 -1100 80
rect -1240 30 -1100 40
rect -890 20 -810 330
rect 110 320 120 360
rect 330 320 340 360
rect 110 310 340 320
rect 410 680 640 690
rect 410 640 420 680
rect 630 640 640 680
rect 410 630 640 640
rect -410 200 -200 210
rect -410 80 -400 200
rect -210 80 -200 200
rect -410 70 -200 80
rect 410 20 470 630
rect 580 20 640 630
rect 710 370 770 970
rect 880 370 940 970
rect 710 360 940 370
rect 710 320 720 360
rect 930 320 940 360
rect 710 310 940 320
rect 1010 680 1240 690
rect 1010 640 1020 680
rect 1230 640 1240 680
rect 1010 630 1240 640
rect 1010 20 1070 630
rect 1180 20 1240 630
rect 1310 370 1370 970
rect 1480 370 1540 970
rect 1310 360 1540 370
rect 1310 320 1320 360
rect 1530 320 1540 360
rect 1310 310 1540 320
rect 1610 680 1840 690
rect 1610 640 1620 680
rect 1830 640 1840 680
rect 1610 630 1840 640
rect 1610 20 1670 630
rect 1780 20 1840 630
rect 1910 370 1970 970
rect 2080 370 2140 970
rect 1910 360 2140 370
rect 1910 320 1920 360
rect 2130 320 2140 360
rect 1910 310 2140 320
rect 2210 680 2440 690
rect 2210 640 2220 680
rect 2430 640 2440 680
rect 2210 630 2440 640
rect 2210 20 2270 630
rect 2380 20 2440 630
rect -890 10 2440 20
rect -1240 -10 -1010 0
rect -1240 -50 -1060 -10
rect -1020 -50 -1010 -10
rect -1240 -60 -1010 -50
rect -890 -30 420 10
rect 630 -30 1020 10
rect 1230 -30 1620 10
rect 1830 -30 2220 10
rect 2430 -30 2440 10
rect -890 -40 2440 -30
rect -890 -149 -810 -40
rect -890 -159 -684 -149
rect -890 -219 -719 -159
rect -890 -269 -810 -219
rect -724 -269 -719 -219
rect -890 -339 -719 -269
rect -689 -339 -684 -159
rect -890 -508 -810 -339
rect -724 -344 -684 -339
rect -653 -152 362 -147
rect -653 -167 -628 -152
rect -578 -167 362 -152
rect -653 -327 -633 -167
rect -513 -327 362 -167
rect -653 -337 -628 -327
rect -578 -337 362 -327
rect -653 -344 362 -337
rect -890 -518 -684 -508
rect -890 -578 -739 -518
rect -890 -628 -810 -578
rect -744 -628 -739 -578
rect -890 -693 -739 -628
rect -689 -693 -684 -518
rect -890 -698 -684 -693
rect -653 -514 1147 -504
rect -653 -524 -628 -514
rect -578 -524 1147 -514
rect -653 -684 -633 -524
rect -513 -684 1147 -524
rect -890 -790 -810 -698
rect -653 -699 -628 -684
rect -578 -699 1147 -684
rect -653 -701 1147 -699
rect -633 -704 -573 -701
<< via3 >>
rect -989 1557 -924 1717
rect -924 1557 -874 1717
rect -874 1557 -869 1717
rect -416 1557 -411 1717
rect -411 1557 -361 1717
rect -361 1557 -296 1717
rect -989 1200 -924 1360
rect -924 1200 -874 1360
rect -874 1200 -869 1360
rect -416 1200 -411 1360
rect -411 1200 -361 1360
rect -361 1200 -296 1360
rect -980 750 -790 860
rect -980 470 -790 580
rect -400 80 -210 200
rect -633 -327 -628 -167
rect -628 -327 -578 -167
rect -578 -327 -513 -167
rect -633 -684 -628 -524
rect -628 -684 -578 -524
rect -578 -684 -513 -524
<< mimcap >>
rect -1844 1707 -1059 1717
rect -1844 1567 -1834 1707
rect -1069 1567 -1059 1707
rect -1844 1557 -1059 1567
rect -226 1707 558 1717
rect -226 1567 -216 1707
rect 548 1567 558 1707
rect -226 1557 558 1567
rect -2629 1350 -1059 1360
rect -2629 1210 -2619 1350
rect -1069 1210 -1059 1350
rect -2629 1200 -1059 1210
rect -226 1350 1343 1360
rect -226 1210 -216 1350
rect 1333 1210 1343 1350
rect -226 1200 1343 1210
rect -443 -177 342 -167
rect -443 -317 -433 -177
rect 332 -317 342 -177
rect -443 -327 342 -317
rect -443 -534 1127 -524
rect -443 -674 -433 -534
rect 1117 -674 1127 -534
rect -443 -684 1127 -674
<< mimcapcontact >>
rect -1834 1567 -1069 1707
rect -216 1567 548 1707
rect -2619 1210 -1069 1350
rect -216 1210 1333 1350
rect -433 -317 332 -177
rect -433 -674 1117 -534
<< metal4 >>
rect -1864 1732 -1039 1737
rect -1869 1707 -1039 1732
rect -1869 1567 -1834 1707
rect -1069 1567 -1039 1707
rect -1869 1542 -1039 1567
rect -1864 1540 -1039 1542
rect -1009 1717 -849 1737
rect -1009 1557 -989 1717
rect -869 1557 -849 1717
rect -1009 1540 -849 1557
rect -436 1717 -276 1737
rect -436 1557 -416 1717
rect -296 1557 -276 1717
rect -436 1540 -276 1557
rect -246 1732 578 1737
rect -246 1707 583 1732
rect -246 1567 -216 1707
rect 548 1567 583 1707
rect -246 1542 583 1567
rect -246 1540 578 1542
rect -1200 1380 -1100 1540
rect -180 1380 -80 1540
rect -2649 1375 -1039 1380
rect -2654 1350 -1039 1375
rect -2654 1210 -2619 1350
rect -1069 1210 -1039 1350
rect -2654 1185 -1039 1210
rect -2649 1183 -1039 1185
rect -1009 1360 -849 1380
rect -1009 1200 -989 1360
rect -869 1200 -849 1360
rect -1009 1183 -849 1200
rect -436 1360 -276 1380
rect -436 1200 -416 1360
rect -296 1200 -276 1360
rect -436 1183 -276 1200
rect -246 1375 1363 1380
rect -246 1350 1368 1375
rect -246 1210 -216 1350
rect 1333 1210 1368 1350
rect -246 1185 1368 1210
rect -246 1183 1363 1185
rect -1200 600 -1100 1183
rect -180 880 -80 1183
rect -1000 860 -80 880
rect -1000 750 -980 860
rect -790 780 -80 860
rect -790 750 -750 780
rect -1000 730 -750 750
rect -1200 580 -750 600
rect -1200 500 -980 580
rect -1000 470 -980 500
rect -790 470 -750 580
rect -1000 450 -750 470
rect -410 200 -200 210
rect -410 80 -400 200
rect -210 80 -200 200
rect -410 70 -200 80
rect -340 -147 -240 70
rect -653 -167 -493 -147
rect -653 -327 -633 -167
rect -513 -327 -493 -167
rect -653 -344 -493 -327
rect -463 -152 362 -147
rect -463 -177 367 -152
rect -463 -317 -433 -177
rect 332 -317 367 -177
rect -463 -342 367 -317
rect -463 -344 362 -342
rect -340 -504 -240 -344
rect -653 -524 -493 -504
rect -653 -684 -633 -524
rect -513 -684 -493 -524
rect -653 -701 -493 -684
rect -463 -509 1147 -504
rect -463 -534 1152 -509
rect -463 -674 -433 -534
rect 1117 -674 1152 -534
rect -463 -699 1152 -674
rect -463 -701 1147 -699
<< via4 >>
rect -989 1557 -869 1717
rect -416 1557 -296 1717
rect -989 1200 -869 1360
rect -416 1200 -296 1360
rect -633 -327 -513 -167
rect -633 -684 -513 -524
<< mimcap2 >>
rect -1844 1707 -1059 1717
rect -1844 1567 -1834 1707
rect -1069 1567 -1059 1707
rect -1844 1557 -1059 1567
rect -226 1707 558 1717
rect -226 1567 -216 1707
rect 548 1567 558 1707
rect -226 1557 558 1567
rect -2629 1350 -1059 1360
rect -2629 1210 -2619 1350
rect -1069 1210 -1059 1350
rect -2629 1200 -1059 1210
rect -226 1350 1343 1360
rect -226 1210 -216 1350
rect 1333 1210 1343 1350
rect -226 1200 1343 1210
rect -443 -177 342 -167
rect -443 -317 -433 -177
rect 332 -317 342 -177
rect -443 -327 342 -317
rect -443 -534 1127 -524
rect -443 -674 -433 -534
rect 1117 -674 1127 -534
rect -443 -684 1127 -674
<< mimcap2contact >>
rect -1834 1567 -1069 1707
rect -216 1567 548 1707
rect -2619 1210 -1069 1350
rect -216 1210 1333 1350
rect -433 -317 332 -177
rect -433 -674 1117 -534
<< metal5 >>
rect -1864 1717 -849 1737
rect -1864 1707 -989 1717
rect -1864 1567 -1834 1707
rect -1069 1567 -989 1707
rect -1864 1557 -989 1567
rect -869 1557 -849 1717
rect -1864 1540 -849 1557
rect -436 1717 578 1737
rect -436 1557 -416 1717
rect -296 1707 578 1717
rect -296 1567 -216 1707
rect 548 1567 578 1707
rect -296 1557 578 1567
rect -436 1540 578 1557
rect -2649 1360 -849 1380
rect -2649 1350 -989 1360
rect -2649 1210 -2619 1350
rect -1069 1210 -989 1350
rect -2649 1200 -989 1210
rect -869 1200 -849 1360
rect -2649 1183 -849 1200
rect -436 1360 1363 1380
rect -436 1200 -416 1360
rect -296 1350 1363 1360
rect -296 1210 -216 1350
rect 1333 1210 1363 1350
rect -296 1200 1363 1210
rect -436 1183 1363 1200
rect -653 -167 362 -147
rect -653 -327 -633 -167
rect -513 -177 362 -167
rect -513 -317 -433 -177
rect 332 -317 362 -177
rect -513 -327 362 -317
rect -653 -344 362 -327
rect -653 -524 1147 -504
rect -653 -684 -633 -524
rect -513 -534 1147 -524
rect -513 -674 -433 -534
rect 1117 -674 1147 -534
rect -513 -684 1147 -674
rect -653 -701 1147 -684
<< res1p41 >>
rect -1043 732 -991 875
rect -1043 456 -991 599
rect -467 66 -415 209
<< labels >>
rlabel metal2 1860 185 1879 211 1 UPDN
rlabel metal3 -1240 120 -1210 180 1 CLKIN
rlabel metal2 -1470 500 -1420 540 1 A0
rlabel metal2 -1460 790 -1410 830 1 A1
rlabel locali 2450 500 2470 540 1 GP
rlabel metal2 1491 137 1523 181 1 RSTB
rlabel metal3 360 1018 394 1030 1 VHI
rlabel metal3 -219 698 -185 709 1 VLO
rlabel metal3 -1240 30 -1210 90 1 C100
rlabel metal3 -1240 -60 -1210 0 1 C50
rlabel metal2 1 435 16 453 1 MUX_OUT
rlabel metal2 90 396 105 414 1 ENCLK
rlabel locali 2467 132 2487 172 1 GN
rlabel metal2 87 46 104 60 1 UDCLK
<< end >>
