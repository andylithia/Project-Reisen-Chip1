magic
tech sky130A
magscale 1 2
timestamp 1671673121
<< poly >>
rect -3066 94 -3004 103
rect -3066 60 -3052 94
rect -3018 60 -3004 94
rect -3066 51 -3004 60
rect -3000 51 -2999 103
<< locali >>
rect -3067 94 -2931 103
rect -3067 60 -3052 94
rect -3018 60 -2980 94
rect -2946 60 -2931 94
rect -3067 51 -2931 60
rect -2845 52 -2703 111
rect -1801 28 -1566 94
rect -1451 78 -1387 87
rect -1451 44 -1436 78
rect -1402 44 -1387 78
rect -1451 35 -1387 44
rect -1455 -90 -1403 -70
rect -1455 -124 -1446 -90
rect -1412 -124 -1403 -90
rect -1455 -139 -1403 -124
<< viali >>
rect -3052 60 -3018 94
rect -2980 60 -2946 94
rect -1436 44 -1402 78
rect -1446 -124 -1412 -90
<< metal1 >>
rect -2890 242 -1386 308
rect -2890 125 -2824 242
rect -2994 103 -2824 125
rect -3067 51 -3061 103
rect -3009 51 -2989 103
rect -2937 59 -2824 103
rect -2937 51 -2931 59
rect -1452 78 -1386 242
rect -1452 44 -1436 78
rect -1402 44 -1386 78
rect -1452 28 -1386 44
rect -1455 -81 -1403 -70
rect -1455 -139 -1403 -133
<< via1 >>
rect -3061 94 -3009 103
rect -3061 60 -3052 94
rect -3052 60 -3018 94
rect -3018 60 -3009 94
rect -3061 51 -3009 60
rect -2989 94 -2937 103
rect -2989 60 -2980 94
rect -2980 60 -2946 94
rect -2946 60 -2937 94
rect -2989 51 -2937 60
rect -2170 -60 -1790 180
rect -1455 -90 -1403 -81
rect -1455 -124 -1446 -90
rect -1446 -124 -1412 -90
rect -1412 -124 -1403 -90
rect -1455 -133 -1403 -124
<< metal2 >>
rect -2180 180 -1780 190
rect -3067 51 -3061 103
rect -3009 51 -2989 103
rect -2937 51 -2931 103
rect -2180 -60 -2170 180
rect -1790 -60 -1780 180
rect -2180 -70 -1780 -60
rect -1455 -81 -1403 -70
rect -1455 -139 -1403 -133
use sky130_fd_pr__res_xhigh_po_1p41_GKKP9B  sky130_fd_pr__res_xhigh_po_1p41_GKKP9B_0
timestamp 1671381513
transform 0 1 -2247 -1 0 60
box -143 -482 143 482
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -2037 0 1 -216
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -2805 0 1 -216
box -38 -49 806 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -3093 0 1 -216
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_2 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -1653 0 1 -216
box -38 -49 326 715
<< labels >>
rlabel metal2 -3067 51 -3061 103 1 A
rlabel metal2 -2180 -70 -1780 -60 1 C
rlabel metal2 -1455 -80 -1403 -70 1 Y
<< end >>
