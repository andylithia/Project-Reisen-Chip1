RC circuit
v1 1 0 dc 0 ac 1
r1 1 2 1k 
c1 2 0 100n
r2 2 0 1MEG
.control
ac dec 10 10Hz 100kHz
display
print vdb(2) vp(2)> export-1.txt
.endc
.end
