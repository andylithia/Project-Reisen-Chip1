magic
tech sky130B
magscale 1 2
timestamp 1668574539
<< error_p >>
rect 1456 0 1524 30
rect 1460 -60 1520 -30
rect 1396 -1320 1440 -1060
rect 1456 -1380 1500 -1000
rect 4276 -1204 4284 -266
rect 4336 -1144 4344 -206
rect 4276 -1436 4284 -1360
rect 4336 -1436 4344 -1420
rect 4216 -1504 4336 -1480
rect 4180 -1564 4336 -1540
<< nwell >>
rect -20 1080 6072 2094
rect -20 -3514 6072 -2500
<< pwell >>
rect 12 924 6040 962
rect 12 890 353 924
rect 356 890 414 924
rect 419 890 2753 924
rect 2758 890 2816 924
rect 2819 890 3233 924
rect 3236 890 3294 924
rect 3299 890 5633 924
rect 5638 890 5696 924
rect 5699 890 6040 924
rect 12 306 6040 890
rect 12 -2310 6040 -1726
rect 12 -2344 353 -2310
rect 356 -2344 414 -2310
rect 419 -2344 2753 -2310
rect 2758 -2344 2816 -2310
rect 2819 -2344 3233 -2310
rect 3236 -2344 3294 -2310
rect 3299 -2344 5633 -2310
rect 5638 -2344 5696 -2310
rect 5699 -2344 6040 -2310
rect 12 -2382 6040 -2344
<< nmos >>
rect 83 452 113 852
rect 179 452 209 852
rect 275 452 305 852
rect 371 452 401 852
rect 467 452 497 852
rect 563 452 593 852
rect 659 452 689 852
rect 755 452 785 852
rect 851 452 881 852
rect 947 452 977 852
rect 1043 452 1073 852
rect 1139 452 1169 852
rect 1235 452 1265 852
rect 1331 452 1361 852
rect 1427 452 1457 852
rect 1523 452 1553 852
rect 1619 452 1649 852
rect 1715 452 1745 852
rect 1811 452 1841 852
rect 1907 452 1937 852
rect 2003 452 2033 852
rect 2099 452 2129 852
rect 2195 452 2225 852
rect 2291 452 2321 852
rect 2387 452 2417 852
rect 2483 452 2513 852
rect 2579 452 2609 852
rect 2675 452 2705 852
rect 2771 452 2801 852
rect 2867 452 2897 852
rect 2963 452 2993 852
rect 3059 452 3089 852
rect 3155 452 3185 852
rect 3251 452 3281 852
rect 3347 452 3377 852
rect 3443 452 3473 852
rect 3539 452 3569 852
rect 3635 452 3665 852
rect 3731 452 3761 852
rect 3827 452 3857 852
rect 3923 452 3953 852
rect 4019 452 4049 852
rect 4115 452 4145 852
rect 4211 452 4241 852
rect 4307 452 4337 852
rect 4403 452 4433 852
rect 4499 452 4529 852
rect 4595 452 4625 852
rect 4691 452 4721 852
rect 4787 452 4817 852
rect 4883 452 4913 852
rect 4979 452 5009 852
rect 5075 452 5105 852
rect 5171 452 5201 852
rect 5267 452 5297 852
rect 5363 452 5393 852
rect 5459 452 5489 852
rect 5555 452 5585 852
rect 5651 452 5681 852
rect 5747 452 5777 852
rect 5843 452 5873 852
rect 5939 452 5969 852
rect 83 -2272 113 -1872
rect 179 -2272 209 -1872
rect 275 -2272 305 -1872
rect 371 -2272 401 -1872
rect 467 -2272 497 -1872
rect 563 -2272 593 -1872
rect 659 -2272 689 -1872
rect 755 -2272 785 -1872
rect 851 -2272 881 -1872
rect 947 -2272 977 -1872
rect 1043 -2272 1073 -1872
rect 1139 -2272 1169 -1872
rect 1235 -2272 1265 -1872
rect 1331 -2272 1361 -1872
rect 1427 -2272 1457 -1872
rect 1523 -2272 1553 -1872
rect 1619 -2272 1649 -1872
rect 1715 -2272 1745 -1872
rect 1811 -2272 1841 -1872
rect 1907 -2272 1937 -1872
rect 2003 -2272 2033 -1872
rect 2099 -2272 2129 -1872
rect 2195 -2272 2225 -1872
rect 2291 -2272 2321 -1872
rect 2387 -2272 2417 -1872
rect 2483 -2272 2513 -1872
rect 2579 -2272 2609 -1872
rect 2675 -2272 2705 -1872
rect 2771 -2272 2801 -1872
rect 2867 -2272 2897 -1872
rect 2963 -2272 2993 -1872
rect 3059 -2272 3089 -1872
rect 3155 -2272 3185 -1872
rect 3251 -2272 3281 -1872
rect 3347 -2272 3377 -1872
rect 3443 -2272 3473 -1872
rect 3539 -2272 3569 -1872
rect 3635 -2272 3665 -1872
rect 3731 -2272 3761 -1872
rect 3827 -2272 3857 -1872
rect 3923 -2272 3953 -1872
rect 4019 -2272 4049 -1872
rect 4115 -2272 4145 -1872
rect 4211 -2272 4241 -1872
rect 4307 -2272 4337 -1872
rect 4403 -2272 4433 -1872
rect 4499 -2272 4529 -1872
rect 4595 -2272 4625 -1872
rect 4691 -2272 4721 -1872
rect 4787 -2272 4817 -1872
rect 4883 -2272 4913 -1872
rect 4979 -2272 5009 -1872
rect 5075 -2272 5105 -1872
rect 5171 -2272 5201 -1872
rect 5267 -2272 5297 -1872
rect 5363 -2272 5393 -1872
rect 5459 -2272 5489 -1872
rect 5555 -2272 5585 -1872
rect 5651 -2272 5681 -1872
rect 5747 -2272 5777 -1872
rect 5843 -2272 5873 -1872
rect 5939 -2272 5969 -1872
<< pmos >>
rect 83 1207 113 1927
rect 179 1207 209 1927
rect 275 1207 305 1927
rect 371 1207 401 1927
rect 467 1207 497 1927
rect 563 1207 593 1927
rect 659 1207 689 1927
rect 755 1207 785 1927
rect 851 1207 881 1927
rect 947 1207 977 1927
rect 1043 1207 1073 1927
rect 1139 1207 1169 1927
rect 1235 1207 1265 1927
rect 1331 1207 1361 1927
rect 1427 1207 1457 1927
rect 1523 1207 1553 1927
rect 1619 1207 1649 1927
rect 1715 1207 1745 1927
rect 1811 1207 1841 1927
rect 1907 1207 1937 1927
rect 2003 1207 2033 1927
rect 2099 1207 2129 1927
rect 2195 1207 2225 1927
rect 2291 1207 2321 1927
rect 2387 1207 2417 1927
rect 2483 1207 2513 1927
rect 2579 1207 2609 1927
rect 2675 1207 2705 1927
rect 2771 1207 2801 1927
rect 2867 1207 2897 1927
rect 2963 1207 2993 1927
rect 3059 1207 3089 1927
rect 3155 1207 3185 1927
rect 3251 1207 3281 1927
rect 3347 1207 3377 1927
rect 3443 1207 3473 1927
rect 3539 1207 3569 1927
rect 3635 1207 3665 1927
rect 3731 1207 3761 1927
rect 3827 1207 3857 1927
rect 3923 1207 3953 1927
rect 4019 1207 4049 1927
rect 4115 1207 4145 1927
rect 4211 1207 4241 1927
rect 4307 1207 4337 1927
rect 4403 1207 4433 1927
rect 4499 1207 4529 1927
rect 4595 1207 4625 1927
rect 4691 1207 4721 1927
rect 4787 1207 4817 1927
rect 4883 1207 4913 1927
rect 4979 1207 5009 1927
rect 5075 1207 5105 1927
rect 5171 1207 5201 1927
rect 5267 1207 5297 1927
rect 5363 1207 5393 1927
rect 5459 1207 5489 1927
rect 5555 1207 5585 1927
rect 5651 1207 5681 1927
rect 5747 1207 5777 1927
rect 5843 1207 5873 1927
rect 5939 1207 5969 1927
rect 83 -3347 113 -2627
rect 179 -3347 209 -2627
rect 275 -3347 305 -2627
rect 371 -3347 401 -2627
rect 467 -3347 497 -2627
rect 563 -3347 593 -2627
rect 659 -3347 689 -2627
rect 755 -3347 785 -2627
rect 851 -3347 881 -2627
rect 947 -3347 977 -2627
rect 1043 -3347 1073 -2627
rect 1139 -3347 1169 -2627
rect 1235 -3347 1265 -2627
rect 1331 -3347 1361 -2627
rect 1427 -3347 1457 -2627
rect 1523 -3347 1553 -2627
rect 1619 -3347 1649 -2627
rect 1715 -3347 1745 -2627
rect 1811 -3347 1841 -2627
rect 1907 -3347 1937 -2627
rect 2003 -3347 2033 -2627
rect 2099 -3347 2129 -2627
rect 2195 -3347 2225 -2627
rect 2291 -3347 2321 -2627
rect 2387 -3347 2417 -2627
rect 2483 -3347 2513 -2627
rect 2579 -3347 2609 -2627
rect 2675 -3347 2705 -2627
rect 2771 -3347 2801 -2627
rect 2867 -3347 2897 -2627
rect 2963 -3347 2993 -2627
rect 3059 -3347 3089 -2627
rect 3155 -3347 3185 -2627
rect 3251 -3347 3281 -2627
rect 3347 -3347 3377 -2627
rect 3443 -3347 3473 -2627
rect 3539 -3347 3569 -2627
rect 3635 -3347 3665 -2627
rect 3731 -3347 3761 -2627
rect 3827 -3347 3857 -2627
rect 3923 -3347 3953 -2627
rect 4019 -3347 4049 -2627
rect 4115 -3347 4145 -2627
rect 4211 -3347 4241 -2627
rect 4307 -3347 4337 -2627
rect 4403 -3347 4433 -2627
rect 4499 -3347 4529 -2627
rect 4595 -3347 4625 -2627
rect 4691 -3347 4721 -2627
rect 4787 -3347 4817 -2627
rect 4883 -3347 4913 -2627
rect 4979 -3347 5009 -2627
rect 5075 -3347 5105 -2627
rect 5171 -3347 5201 -2627
rect 5267 -3347 5297 -2627
rect 5363 -3347 5393 -2627
rect 5459 -3347 5489 -2627
rect 5555 -3347 5585 -2627
rect 5651 -3347 5681 -2627
rect 5747 -3347 5777 -2627
rect 5843 -3347 5873 -2627
rect 5939 -3347 5969 -2627
<< ndiff >>
rect 21 840 83 852
rect 21 464 33 840
rect 67 464 83 840
rect 21 452 83 464
rect 113 840 179 852
rect 113 464 129 840
rect 163 464 179 840
rect 113 452 179 464
rect 209 840 275 852
rect 209 464 225 840
rect 259 464 275 840
rect 209 452 275 464
rect 305 840 371 852
rect 305 464 321 840
rect 355 464 371 840
rect 305 452 371 464
rect 401 840 467 852
rect 401 464 417 840
rect 451 464 467 840
rect 401 452 467 464
rect 497 840 563 852
rect 497 464 513 840
rect 547 464 563 840
rect 497 452 563 464
rect 593 840 659 852
rect 593 464 609 840
rect 643 464 659 840
rect 593 452 659 464
rect 689 840 755 852
rect 689 464 705 840
rect 739 464 755 840
rect 689 452 755 464
rect 785 840 851 852
rect 785 464 801 840
rect 835 464 851 840
rect 785 452 851 464
rect 881 840 947 852
rect 881 464 897 840
rect 931 464 947 840
rect 881 452 947 464
rect 977 840 1043 852
rect 977 464 993 840
rect 1027 464 1043 840
rect 977 452 1043 464
rect 1073 840 1139 852
rect 1073 464 1089 840
rect 1123 464 1139 840
rect 1073 452 1139 464
rect 1169 840 1235 852
rect 1169 464 1185 840
rect 1219 464 1235 840
rect 1169 452 1235 464
rect 1265 840 1331 852
rect 1265 464 1281 840
rect 1315 464 1331 840
rect 1265 452 1331 464
rect 1361 840 1427 852
rect 1361 464 1377 840
rect 1411 464 1427 840
rect 1361 452 1427 464
rect 1457 840 1523 852
rect 1457 464 1473 840
rect 1507 464 1523 840
rect 1457 452 1523 464
rect 1553 840 1619 852
rect 1553 464 1569 840
rect 1603 464 1619 840
rect 1553 452 1619 464
rect 1649 840 1715 852
rect 1649 464 1665 840
rect 1699 464 1715 840
rect 1649 452 1715 464
rect 1745 840 1811 852
rect 1745 464 1761 840
rect 1795 464 1811 840
rect 1745 452 1811 464
rect 1841 840 1907 852
rect 1841 464 1857 840
rect 1891 464 1907 840
rect 1841 452 1907 464
rect 1937 840 2003 852
rect 1937 464 1953 840
rect 1987 464 2003 840
rect 1937 452 2003 464
rect 2033 840 2099 852
rect 2033 464 2049 840
rect 2083 464 2099 840
rect 2033 452 2099 464
rect 2129 840 2195 852
rect 2129 464 2145 840
rect 2179 464 2195 840
rect 2129 452 2195 464
rect 2225 840 2291 852
rect 2225 464 2241 840
rect 2275 464 2291 840
rect 2225 452 2291 464
rect 2321 840 2387 852
rect 2321 464 2337 840
rect 2371 464 2387 840
rect 2321 452 2387 464
rect 2417 840 2483 852
rect 2417 464 2433 840
rect 2467 464 2483 840
rect 2417 452 2483 464
rect 2513 840 2579 852
rect 2513 464 2529 840
rect 2563 464 2579 840
rect 2513 452 2579 464
rect 2609 840 2675 852
rect 2609 464 2625 840
rect 2659 464 2675 840
rect 2609 452 2675 464
rect 2705 840 2771 852
rect 2705 464 2721 840
rect 2755 464 2771 840
rect 2705 452 2771 464
rect 2801 840 2867 852
rect 2801 464 2817 840
rect 2851 464 2867 840
rect 2801 452 2867 464
rect 2897 840 2963 852
rect 2897 464 2913 840
rect 2947 464 2963 840
rect 2897 452 2963 464
rect 2993 840 3059 852
rect 2993 464 3009 840
rect 3043 464 3059 840
rect 2993 452 3059 464
rect 3089 840 3155 852
rect 3089 464 3105 840
rect 3139 464 3155 840
rect 3089 452 3155 464
rect 3185 840 3251 852
rect 3185 464 3201 840
rect 3235 464 3251 840
rect 3185 452 3251 464
rect 3281 840 3347 852
rect 3281 464 3297 840
rect 3331 464 3347 840
rect 3281 452 3347 464
rect 3377 840 3443 852
rect 3377 464 3393 840
rect 3427 464 3443 840
rect 3377 452 3443 464
rect 3473 840 3539 852
rect 3473 464 3489 840
rect 3523 464 3539 840
rect 3473 452 3539 464
rect 3569 840 3635 852
rect 3569 464 3585 840
rect 3619 464 3635 840
rect 3569 452 3635 464
rect 3665 840 3731 852
rect 3665 464 3681 840
rect 3715 464 3731 840
rect 3665 452 3731 464
rect 3761 840 3827 852
rect 3761 464 3777 840
rect 3811 464 3827 840
rect 3761 452 3827 464
rect 3857 840 3923 852
rect 3857 464 3873 840
rect 3907 464 3923 840
rect 3857 452 3923 464
rect 3953 840 4019 852
rect 3953 464 3969 840
rect 4003 464 4019 840
rect 3953 452 4019 464
rect 4049 840 4115 852
rect 4049 464 4065 840
rect 4099 464 4115 840
rect 4049 452 4115 464
rect 4145 840 4211 852
rect 4145 464 4161 840
rect 4195 464 4211 840
rect 4145 452 4211 464
rect 4241 840 4307 852
rect 4241 464 4257 840
rect 4291 464 4307 840
rect 4241 452 4307 464
rect 4337 840 4403 852
rect 4337 464 4353 840
rect 4387 464 4403 840
rect 4337 452 4403 464
rect 4433 840 4499 852
rect 4433 464 4449 840
rect 4483 464 4499 840
rect 4433 452 4499 464
rect 4529 840 4595 852
rect 4529 464 4545 840
rect 4579 464 4595 840
rect 4529 452 4595 464
rect 4625 840 4691 852
rect 4625 464 4641 840
rect 4675 464 4691 840
rect 4625 452 4691 464
rect 4721 840 4787 852
rect 4721 464 4737 840
rect 4771 464 4787 840
rect 4721 452 4787 464
rect 4817 840 4883 852
rect 4817 464 4833 840
rect 4867 464 4883 840
rect 4817 452 4883 464
rect 4913 840 4979 852
rect 4913 464 4929 840
rect 4963 464 4979 840
rect 4913 452 4979 464
rect 5009 840 5075 852
rect 5009 464 5025 840
rect 5059 464 5075 840
rect 5009 452 5075 464
rect 5105 840 5171 852
rect 5105 464 5121 840
rect 5155 464 5171 840
rect 5105 452 5171 464
rect 5201 840 5267 852
rect 5201 464 5217 840
rect 5251 464 5267 840
rect 5201 452 5267 464
rect 5297 840 5363 852
rect 5297 464 5313 840
rect 5347 464 5363 840
rect 5297 452 5363 464
rect 5393 840 5459 852
rect 5393 464 5409 840
rect 5443 464 5459 840
rect 5393 452 5459 464
rect 5489 840 5555 852
rect 5489 464 5505 840
rect 5539 464 5555 840
rect 5489 452 5555 464
rect 5585 840 5651 852
rect 5585 464 5601 840
rect 5635 464 5651 840
rect 5585 452 5651 464
rect 5681 840 5747 852
rect 5681 464 5697 840
rect 5731 464 5747 840
rect 5681 452 5747 464
rect 5777 840 5843 852
rect 5777 464 5793 840
rect 5827 464 5843 840
rect 5777 452 5843 464
rect 5873 840 5939 852
rect 5873 464 5889 840
rect 5923 464 5939 840
rect 5873 452 5939 464
rect 5969 840 6031 852
rect 5969 464 5985 840
rect 6019 464 6031 840
rect 5969 452 6031 464
rect 21 -1884 83 -1872
rect 21 -2260 33 -1884
rect 67 -2260 83 -1884
rect 21 -2272 83 -2260
rect 113 -1884 179 -1872
rect 113 -2260 129 -1884
rect 163 -2260 179 -1884
rect 113 -2272 179 -2260
rect 209 -1884 275 -1872
rect 209 -2260 225 -1884
rect 259 -2260 275 -1884
rect 209 -2272 275 -2260
rect 305 -1884 371 -1872
rect 305 -2260 321 -1884
rect 355 -2260 371 -1884
rect 305 -2272 371 -2260
rect 401 -1884 467 -1872
rect 401 -2260 417 -1884
rect 451 -2260 467 -1884
rect 401 -2272 467 -2260
rect 497 -1884 563 -1872
rect 497 -2260 513 -1884
rect 547 -2260 563 -1884
rect 497 -2272 563 -2260
rect 593 -1884 659 -1872
rect 593 -2260 609 -1884
rect 643 -2260 659 -1884
rect 593 -2272 659 -2260
rect 689 -1884 755 -1872
rect 689 -2260 705 -1884
rect 739 -2260 755 -1884
rect 689 -2272 755 -2260
rect 785 -1884 851 -1872
rect 785 -2260 801 -1884
rect 835 -2260 851 -1884
rect 785 -2272 851 -2260
rect 881 -1884 947 -1872
rect 881 -2260 897 -1884
rect 931 -2260 947 -1884
rect 881 -2272 947 -2260
rect 977 -1884 1043 -1872
rect 977 -2260 993 -1884
rect 1027 -2260 1043 -1884
rect 977 -2272 1043 -2260
rect 1073 -1884 1139 -1872
rect 1073 -2260 1089 -1884
rect 1123 -2260 1139 -1884
rect 1073 -2272 1139 -2260
rect 1169 -1884 1235 -1872
rect 1169 -2260 1185 -1884
rect 1219 -2260 1235 -1884
rect 1169 -2272 1235 -2260
rect 1265 -1884 1331 -1872
rect 1265 -2260 1281 -1884
rect 1315 -2260 1331 -1884
rect 1265 -2272 1331 -2260
rect 1361 -1884 1427 -1872
rect 1361 -2260 1377 -1884
rect 1411 -2260 1427 -1884
rect 1361 -2272 1427 -2260
rect 1457 -1884 1523 -1872
rect 1457 -2260 1473 -1884
rect 1507 -2260 1523 -1884
rect 1457 -2272 1523 -2260
rect 1553 -1884 1619 -1872
rect 1553 -2260 1569 -1884
rect 1603 -2260 1619 -1884
rect 1553 -2272 1619 -2260
rect 1649 -1884 1715 -1872
rect 1649 -2260 1665 -1884
rect 1699 -2260 1715 -1884
rect 1649 -2272 1715 -2260
rect 1745 -1884 1811 -1872
rect 1745 -2260 1761 -1884
rect 1795 -2260 1811 -1884
rect 1745 -2272 1811 -2260
rect 1841 -1884 1907 -1872
rect 1841 -2260 1857 -1884
rect 1891 -2260 1907 -1884
rect 1841 -2272 1907 -2260
rect 1937 -1884 2003 -1872
rect 1937 -2260 1953 -1884
rect 1987 -2260 2003 -1884
rect 1937 -2272 2003 -2260
rect 2033 -1884 2099 -1872
rect 2033 -2260 2049 -1884
rect 2083 -2260 2099 -1884
rect 2033 -2272 2099 -2260
rect 2129 -1884 2195 -1872
rect 2129 -2260 2145 -1884
rect 2179 -2260 2195 -1884
rect 2129 -2272 2195 -2260
rect 2225 -1884 2291 -1872
rect 2225 -2260 2241 -1884
rect 2275 -2260 2291 -1884
rect 2225 -2272 2291 -2260
rect 2321 -1884 2387 -1872
rect 2321 -2260 2337 -1884
rect 2371 -2260 2387 -1884
rect 2321 -2272 2387 -2260
rect 2417 -1884 2483 -1872
rect 2417 -2260 2433 -1884
rect 2467 -2260 2483 -1884
rect 2417 -2272 2483 -2260
rect 2513 -1884 2579 -1872
rect 2513 -2260 2529 -1884
rect 2563 -2260 2579 -1884
rect 2513 -2272 2579 -2260
rect 2609 -1884 2675 -1872
rect 2609 -2260 2625 -1884
rect 2659 -2260 2675 -1884
rect 2609 -2272 2675 -2260
rect 2705 -1884 2771 -1872
rect 2705 -2260 2721 -1884
rect 2755 -2260 2771 -1884
rect 2705 -2272 2771 -2260
rect 2801 -1884 2867 -1872
rect 2801 -2260 2817 -1884
rect 2851 -2260 2867 -1884
rect 2801 -2272 2867 -2260
rect 2897 -1884 2963 -1872
rect 2897 -2260 2913 -1884
rect 2947 -2260 2963 -1884
rect 2897 -2272 2963 -2260
rect 2993 -1884 3059 -1872
rect 2993 -2260 3009 -1884
rect 3043 -2260 3059 -1884
rect 2993 -2272 3059 -2260
rect 3089 -1884 3155 -1872
rect 3089 -2260 3105 -1884
rect 3139 -2260 3155 -1884
rect 3089 -2272 3155 -2260
rect 3185 -1884 3251 -1872
rect 3185 -2260 3201 -1884
rect 3235 -2260 3251 -1884
rect 3185 -2272 3251 -2260
rect 3281 -1884 3347 -1872
rect 3281 -2260 3297 -1884
rect 3331 -2260 3347 -1884
rect 3281 -2272 3347 -2260
rect 3377 -1884 3443 -1872
rect 3377 -2260 3393 -1884
rect 3427 -2260 3443 -1884
rect 3377 -2272 3443 -2260
rect 3473 -1884 3539 -1872
rect 3473 -2260 3489 -1884
rect 3523 -2260 3539 -1884
rect 3473 -2272 3539 -2260
rect 3569 -1884 3635 -1872
rect 3569 -2260 3585 -1884
rect 3619 -2260 3635 -1884
rect 3569 -2272 3635 -2260
rect 3665 -1884 3731 -1872
rect 3665 -2260 3681 -1884
rect 3715 -2260 3731 -1884
rect 3665 -2272 3731 -2260
rect 3761 -1884 3827 -1872
rect 3761 -2260 3777 -1884
rect 3811 -2260 3827 -1884
rect 3761 -2272 3827 -2260
rect 3857 -1884 3923 -1872
rect 3857 -2260 3873 -1884
rect 3907 -2260 3923 -1884
rect 3857 -2272 3923 -2260
rect 3953 -1884 4019 -1872
rect 3953 -2260 3969 -1884
rect 4003 -2260 4019 -1884
rect 3953 -2272 4019 -2260
rect 4049 -1884 4115 -1872
rect 4049 -2260 4065 -1884
rect 4099 -2260 4115 -1884
rect 4049 -2272 4115 -2260
rect 4145 -1884 4211 -1872
rect 4145 -2260 4161 -1884
rect 4195 -2260 4211 -1884
rect 4145 -2272 4211 -2260
rect 4241 -1884 4307 -1872
rect 4241 -2260 4257 -1884
rect 4291 -2260 4307 -1884
rect 4241 -2272 4307 -2260
rect 4337 -1884 4403 -1872
rect 4337 -2260 4353 -1884
rect 4387 -2260 4403 -1884
rect 4337 -2272 4403 -2260
rect 4433 -1884 4499 -1872
rect 4433 -2260 4449 -1884
rect 4483 -2260 4499 -1884
rect 4433 -2272 4499 -2260
rect 4529 -1884 4595 -1872
rect 4529 -2260 4545 -1884
rect 4579 -2260 4595 -1884
rect 4529 -2272 4595 -2260
rect 4625 -1884 4691 -1872
rect 4625 -2260 4641 -1884
rect 4675 -2260 4691 -1884
rect 4625 -2272 4691 -2260
rect 4721 -1884 4787 -1872
rect 4721 -2260 4737 -1884
rect 4771 -2260 4787 -1884
rect 4721 -2272 4787 -2260
rect 4817 -1884 4883 -1872
rect 4817 -2260 4833 -1884
rect 4867 -2260 4883 -1884
rect 4817 -2272 4883 -2260
rect 4913 -1884 4979 -1872
rect 4913 -2260 4929 -1884
rect 4963 -2260 4979 -1884
rect 4913 -2272 4979 -2260
rect 5009 -1884 5075 -1872
rect 5009 -2260 5025 -1884
rect 5059 -2260 5075 -1884
rect 5009 -2272 5075 -2260
rect 5105 -1884 5171 -1872
rect 5105 -2260 5121 -1884
rect 5155 -2260 5171 -1884
rect 5105 -2272 5171 -2260
rect 5201 -1884 5267 -1872
rect 5201 -2260 5217 -1884
rect 5251 -2260 5267 -1884
rect 5201 -2272 5267 -2260
rect 5297 -1884 5363 -1872
rect 5297 -2260 5313 -1884
rect 5347 -2260 5363 -1884
rect 5297 -2272 5363 -2260
rect 5393 -1884 5459 -1872
rect 5393 -2260 5409 -1884
rect 5443 -2260 5459 -1884
rect 5393 -2272 5459 -2260
rect 5489 -1884 5555 -1872
rect 5489 -2260 5505 -1884
rect 5539 -2260 5555 -1884
rect 5489 -2272 5555 -2260
rect 5585 -1884 5651 -1872
rect 5585 -2260 5601 -1884
rect 5635 -2260 5651 -1884
rect 5585 -2272 5651 -2260
rect 5681 -1884 5747 -1872
rect 5681 -2260 5697 -1884
rect 5731 -2260 5747 -1884
rect 5681 -2272 5747 -2260
rect 5777 -1884 5843 -1872
rect 5777 -2260 5793 -1884
rect 5827 -2260 5843 -1884
rect 5777 -2272 5843 -2260
rect 5873 -1884 5939 -1872
rect 5873 -2260 5889 -1884
rect 5923 -2260 5939 -1884
rect 5873 -2272 5939 -2260
rect 5969 -1884 6031 -1872
rect 5969 -2260 5985 -1884
rect 6019 -2260 6031 -1884
rect 5969 -2272 6031 -2260
<< pdiff >>
rect 21 1915 83 1927
rect 21 1219 33 1915
rect 67 1219 83 1915
rect 21 1207 83 1219
rect 113 1915 179 1927
rect 113 1219 129 1915
rect 163 1219 179 1915
rect 113 1207 179 1219
rect 209 1915 275 1927
rect 209 1219 225 1915
rect 259 1219 275 1915
rect 209 1207 275 1219
rect 305 1915 371 1927
rect 305 1219 321 1915
rect 355 1219 371 1915
rect 305 1207 371 1219
rect 401 1915 467 1927
rect 401 1219 417 1915
rect 451 1219 467 1915
rect 401 1207 467 1219
rect 497 1915 563 1927
rect 497 1219 513 1915
rect 547 1219 563 1915
rect 497 1207 563 1219
rect 593 1915 659 1927
rect 593 1219 609 1915
rect 643 1219 659 1915
rect 593 1207 659 1219
rect 689 1915 755 1927
rect 689 1219 705 1915
rect 739 1219 755 1915
rect 689 1207 755 1219
rect 785 1915 851 1927
rect 785 1219 801 1915
rect 835 1219 851 1915
rect 785 1207 851 1219
rect 881 1915 947 1927
rect 881 1219 897 1915
rect 931 1219 947 1915
rect 881 1207 947 1219
rect 977 1915 1043 1927
rect 977 1219 993 1915
rect 1027 1219 1043 1915
rect 977 1207 1043 1219
rect 1073 1915 1139 1927
rect 1073 1219 1089 1915
rect 1123 1219 1139 1915
rect 1073 1207 1139 1219
rect 1169 1915 1235 1927
rect 1169 1219 1185 1915
rect 1219 1219 1235 1915
rect 1169 1207 1235 1219
rect 1265 1915 1331 1927
rect 1265 1219 1281 1915
rect 1315 1219 1331 1915
rect 1265 1207 1331 1219
rect 1361 1915 1427 1927
rect 1361 1219 1377 1915
rect 1411 1219 1427 1915
rect 1361 1207 1427 1219
rect 1457 1915 1523 1927
rect 1457 1219 1473 1915
rect 1507 1219 1523 1915
rect 1457 1207 1523 1219
rect 1553 1915 1619 1927
rect 1553 1219 1569 1915
rect 1603 1219 1619 1915
rect 1553 1207 1619 1219
rect 1649 1915 1715 1927
rect 1649 1219 1665 1915
rect 1699 1219 1715 1915
rect 1649 1207 1715 1219
rect 1745 1915 1811 1927
rect 1745 1219 1761 1915
rect 1795 1219 1811 1915
rect 1745 1207 1811 1219
rect 1841 1915 1907 1927
rect 1841 1219 1857 1915
rect 1891 1219 1907 1915
rect 1841 1207 1907 1219
rect 1937 1915 2003 1927
rect 1937 1219 1953 1915
rect 1987 1219 2003 1915
rect 1937 1207 2003 1219
rect 2033 1915 2099 1927
rect 2033 1219 2049 1915
rect 2083 1219 2099 1915
rect 2033 1207 2099 1219
rect 2129 1915 2195 1927
rect 2129 1219 2145 1915
rect 2179 1219 2195 1915
rect 2129 1207 2195 1219
rect 2225 1915 2291 1927
rect 2225 1219 2241 1915
rect 2275 1219 2291 1915
rect 2225 1207 2291 1219
rect 2321 1915 2387 1927
rect 2321 1219 2337 1915
rect 2371 1219 2387 1915
rect 2321 1207 2387 1219
rect 2417 1915 2483 1927
rect 2417 1219 2433 1915
rect 2467 1219 2483 1915
rect 2417 1207 2483 1219
rect 2513 1915 2579 1927
rect 2513 1219 2529 1915
rect 2563 1219 2579 1915
rect 2513 1207 2579 1219
rect 2609 1915 2675 1927
rect 2609 1219 2625 1915
rect 2659 1219 2675 1915
rect 2609 1207 2675 1219
rect 2705 1915 2771 1927
rect 2705 1219 2721 1915
rect 2755 1219 2771 1915
rect 2705 1207 2771 1219
rect 2801 1915 2867 1927
rect 2801 1219 2817 1915
rect 2851 1219 2867 1915
rect 2801 1207 2867 1219
rect 2897 1915 2963 1927
rect 2897 1219 2913 1915
rect 2947 1219 2963 1915
rect 2897 1207 2963 1219
rect 2993 1915 3059 1927
rect 2993 1219 3009 1915
rect 3043 1219 3059 1915
rect 2993 1207 3059 1219
rect 3089 1915 3155 1927
rect 3089 1219 3105 1915
rect 3139 1219 3155 1915
rect 3089 1207 3155 1219
rect 3185 1915 3251 1927
rect 3185 1219 3201 1915
rect 3235 1219 3251 1915
rect 3185 1207 3251 1219
rect 3281 1915 3347 1927
rect 3281 1219 3297 1915
rect 3331 1219 3347 1915
rect 3281 1207 3347 1219
rect 3377 1915 3443 1927
rect 3377 1219 3393 1915
rect 3427 1219 3443 1915
rect 3377 1207 3443 1219
rect 3473 1915 3539 1927
rect 3473 1219 3489 1915
rect 3523 1219 3539 1915
rect 3473 1207 3539 1219
rect 3569 1915 3635 1927
rect 3569 1219 3585 1915
rect 3619 1219 3635 1915
rect 3569 1207 3635 1219
rect 3665 1915 3731 1927
rect 3665 1219 3681 1915
rect 3715 1219 3731 1915
rect 3665 1207 3731 1219
rect 3761 1915 3827 1927
rect 3761 1219 3777 1915
rect 3811 1219 3827 1915
rect 3761 1207 3827 1219
rect 3857 1915 3923 1927
rect 3857 1219 3873 1915
rect 3907 1219 3923 1915
rect 3857 1207 3923 1219
rect 3953 1915 4019 1927
rect 3953 1219 3969 1915
rect 4003 1219 4019 1915
rect 3953 1207 4019 1219
rect 4049 1915 4115 1927
rect 4049 1219 4065 1915
rect 4099 1219 4115 1915
rect 4049 1207 4115 1219
rect 4145 1915 4211 1927
rect 4145 1219 4161 1915
rect 4195 1219 4211 1915
rect 4145 1207 4211 1219
rect 4241 1915 4307 1927
rect 4241 1219 4257 1915
rect 4291 1219 4307 1915
rect 4241 1207 4307 1219
rect 4337 1915 4403 1927
rect 4337 1219 4353 1915
rect 4387 1219 4403 1915
rect 4337 1207 4403 1219
rect 4433 1915 4499 1927
rect 4433 1219 4449 1915
rect 4483 1219 4499 1915
rect 4433 1207 4499 1219
rect 4529 1915 4595 1927
rect 4529 1219 4545 1915
rect 4579 1219 4595 1915
rect 4529 1207 4595 1219
rect 4625 1915 4691 1927
rect 4625 1219 4641 1915
rect 4675 1219 4691 1915
rect 4625 1207 4691 1219
rect 4721 1915 4787 1927
rect 4721 1219 4737 1915
rect 4771 1219 4787 1915
rect 4721 1207 4787 1219
rect 4817 1915 4883 1927
rect 4817 1219 4833 1915
rect 4867 1219 4883 1915
rect 4817 1207 4883 1219
rect 4913 1915 4979 1927
rect 4913 1219 4929 1915
rect 4963 1219 4979 1915
rect 4913 1207 4979 1219
rect 5009 1915 5075 1927
rect 5009 1219 5025 1915
rect 5059 1219 5075 1915
rect 5009 1207 5075 1219
rect 5105 1915 5171 1927
rect 5105 1219 5121 1915
rect 5155 1219 5171 1915
rect 5105 1207 5171 1219
rect 5201 1915 5267 1927
rect 5201 1219 5217 1915
rect 5251 1219 5267 1915
rect 5201 1207 5267 1219
rect 5297 1915 5363 1927
rect 5297 1219 5313 1915
rect 5347 1219 5363 1915
rect 5297 1207 5363 1219
rect 5393 1915 5459 1927
rect 5393 1219 5409 1915
rect 5443 1219 5459 1915
rect 5393 1207 5459 1219
rect 5489 1915 5555 1927
rect 5489 1219 5505 1915
rect 5539 1219 5555 1915
rect 5489 1207 5555 1219
rect 5585 1915 5651 1927
rect 5585 1219 5601 1915
rect 5635 1219 5651 1915
rect 5585 1207 5651 1219
rect 5681 1915 5747 1927
rect 5681 1219 5697 1915
rect 5731 1219 5747 1915
rect 5681 1207 5747 1219
rect 5777 1915 5843 1927
rect 5777 1219 5793 1915
rect 5827 1219 5843 1915
rect 5777 1207 5843 1219
rect 5873 1915 5939 1927
rect 5873 1219 5889 1915
rect 5923 1219 5939 1915
rect 5873 1207 5939 1219
rect 5969 1915 6031 1927
rect 5969 1219 5985 1915
rect 6019 1219 6031 1915
rect 5969 1207 6031 1219
rect 21 -2639 83 -2627
rect 21 -3335 33 -2639
rect 67 -3335 83 -2639
rect 21 -3347 83 -3335
rect 113 -2639 179 -2627
rect 113 -3335 129 -2639
rect 163 -3335 179 -2639
rect 113 -3347 179 -3335
rect 209 -2639 275 -2627
rect 209 -3335 225 -2639
rect 259 -3335 275 -2639
rect 209 -3347 275 -3335
rect 305 -2639 371 -2627
rect 305 -3335 321 -2639
rect 355 -3335 371 -2639
rect 305 -3347 371 -3335
rect 401 -2639 467 -2627
rect 401 -3335 417 -2639
rect 451 -3335 467 -2639
rect 401 -3347 467 -3335
rect 497 -2639 563 -2627
rect 497 -3335 513 -2639
rect 547 -3335 563 -2639
rect 497 -3347 563 -3335
rect 593 -2639 659 -2627
rect 593 -3335 609 -2639
rect 643 -3335 659 -2639
rect 593 -3347 659 -3335
rect 689 -2639 755 -2627
rect 689 -3335 705 -2639
rect 739 -3335 755 -2639
rect 689 -3347 755 -3335
rect 785 -2639 851 -2627
rect 785 -3335 801 -2639
rect 835 -3335 851 -2639
rect 785 -3347 851 -3335
rect 881 -2639 947 -2627
rect 881 -3335 897 -2639
rect 931 -3335 947 -2639
rect 881 -3347 947 -3335
rect 977 -2639 1043 -2627
rect 977 -3335 993 -2639
rect 1027 -3335 1043 -2639
rect 977 -3347 1043 -3335
rect 1073 -2639 1139 -2627
rect 1073 -3335 1089 -2639
rect 1123 -3335 1139 -2639
rect 1073 -3347 1139 -3335
rect 1169 -2639 1235 -2627
rect 1169 -3335 1185 -2639
rect 1219 -3335 1235 -2639
rect 1169 -3347 1235 -3335
rect 1265 -2639 1331 -2627
rect 1265 -3335 1281 -2639
rect 1315 -3335 1331 -2639
rect 1265 -3347 1331 -3335
rect 1361 -2639 1427 -2627
rect 1361 -3335 1377 -2639
rect 1411 -3335 1427 -2639
rect 1361 -3347 1427 -3335
rect 1457 -2639 1523 -2627
rect 1457 -3335 1473 -2639
rect 1507 -3335 1523 -2639
rect 1457 -3347 1523 -3335
rect 1553 -2639 1619 -2627
rect 1553 -3335 1569 -2639
rect 1603 -3335 1619 -2639
rect 1553 -3347 1619 -3335
rect 1649 -2639 1715 -2627
rect 1649 -3335 1665 -2639
rect 1699 -3335 1715 -2639
rect 1649 -3347 1715 -3335
rect 1745 -2639 1811 -2627
rect 1745 -3335 1761 -2639
rect 1795 -3335 1811 -2639
rect 1745 -3347 1811 -3335
rect 1841 -2639 1907 -2627
rect 1841 -3335 1857 -2639
rect 1891 -3335 1907 -2639
rect 1841 -3347 1907 -3335
rect 1937 -2639 2003 -2627
rect 1937 -3335 1953 -2639
rect 1987 -3335 2003 -2639
rect 1937 -3347 2003 -3335
rect 2033 -2639 2099 -2627
rect 2033 -3335 2049 -2639
rect 2083 -3335 2099 -2639
rect 2033 -3347 2099 -3335
rect 2129 -2639 2195 -2627
rect 2129 -3335 2145 -2639
rect 2179 -3335 2195 -2639
rect 2129 -3347 2195 -3335
rect 2225 -2639 2291 -2627
rect 2225 -3335 2241 -2639
rect 2275 -3335 2291 -2639
rect 2225 -3347 2291 -3335
rect 2321 -2639 2387 -2627
rect 2321 -3335 2337 -2639
rect 2371 -3335 2387 -2639
rect 2321 -3347 2387 -3335
rect 2417 -2639 2483 -2627
rect 2417 -3335 2433 -2639
rect 2467 -3335 2483 -2639
rect 2417 -3347 2483 -3335
rect 2513 -2639 2579 -2627
rect 2513 -3335 2529 -2639
rect 2563 -3335 2579 -2639
rect 2513 -3347 2579 -3335
rect 2609 -2639 2675 -2627
rect 2609 -3335 2625 -2639
rect 2659 -3335 2675 -2639
rect 2609 -3347 2675 -3335
rect 2705 -2639 2771 -2627
rect 2705 -3335 2721 -2639
rect 2755 -3335 2771 -2639
rect 2705 -3347 2771 -3335
rect 2801 -2639 2867 -2627
rect 2801 -3335 2817 -2639
rect 2851 -3335 2867 -2639
rect 2801 -3347 2867 -3335
rect 2897 -2639 2963 -2627
rect 2897 -3335 2913 -2639
rect 2947 -3335 2963 -2639
rect 2897 -3347 2963 -3335
rect 2993 -2639 3059 -2627
rect 2993 -3335 3009 -2639
rect 3043 -3335 3059 -2639
rect 2993 -3347 3059 -3335
rect 3089 -2639 3155 -2627
rect 3089 -3335 3105 -2639
rect 3139 -3335 3155 -2639
rect 3089 -3347 3155 -3335
rect 3185 -2639 3251 -2627
rect 3185 -3335 3201 -2639
rect 3235 -3335 3251 -2639
rect 3185 -3347 3251 -3335
rect 3281 -2639 3347 -2627
rect 3281 -3335 3297 -2639
rect 3331 -3335 3347 -2639
rect 3281 -3347 3347 -3335
rect 3377 -2639 3443 -2627
rect 3377 -3335 3393 -2639
rect 3427 -3335 3443 -2639
rect 3377 -3347 3443 -3335
rect 3473 -2639 3539 -2627
rect 3473 -3335 3489 -2639
rect 3523 -3335 3539 -2639
rect 3473 -3347 3539 -3335
rect 3569 -2639 3635 -2627
rect 3569 -3335 3585 -2639
rect 3619 -3335 3635 -2639
rect 3569 -3347 3635 -3335
rect 3665 -2639 3731 -2627
rect 3665 -3335 3681 -2639
rect 3715 -3335 3731 -2639
rect 3665 -3347 3731 -3335
rect 3761 -2639 3827 -2627
rect 3761 -3335 3777 -2639
rect 3811 -3335 3827 -2639
rect 3761 -3347 3827 -3335
rect 3857 -2639 3923 -2627
rect 3857 -3335 3873 -2639
rect 3907 -3335 3923 -2639
rect 3857 -3347 3923 -3335
rect 3953 -2639 4019 -2627
rect 3953 -3335 3969 -2639
rect 4003 -3335 4019 -2639
rect 3953 -3347 4019 -3335
rect 4049 -2639 4115 -2627
rect 4049 -3335 4065 -2639
rect 4099 -3335 4115 -2639
rect 4049 -3347 4115 -3335
rect 4145 -2639 4211 -2627
rect 4145 -3335 4161 -2639
rect 4195 -3335 4211 -2639
rect 4145 -3347 4211 -3335
rect 4241 -2639 4307 -2627
rect 4241 -3335 4257 -2639
rect 4291 -3335 4307 -2639
rect 4241 -3347 4307 -3335
rect 4337 -2639 4403 -2627
rect 4337 -3335 4353 -2639
rect 4387 -3335 4403 -2639
rect 4337 -3347 4403 -3335
rect 4433 -2639 4499 -2627
rect 4433 -3335 4449 -2639
rect 4483 -3335 4499 -2639
rect 4433 -3347 4499 -3335
rect 4529 -2639 4595 -2627
rect 4529 -3335 4545 -2639
rect 4579 -3335 4595 -2639
rect 4529 -3347 4595 -3335
rect 4625 -2639 4691 -2627
rect 4625 -3335 4641 -2639
rect 4675 -3335 4691 -2639
rect 4625 -3347 4691 -3335
rect 4721 -2639 4787 -2627
rect 4721 -3335 4737 -2639
rect 4771 -3335 4787 -2639
rect 4721 -3347 4787 -3335
rect 4817 -2639 4883 -2627
rect 4817 -3335 4833 -2639
rect 4867 -3335 4883 -2639
rect 4817 -3347 4883 -3335
rect 4913 -2639 4979 -2627
rect 4913 -3335 4929 -2639
rect 4963 -3335 4979 -2639
rect 4913 -3347 4979 -3335
rect 5009 -2639 5075 -2627
rect 5009 -3335 5025 -2639
rect 5059 -3335 5075 -2639
rect 5009 -3347 5075 -3335
rect 5105 -2639 5171 -2627
rect 5105 -3335 5121 -2639
rect 5155 -3335 5171 -2639
rect 5105 -3347 5171 -3335
rect 5201 -2639 5267 -2627
rect 5201 -3335 5217 -2639
rect 5251 -3335 5267 -2639
rect 5201 -3347 5267 -3335
rect 5297 -2639 5363 -2627
rect 5297 -3335 5313 -2639
rect 5347 -3335 5363 -2639
rect 5297 -3347 5363 -3335
rect 5393 -2639 5459 -2627
rect 5393 -3335 5409 -2639
rect 5443 -3335 5459 -2639
rect 5393 -3347 5459 -3335
rect 5489 -2639 5555 -2627
rect 5489 -3335 5505 -2639
rect 5539 -3335 5555 -2639
rect 5489 -3347 5555 -3335
rect 5585 -2639 5651 -2627
rect 5585 -3335 5601 -2639
rect 5635 -3335 5651 -2639
rect 5585 -3347 5651 -3335
rect 5681 -2639 5747 -2627
rect 5681 -3335 5697 -2639
rect 5731 -3335 5747 -2639
rect 5681 -3347 5747 -3335
rect 5777 -2639 5843 -2627
rect 5777 -3335 5793 -2639
rect 5827 -3335 5843 -2639
rect 5777 -3347 5843 -3335
rect 5873 -2639 5939 -2627
rect 5873 -3335 5889 -2639
rect 5923 -3335 5939 -2639
rect 5873 -3347 5939 -3335
rect 5969 -2639 6031 -2627
rect 5969 -3335 5985 -2639
rect 6019 -3335 6031 -2639
rect 5969 -3347 6031 -3335
<< ndiffc >>
rect 33 464 67 840
rect 129 464 163 840
rect 225 464 259 840
rect 321 464 355 840
rect 417 464 451 840
rect 513 464 547 840
rect 609 464 643 840
rect 705 464 739 840
rect 801 464 835 840
rect 897 464 931 840
rect 993 464 1027 840
rect 1089 464 1123 840
rect 1185 464 1219 840
rect 1281 464 1315 840
rect 1377 464 1411 840
rect 1473 464 1507 840
rect 1569 464 1603 840
rect 1665 464 1699 840
rect 1761 464 1795 840
rect 1857 464 1891 840
rect 1953 464 1987 840
rect 2049 464 2083 840
rect 2145 464 2179 840
rect 2241 464 2275 840
rect 2337 464 2371 840
rect 2433 464 2467 840
rect 2529 464 2563 840
rect 2625 464 2659 840
rect 2721 464 2755 840
rect 2817 464 2851 840
rect 2913 464 2947 840
rect 3009 464 3043 840
rect 3105 464 3139 840
rect 3201 464 3235 840
rect 3297 464 3331 840
rect 3393 464 3427 840
rect 3489 464 3523 840
rect 3585 464 3619 840
rect 3681 464 3715 840
rect 3777 464 3811 840
rect 3873 464 3907 840
rect 3969 464 4003 840
rect 4065 464 4099 840
rect 4161 464 4195 840
rect 4257 464 4291 840
rect 4353 464 4387 840
rect 4449 464 4483 840
rect 4545 464 4579 840
rect 4641 464 4675 840
rect 4737 464 4771 840
rect 4833 464 4867 840
rect 4929 464 4963 840
rect 5025 464 5059 840
rect 5121 464 5155 840
rect 5217 464 5251 840
rect 5313 464 5347 840
rect 5409 464 5443 840
rect 5505 464 5539 840
rect 5601 464 5635 840
rect 5697 464 5731 840
rect 5793 464 5827 840
rect 5889 464 5923 840
rect 5985 464 6019 840
rect 33 -2260 67 -1884
rect 129 -2260 163 -1884
rect 225 -2260 259 -1884
rect 321 -2260 355 -1884
rect 417 -2260 451 -1884
rect 513 -2260 547 -1884
rect 609 -2260 643 -1884
rect 705 -2260 739 -1884
rect 801 -2260 835 -1884
rect 897 -2260 931 -1884
rect 993 -2260 1027 -1884
rect 1089 -2260 1123 -1884
rect 1185 -2260 1219 -1884
rect 1281 -2260 1315 -1884
rect 1377 -2260 1411 -1884
rect 1473 -2260 1507 -1884
rect 1569 -2260 1603 -1884
rect 1665 -2260 1699 -1884
rect 1761 -2260 1795 -1884
rect 1857 -2260 1891 -1884
rect 1953 -2260 1987 -1884
rect 2049 -2260 2083 -1884
rect 2145 -2260 2179 -1884
rect 2241 -2260 2275 -1884
rect 2337 -2260 2371 -1884
rect 2433 -2260 2467 -1884
rect 2529 -2260 2563 -1884
rect 2625 -2260 2659 -1884
rect 2721 -2260 2755 -1884
rect 2817 -2260 2851 -1884
rect 2913 -2260 2947 -1884
rect 3009 -2260 3043 -1884
rect 3105 -2260 3139 -1884
rect 3201 -2260 3235 -1884
rect 3297 -2260 3331 -1884
rect 3393 -2260 3427 -1884
rect 3489 -2260 3523 -1884
rect 3585 -2260 3619 -1884
rect 3681 -2260 3715 -1884
rect 3777 -2260 3811 -1884
rect 3873 -2260 3907 -1884
rect 3969 -2260 4003 -1884
rect 4065 -2260 4099 -1884
rect 4161 -2260 4195 -1884
rect 4257 -2260 4291 -1884
rect 4353 -2260 4387 -1884
rect 4449 -2260 4483 -1884
rect 4545 -2260 4579 -1884
rect 4641 -2260 4675 -1884
rect 4737 -2260 4771 -1884
rect 4833 -2260 4867 -1884
rect 4929 -2260 4963 -1884
rect 5025 -2260 5059 -1884
rect 5121 -2260 5155 -1884
rect 5217 -2260 5251 -1884
rect 5313 -2260 5347 -1884
rect 5409 -2260 5443 -1884
rect 5505 -2260 5539 -1884
rect 5601 -2260 5635 -1884
rect 5697 -2260 5731 -1884
rect 5793 -2260 5827 -1884
rect 5889 -2260 5923 -1884
rect 5985 -2260 6019 -1884
<< pdiffc >>
rect 33 1219 67 1915
rect 129 1219 163 1915
rect 225 1219 259 1915
rect 321 1219 355 1915
rect 417 1219 451 1915
rect 513 1219 547 1915
rect 609 1219 643 1915
rect 705 1219 739 1915
rect 801 1219 835 1915
rect 897 1219 931 1915
rect 993 1219 1027 1915
rect 1089 1219 1123 1915
rect 1185 1219 1219 1915
rect 1281 1219 1315 1915
rect 1377 1219 1411 1915
rect 1473 1219 1507 1915
rect 1569 1219 1603 1915
rect 1665 1219 1699 1915
rect 1761 1219 1795 1915
rect 1857 1219 1891 1915
rect 1953 1219 1987 1915
rect 2049 1219 2083 1915
rect 2145 1219 2179 1915
rect 2241 1219 2275 1915
rect 2337 1219 2371 1915
rect 2433 1219 2467 1915
rect 2529 1219 2563 1915
rect 2625 1219 2659 1915
rect 2721 1219 2755 1915
rect 2817 1219 2851 1915
rect 2913 1219 2947 1915
rect 3009 1219 3043 1915
rect 3105 1219 3139 1915
rect 3201 1219 3235 1915
rect 3297 1219 3331 1915
rect 3393 1219 3427 1915
rect 3489 1219 3523 1915
rect 3585 1219 3619 1915
rect 3681 1219 3715 1915
rect 3777 1219 3811 1915
rect 3873 1219 3907 1915
rect 3969 1219 4003 1915
rect 4065 1219 4099 1915
rect 4161 1219 4195 1915
rect 4257 1219 4291 1915
rect 4353 1219 4387 1915
rect 4449 1219 4483 1915
rect 4545 1219 4579 1915
rect 4641 1219 4675 1915
rect 4737 1219 4771 1915
rect 4833 1219 4867 1915
rect 4929 1219 4963 1915
rect 5025 1219 5059 1915
rect 5121 1219 5155 1915
rect 5217 1219 5251 1915
rect 5313 1219 5347 1915
rect 5409 1219 5443 1915
rect 5505 1219 5539 1915
rect 5601 1219 5635 1915
rect 5697 1219 5731 1915
rect 5793 1219 5827 1915
rect 5889 1219 5923 1915
rect 5985 1219 6019 1915
rect 33 -3335 67 -2639
rect 129 -3335 163 -2639
rect 225 -3335 259 -2639
rect 321 -3335 355 -2639
rect 417 -3335 451 -2639
rect 513 -3335 547 -2639
rect 609 -3335 643 -2639
rect 705 -3335 739 -2639
rect 801 -3335 835 -2639
rect 897 -3335 931 -2639
rect 993 -3335 1027 -2639
rect 1089 -3335 1123 -2639
rect 1185 -3335 1219 -2639
rect 1281 -3335 1315 -2639
rect 1377 -3335 1411 -2639
rect 1473 -3335 1507 -2639
rect 1569 -3335 1603 -2639
rect 1665 -3335 1699 -2639
rect 1761 -3335 1795 -2639
rect 1857 -3335 1891 -2639
rect 1953 -3335 1987 -2639
rect 2049 -3335 2083 -2639
rect 2145 -3335 2179 -2639
rect 2241 -3335 2275 -2639
rect 2337 -3335 2371 -2639
rect 2433 -3335 2467 -2639
rect 2529 -3335 2563 -2639
rect 2625 -3335 2659 -2639
rect 2721 -3335 2755 -2639
rect 2817 -3335 2851 -2639
rect 2913 -3335 2947 -2639
rect 3009 -3335 3043 -2639
rect 3105 -3335 3139 -2639
rect 3201 -3335 3235 -2639
rect 3297 -3335 3331 -2639
rect 3393 -3335 3427 -2639
rect 3489 -3335 3523 -2639
rect 3585 -3335 3619 -2639
rect 3681 -3335 3715 -2639
rect 3777 -3335 3811 -2639
rect 3873 -3335 3907 -2639
rect 3969 -3335 4003 -2639
rect 4065 -3335 4099 -2639
rect 4161 -3335 4195 -2639
rect 4257 -3335 4291 -2639
rect 4353 -3335 4387 -2639
rect 4449 -3335 4483 -2639
rect 4545 -3335 4579 -2639
rect 4641 -3335 4675 -2639
rect 4737 -3335 4771 -2639
rect 4833 -3335 4867 -2639
rect 4929 -3335 4963 -2639
rect 5025 -3335 5059 -2639
rect 5121 -3335 5155 -2639
rect 5217 -3335 5251 -2639
rect 5313 -3335 5347 -2639
rect 5409 -3335 5443 -2639
rect 5505 -3335 5539 -2639
rect 5601 -3335 5635 -2639
rect 5697 -3335 5731 -2639
rect 5793 -3335 5827 -2639
rect 5889 -3335 5923 -2639
rect 5985 -3335 6019 -2639
<< psubdiff >>
rect 26 322 126 356
rect 5926 322 6026 356
rect 26 -1776 126 -1742
rect 5926 -1776 6026 -1742
<< nsubdiff >>
rect 26 2024 126 2058
rect 5926 2024 6026 2058
rect 26 -3478 126 -3444
rect 5926 -3478 6026 -3444
<< psubdiffcont >>
rect 126 322 5926 356
rect 126 -1776 5926 -1742
<< nsubdiffcont >>
rect 126 2024 5926 2058
rect 126 -3478 5926 -3444
<< poly >>
rect 83 1927 113 1958
rect 179 1927 209 1958
rect 275 1927 305 1958
rect 371 1927 401 1958
rect 467 1927 497 1958
rect 563 1927 593 1958
rect 659 1927 689 1958
rect 755 1927 785 1958
rect 851 1927 881 1958
rect 947 1927 977 1958
rect 1043 1927 1073 1958
rect 1139 1927 1169 1958
rect 1235 1927 1265 1958
rect 1331 1927 1361 1958
rect 1427 1927 1457 1958
rect 1523 1927 1553 1958
rect 1619 1927 1649 1958
rect 1715 1927 1745 1958
rect 1811 1927 1841 1958
rect 1907 1927 1937 1958
rect 2003 1927 2033 1958
rect 2099 1927 2129 1958
rect 2195 1927 2225 1958
rect 2291 1927 2321 1958
rect 2387 1927 2417 1958
rect 2483 1927 2513 1958
rect 2579 1927 2609 1958
rect 2675 1927 2705 1958
rect 2771 1927 2801 1958
rect 2867 1927 2897 1958
rect 2963 1927 2993 1958
rect 3059 1927 3089 1958
rect 3155 1927 3185 1958
rect 3251 1927 3281 1958
rect 3347 1927 3377 1958
rect 3443 1927 3473 1958
rect 3539 1927 3569 1958
rect 3635 1927 3665 1958
rect 3731 1927 3761 1958
rect 3827 1927 3857 1958
rect 3923 1927 3953 1958
rect 4019 1927 4049 1958
rect 4115 1927 4145 1958
rect 4211 1927 4241 1958
rect 4307 1927 4337 1958
rect 4403 1927 4433 1958
rect 4499 1927 4529 1958
rect 4595 1927 4625 1958
rect 4691 1927 4721 1958
rect 4787 1927 4817 1958
rect 4883 1927 4913 1958
rect 4979 1927 5009 1958
rect 5075 1927 5105 1958
rect 5171 1927 5201 1958
rect 5267 1927 5297 1958
rect 5363 1927 5393 1958
rect 5459 1927 5489 1958
rect 5555 1927 5585 1958
rect 5651 1927 5681 1958
rect 5747 1927 5777 1958
rect 5843 1927 5873 1958
rect 5939 1927 5969 1958
rect 83 1176 113 1207
rect 179 1176 209 1207
rect 83 1160 209 1176
rect 83 1126 93 1160
rect 198 1126 209 1160
rect 83 1110 209 1126
rect 275 1176 305 1207
rect 371 1176 401 1207
rect 275 1160 401 1176
rect 275 1126 285 1160
rect 390 1126 401 1160
rect 275 1110 401 1126
rect 467 1176 497 1207
rect 563 1176 593 1207
rect 467 1160 593 1176
rect 467 1126 477 1160
rect 582 1126 593 1160
rect 467 1110 593 1126
rect 659 1176 689 1207
rect 755 1176 785 1207
rect 659 1160 785 1176
rect 659 1126 669 1160
rect 774 1126 785 1160
rect 659 1110 785 1126
rect 851 1176 881 1207
rect 947 1176 977 1207
rect 851 1160 977 1176
rect 851 1126 861 1160
rect 966 1126 977 1160
rect 851 1110 977 1126
rect 1043 1176 1073 1207
rect 1139 1176 1169 1207
rect 1043 1160 1169 1176
rect 1043 1126 1053 1160
rect 1158 1126 1169 1160
rect 1043 1110 1169 1126
rect 1235 1176 1265 1207
rect 1331 1176 1361 1207
rect 1235 1160 1361 1176
rect 1235 1126 1245 1160
rect 1350 1126 1361 1160
rect 1235 1110 1361 1126
rect 1427 1176 1457 1207
rect 1523 1176 1553 1207
rect 1427 1160 1553 1176
rect 1427 1126 1437 1160
rect 1542 1126 1553 1160
rect 1427 1110 1553 1126
rect 1619 1176 1649 1207
rect 1715 1176 1745 1207
rect 1619 1160 1745 1176
rect 1619 1126 1630 1160
rect 1735 1126 1745 1160
rect 1619 1110 1745 1126
rect 1811 1176 1841 1207
rect 1907 1176 1937 1207
rect 1811 1160 1937 1176
rect 1811 1126 1822 1160
rect 1927 1126 1937 1160
rect 1811 1110 1937 1126
rect 2003 1176 2033 1207
rect 2099 1176 2129 1207
rect 2003 1160 2129 1176
rect 2003 1126 2014 1160
rect 2119 1126 2129 1160
rect 2003 1110 2129 1126
rect 2195 1176 2225 1207
rect 2291 1176 2321 1207
rect 2195 1160 2321 1176
rect 2195 1126 2206 1160
rect 2311 1126 2321 1160
rect 2195 1110 2321 1126
rect 2387 1176 2417 1207
rect 2483 1176 2513 1207
rect 2387 1160 2513 1176
rect 2387 1126 2398 1160
rect 2503 1126 2513 1160
rect 2387 1110 2513 1126
rect 2579 1176 2609 1207
rect 2675 1176 2705 1207
rect 2579 1160 2705 1176
rect 2579 1126 2590 1160
rect 2695 1126 2705 1160
rect 2579 1110 2705 1126
rect 2771 1176 2801 1207
rect 2867 1176 2897 1207
rect 2771 1160 2897 1176
rect 2771 1126 2782 1160
rect 2887 1126 2897 1160
rect 2771 1110 2897 1126
rect 2963 1176 2993 1207
rect 3059 1176 3089 1207
rect 2963 1160 3089 1176
rect 2963 1126 2973 1160
rect 3079 1126 3089 1160
rect 2963 1110 3089 1126
rect 3155 1176 3185 1207
rect 3251 1176 3281 1207
rect 3155 1160 3281 1176
rect 3155 1126 3165 1160
rect 3270 1126 3281 1160
rect 3155 1110 3281 1126
rect 3347 1176 3377 1207
rect 3443 1176 3473 1207
rect 3347 1160 3473 1176
rect 3347 1126 3357 1160
rect 3462 1126 3473 1160
rect 3347 1110 3473 1126
rect 3539 1176 3569 1207
rect 3635 1176 3665 1207
rect 3539 1160 3665 1176
rect 3539 1126 3549 1160
rect 3654 1126 3665 1160
rect 3539 1110 3665 1126
rect 3731 1176 3761 1207
rect 3827 1176 3857 1207
rect 3731 1160 3857 1176
rect 3731 1126 3741 1160
rect 3846 1126 3857 1160
rect 3731 1110 3857 1126
rect 3923 1176 3953 1207
rect 4019 1176 4049 1207
rect 3923 1160 4049 1176
rect 3923 1126 3933 1160
rect 4038 1126 4049 1160
rect 3923 1110 4049 1126
rect 4115 1176 4145 1207
rect 4211 1176 4241 1207
rect 4115 1160 4241 1176
rect 4115 1126 4125 1160
rect 4230 1126 4241 1160
rect 4115 1110 4241 1126
rect 4307 1176 4337 1207
rect 4403 1176 4433 1207
rect 4307 1160 4433 1176
rect 4307 1126 4317 1160
rect 4422 1126 4433 1160
rect 4307 1110 4433 1126
rect 4499 1176 4529 1207
rect 4595 1176 4625 1207
rect 4499 1160 4625 1176
rect 4499 1126 4510 1160
rect 4615 1126 4625 1160
rect 4499 1110 4625 1126
rect 4691 1176 4721 1207
rect 4787 1176 4817 1207
rect 4691 1160 4817 1176
rect 4691 1126 4702 1160
rect 4807 1126 4817 1160
rect 4691 1110 4817 1126
rect 4883 1176 4913 1207
rect 4979 1176 5009 1207
rect 4883 1160 5009 1176
rect 4883 1126 4894 1160
rect 4999 1126 5009 1160
rect 4883 1110 5009 1126
rect 5075 1176 5105 1207
rect 5171 1176 5201 1207
rect 5075 1160 5201 1176
rect 5075 1126 5086 1160
rect 5191 1126 5201 1160
rect 5075 1110 5201 1126
rect 5267 1176 5297 1207
rect 5363 1176 5393 1207
rect 5267 1160 5393 1176
rect 5267 1126 5278 1160
rect 5383 1126 5393 1160
rect 5267 1110 5393 1126
rect 5459 1176 5489 1207
rect 5555 1176 5585 1207
rect 5459 1160 5585 1176
rect 5459 1126 5470 1160
rect 5575 1126 5585 1160
rect 5459 1110 5585 1126
rect 5651 1176 5681 1207
rect 5747 1176 5777 1207
rect 5651 1160 5777 1176
rect 5651 1126 5662 1160
rect 5767 1126 5777 1160
rect 5651 1110 5777 1126
rect 5843 1176 5873 1207
rect 5939 1176 5969 1207
rect 5843 1160 5969 1176
rect 5843 1126 5854 1160
rect 5959 1126 5969 1160
rect 5843 1110 5969 1126
rect 83 924 305 940
rect 83 890 93 924
rect 198 890 305 924
rect 83 874 305 890
rect 350 930 422 940
rect 350 896 368 930
rect 402 896 422 930
rect 350 874 422 896
rect 467 924 593 940
rect 467 890 477 924
rect 582 890 593 924
rect 467 874 593 890
rect 83 852 113 874
rect 179 852 209 874
rect 275 852 305 874
rect 371 852 401 874
rect 467 852 497 874
rect 563 852 593 874
rect 659 924 785 940
rect 659 890 669 924
rect 774 890 785 924
rect 659 874 785 890
rect 659 852 689 874
rect 755 852 785 874
rect 851 924 977 940
rect 851 890 861 924
rect 966 890 977 924
rect 851 874 977 890
rect 851 852 881 874
rect 947 852 977 874
rect 1043 924 1169 940
rect 1043 890 1053 924
rect 1158 890 1169 924
rect 1043 874 1169 890
rect 1043 852 1073 874
rect 1139 852 1169 874
rect 1235 924 1361 940
rect 1235 890 1245 924
rect 1350 890 1361 924
rect 1235 874 1361 890
rect 1235 852 1265 874
rect 1331 852 1361 874
rect 1427 924 1553 940
rect 1427 890 1437 924
rect 1542 890 1553 924
rect 1427 874 1553 890
rect 1427 852 1457 874
rect 1523 852 1553 874
rect 1619 924 1745 940
rect 1619 890 1630 924
rect 1735 890 1745 924
rect 1619 874 1745 890
rect 1619 852 1649 874
rect 1715 852 1745 874
rect 1811 924 1937 940
rect 1811 890 1822 924
rect 1927 890 1937 924
rect 1811 874 1937 890
rect 1811 852 1841 874
rect 1907 852 1937 874
rect 2003 924 2129 940
rect 2003 890 2014 924
rect 2119 890 2129 924
rect 2003 874 2129 890
rect 2003 852 2033 874
rect 2099 852 2129 874
rect 2195 924 2321 940
rect 2195 890 2206 924
rect 2311 890 2321 924
rect 2195 874 2321 890
rect 2195 852 2225 874
rect 2291 852 2321 874
rect 2387 924 2513 940
rect 2387 890 2398 924
rect 2503 890 2513 924
rect 2387 874 2513 890
rect 2387 852 2417 874
rect 2483 852 2513 874
rect 2579 924 2705 940
rect 2579 890 2590 924
rect 2695 890 2705 924
rect 2579 874 2705 890
rect 2750 930 2822 940
rect 2750 896 2770 930
rect 2804 896 2822 930
rect 2750 874 2822 896
rect 2867 924 3185 940
rect 2867 890 2973 924
rect 3079 890 3185 924
rect 2867 874 3185 890
rect 3230 930 3302 940
rect 3230 896 3248 930
rect 3282 896 3302 930
rect 3230 874 3302 896
rect 3347 924 3473 940
rect 3347 890 3357 924
rect 3462 890 3473 924
rect 3347 874 3473 890
rect 2579 852 2609 874
rect 2675 852 2705 874
rect 2771 852 2801 874
rect 2867 852 2897 874
rect 2963 852 2993 874
rect 3059 852 3089 874
rect 3155 852 3185 874
rect 3251 852 3281 874
rect 3347 852 3377 874
rect 3443 852 3473 874
rect 3539 924 3665 940
rect 3539 890 3549 924
rect 3654 890 3665 924
rect 3539 874 3665 890
rect 3539 852 3569 874
rect 3635 852 3665 874
rect 3731 924 3857 940
rect 3731 890 3741 924
rect 3846 890 3857 924
rect 3731 874 3857 890
rect 3731 852 3761 874
rect 3827 852 3857 874
rect 3923 924 4049 940
rect 3923 890 3933 924
rect 4038 890 4049 924
rect 3923 874 4049 890
rect 3923 852 3953 874
rect 4019 852 4049 874
rect 4115 924 4241 940
rect 4115 890 4125 924
rect 4230 890 4241 924
rect 4115 874 4241 890
rect 4115 852 4145 874
rect 4211 852 4241 874
rect 4307 924 4433 940
rect 4307 890 4317 924
rect 4422 890 4433 924
rect 4307 874 4433 890
rect 4307 852 4337 874
rect 4403 852 4433 874
rect 4499 924 4625 940
rect 4499 890 4510 924
rect 4615 890 4625 924
rect 4499 874 4625 890
rect 4499 852 4529 874
rect 4595 852 4625 874
rect 4691 924 4817 940
rect 4691 890 4702 924
rect 4807 890 4817 924
rect 4691 874 4817 890
rect 4691 852 4721 874
rect 4787 852 4817 874
rect 4883 924 5009 940
rect 4883 890 4894 924
rect 4999 890 5009 924
rect 4883 874 5009 890
rect 4883 852 4913 874
rect 4979 852 5009 874
rect 5075 924 5201 940
rect 5075 890 5086 924
rect 5191 890 5201 924
rect 5075 874 5201 890
rect 5075 852 5105 874
rect 5171 852 5201 874
rect 5267 924 5393 940
rect 5267 890 5278 924
rect 5383 890 5393 924
rect 5267 874 5393 890
rect 5267 852 5297 874
rect 5363 852 5393 874
rect 5459 924 5585 940
rect 5459 890 5470 924
rect 5575 890 5585 924
rect 5459 874 5585 890
rect 5630 930 5702 940
rect 5630 896 5650 930
rect 5684 896 5702 930
rect 5630 874 5702 896
rect 5747 924 5969 940
rect 5747 890 5854 924
rect 5959 890 5969 924
rect 5747 874 5969 890
rect 5459 852 5489 874
rect 5555 852 5585 874
rect 5651 852 5681 874
rect 5747 852 5777 874
rect 5843 852 5873 874
rect 5939 852 5969 874
rect 83 426 113 452
rect 179 426 209 452
rect 275 426 305 452
rect 371 426 401 452
rect 467 426 497 452
rect 563 426 593 452
rect 659 426 689 452
rect 755 426 785 452
rect 851 426 881 452
rect 947 426 977 452
rect 1043 426 1073 452
rect 1139 426 1169 452
rect 1235 426 1265 452
rect 1331 426 1361 452
rect 1427 426 1457 452
rect 1523 426 1553 452
rect 1619 426 1649 452
rect 1715 426 1745 452
rect 1811 426 1841 452
rect 1907 426 1937 452
rect 2003 426 2033 452
rect 2099 426 2129 452
rect 2195 426 2225 452
rect 2291 426 2321 452
rect 2387 426 2417 452
rect 2483 426 2513 452
rect 2579 426 2609 452
rect 2675 426 2705 452
rect 2771 426 2801 452
rect 2867 426 2897 452
rect 2963 426 2993 452
rect 3059 426 3089 452
rect 3155 426 3185 452
rect 3251 426 3281 452
rect 3347 426 3377 452
rect 3443 426 3473 452
rect 3539 426 3569 452
rect 3635 426 3665 452
rect 3731 426 3761 452
rect 3827 426 3857 452
rect 3923 426 3953 452
rect 4019 426 4049 452
rect 4115 426 4145 452
rect 4211 426 4241 452
rect 4307 426 4337 452
rect 4403 426 4433 452
rect 4499 426 4529 452
rect 4595 426 4625 452
rect 4691 426 4721 452
rect 4787 426 4817 452
rect 4883 426 4913 452
rect 4979 426 5009 452
rect 5075 426 5105 452
rect 5171 426 5201 452
rect 5267 426 5297 452
rect 5363 426 5393 452
rect 5459 426 5489 452
rect 5555 426 5585 452
rect 5651 426 5681 452
rect 5747 426 5777 452
rect 5843 426 5873 452
rect 5939 426 5969 452
rect 83 -1872 113 -1846
rect 179 -1872 209 -1846
rect 275 -1872 305 -1846
rect 371 -1872 401 -1846
rect 467 -1872 497 -1846
rect 563 -1872 593 -1846
rect 659 -1872 689 -1846
rect 755 -1872 785 -1846
rect 851 -1872 881 -1846
rect 947 -1872 977 -1846
rect 1043 -1872 1073 -1846
rect 1139 -1872 1169 -1846
rect 1235 -1872 1265 -1846
rect 1331 -1872 1361 -1846
rect 1427 -1872 1457 -1846
rect 1523 -1872 1553 -1846
rect 1619 -1872 1649 -1846
rect 1715 -1872 1745 -1846
rect 1811 -1872 1841 -1846
rect 1907 -1872 1937 -1846
rect 2003 -1872 2033 -1846
rect 2099 -1872 2129 -1846
rect 2195 -1872 2225 -1846
rect 2291 -1872 2321 -1846
rect 2387 -1872 2417 -1846
rect 2483 -1872 2513 -1846
rect 2579 -1872 2609 -1846
rect 2675 -1872 2705 -1846
rect 2771 -1872 2801 -1846
rect 2867 -1872 2897 -1846
rect 2963 -1872 2993 -1846
rect 3059 -1872 3089 -1846
rect 3155 -1872 3185 -1846
rect 3251 -1872 3281 -1846
rect 3347 -1872 3377 -1846
rect 3443 -1872 3473 -1846
rect 3539 -1872 3569 -1846
rect 3635 -1872 3665 -1846
rect 3731 -1872 3761 -1846
rect 3827 -1872 3857 -1846
rect 3923 -1872 3953 -1846
rect 4019 -1872 4049 -1846
rect 4115 -1872 4145 -1846
rect 4211 -1872 4241 -1846
rect 4307 -1872 4337 -1846
rect 4403 -1872 4433 -1846
rect 4499 -1872 4529 -1846
rect 4595 -1872 4625 -1846
rect 4691 -1872 4721 -1846
rect 4787 -1872 4817 -1846
rect 4883 -1872 4913 -1846
rect 4979 -1872 5009 -1846
rect 5075 -1872 5105 -1846
rect 5171 -1872 5201 -1846
rect 5267 -1872 5297 -1846
rect 5363 -1872 5393 -1846
rect 5459 -1872 5489 -1846
rect 5555 -1872 5585 -1846
rect 5651 -1872 5681 -1846
rect 5747 -1872 5777 -1846
rect 5843 -1872 5873 -1846
rect 5939 -1872 5969 -1846
rect 83 -2294 113 -2272
rect 179 -2294 209 -2272
rect 275 -2294 305 -2272
rect 371 -2294 401 -2272
rect 467 -2294 497 -2272
rect 563 -2294 593 -2272
rect 83 -2310 305 -2294
rect 83 -2344 93 -2310
rect 198 -2344 305 -2310
rect 83 -2360 305 -2344
rect 350 -2316 422 -2294
rect 350 -2350 368 -2316
rect 402 -2350 422 -2316
rect 350 -2360 422 -2350
rect 467 -2310 593 -2294
rect 467 -2344 477 -2310
rect 582 -2344 593 -2310
rect 467 -2360 593 -2344
rect 659 -2294 689 -2272
rect 755 -2294 785 -2272
rect 659 -2310 785 -2294
rect 659 -2344 669 -2310
rect 774 -2344 785 -2310
rect 659 -2360 785 -2344
rect 851 -2294 881 -2272
rect 947 -2294 977 -2272
rect 851 -2310 977 -2294
rect 851 -2344 861 -2310
rect 966 -2344 977 -2310
rect 851 -2360 977 -2344
rect 1043 -2294 1073 -2272
rect 1139 -2294 1169 -2272
rect 1043 -2310 1169 -2294
rect 1043 -2344 1053 -2310
rect 1158 -2344 1169 -2310
rect 1043 -2360 1169 -2344
rect 1235 -2294 1265 -2272
rect 1331 -2294 1361 -2272
rect 1235 -2310 1361 -2294
rect 1235 -2344 1245 -2310
rect 1350 -2344 1361 -2310
rect 1235 -2360 1361 -2344
rect 1427 -2294 1457 -2272
rect 1523 -2294 1553 -2272
rect 1427 -2310 1553 -2294
rect 1427 -2344 1437 -2310
rect 1542 -2344 1553 -2310
rect 1427 -2360 1553 -2344
rect 1619 -2294 1649 -2272
rect 1715 -2294 1745 -2272
rect 1619 -2310 1745 -2294
rect 1619 -2344 1630 -2310
rect 1735 -2344 1745 -2310
rect 1619 -2360 1745 -2344
rect 1811 -2294 1841 -2272
rect 1907 -2294 1937 -2272
rect 1811 -2310 1937 -2294
rect 1811 -2344 1822 -2310
rect 1927 -2344 1937 -2310
rect 1811 -2360 1937 -2344
rect 2003 -2294 2033 -2272
rect 2099 -2294 2129 -2272
rect 2003 -2310 2129 -2294
rect 2003 -2344 2014 -2310
rect 2119 -2344 2129 -2310
rect 2003 -2360 2129 -2344
rect 2195 -2294 2225 -2272
rect 2291 -2294 2321 -2272
rect 2195 -2310 2321 -2294
rect 2195 -2344 2206 -2310
rect 2311 -2344 2321 -2310
rect 2195 -2360 2321 -2344
rect 2387 -2294 2417 -2272
rect 2483 -2294 2513 -2272
rect 2387 -2310 2513 -2294
rect 2387 -2344 2398 -2310
rect 2503 -2344 2513 -2310
rect 2387 -2360 2513 -2344
rect 2579 -2294 2609 -2272
rect 2675 -2294 2705 -2272
rect 2771 -2294 2801 -2272
rect 2867 -2294 2897 -2272
rect 2963 -2294 2993 -2272
rect 3059 -2294 3089 -2272
rect 3155 -2294 3185 -2272
rect 3251 -2294 3281 -2272
rect 3347 -2294 3377 -2272
rect 3443 -2294 3473 -2272
rect 2579 -2310 2705 -2294
rect 2579 -2344 2590 -2310
rect 2695 -2344 2705 -2310
rect 2579 -2360 2705 -2344
rect 2750 -2316 2822 -2294
rect 2750 -2350 2770 -2316
rect 2804 -2350 2822 -2316
rect 2750 -2360 2822 -2350
rect 2867 -2310 3185 -2294
rect 2867 -2344 2973 -2310
rect 3079 -2344 3185 -2310
rect 2867 -2360 3185 -2344
rect 3230 -2316 3302 -2294
rect 3230 -2350 3248 -2316
rect 3282 -2350 3302 -2316
rect 3230 -2360 3302 -2350
rect 3347 -2310 3473 -2294
rect 3347 -2344 3357 -2310
rect 3462 -2344 3473 -2310
rect 3347 -2360 3473 -2344
rect 3539 -2294 3569 -2272
rect 3635 -2294 3665 -2272
rect 3539 -2310 3665 -2294
rect 3539 -2344 3549 -2310
rect 3654 -2344 3665 -2310
rect 3539 -2360 3665 -2344
rect 3731 -2294 3761 -2272
rect 3827 -2294 3857 -2272
rect 3731 -2310 3857 -2294
rect 3731 -2344 3741 -2310
rect 3846 -2344 3857 -2310
rect 3731 -2360 3857 -2344
rect 3923 -2294 3953 -2272
rect 4019 -2294 4049 -2272
rect 3923 -2310 4049 -2294
rect 3923 -2344 3933 -2310
rect 4038 -2344 4049 -2310
rect 3923 -2360 4049 -2344
rect 4115 -2294 4145 -2272
rect 4211 -2294 4241 -2272
rect 4115 -2310 4241 -2294
rect 4115 -2344 4125 -2310
rect 4230 -2344 4241 -2310
rect 4115 -2360 4241 -2344
rect 4307 -2294 4337 -2272
rect 4403 -2294 4433 -2272
rect 4307 -2310 4433 -2294
rect 4307 -2344 4317 -2310
rect 4422 -2344 4433 -2310
rect 4307 -2360 4433 -2344
rect 4499 -2294 4529 -2272
rect 4595 -2294 4625 -2272
rect 4499 -2310 4625 -2294
rect 4499 -2344 4510 -2310
rect 4615 -2344 4625 -2310
rect 4499 -2360 4625 -2344
rect 4691 -2294 4721 -2272
rect 4787 -2294 4817 -2272
rect 4691 -2310 4817 -2294
rect 4691 -2344 4702 -2310
rect 4807 -2344 4817 -2310
rect 4691 -2360 4817 -2344
rect 4883 -2294 4913 -2272
rect 4979 -2294 5009 -2272
rect 4883 -2310 5009 -2294
rect 4883 -2344 4894 -2310
rect 4999 -2344 5009 -2310
rect 4883 -2360 5009 -2344
rect 5075 -2294 5105 -2272
rect 5171 -2294 5201 -2272
rect 5075 -2310 5201 -2294
rect 5075 -2344 5086 -2310
rect 5191 -2344 5201 -2310
rect 5075 -2360 5201 -2344
rect 5267 -2294 5297 -2272
rect 5363 -2294 5393 -2272
rect 5267 -2310 5393 -2294
rect 5267 -2344 5278 -2310
rect 5383 -2344 5393 -2310
rect 5267 -2360 5393 -2344
rect 5459 -2294 5489 -2272
rect 5555 -2294 5585 -2272
rect 5651 -2294 5681 -2272
rect 5747 -2294 5777 -2272
rect 5843 -2294 5873 -2272
rect 5939 -2294 5969 -2272
rect 5459 -2310 5585 -2294
rect 5459 -2344 5470 -2310
rect 5575 -2344 5585 -2310
rect 5459 -2360 5585 -2344
rect 5630 -2316 5702 -2294
rect 5630 -2350 5650 -2316
rect 5684 -2350 5702 -2316
rect 5630 -2360 5702 -2350
rect 5747 -2310 5969 -2294
rect 5747 -2344 5854 -2310
rect 5959 -2344 5969 -2310
rect 5747 -2360 5969 -2344
rect 83 -2546 209 -2530
rect 83 -2580 93 -2546
rect 198 -2580 209 -2546
rect 83 -2596 209 -2580
rect 83 -2627 113 -2596
rect 179 -2627 209 -2596
rect 275 -2546 401 -2530
rect 275 -2580 285 -2546
rect 390 -2580 401 -2546
rect 275 -2596 401 -2580
rect 275 -2627 305 -2596
rect 371 -2627 401 -2596
rect 467 -2546 593 -2530
rect 467 -2580 477 -2546
rect 582 -2580 593 -2546
rect 467 -2596 593 -2580
rect 467 -2627 497 -2596
rect 563 -2627 593 -2596
rect 659 -2546 785 -2530
rect 659 -2580 669 -2546
rect 774 -2580 785 -2546
rect 659 -2596 785 -2580
rect 659 -2627 689 -2596
rect 755 -2627 785 -2596
rect 851 -2546 977 -2530
rect 851 -2580 861 -2546
rect 966 -2580 977 -2546
rect 851 -2596 977 -2580
rect 851 -2627 881 -2596
rect 947 -2627 977 -2596
rect 1043 -2546 1169 -2530
rect 1043 -2580 1053 -2546
rect 1158 -2580 1169 -2546
rect 1043 -2596 1169 -2580
rect 1043 -2627 1073 -2596
rect 1139 -2627 1169 -2596
rect 1235 -2546 1361 -2530
rect 1235 -2580 1245 -2546
rect 1350 -2580 1361 -2546
rect 1235 -2596 1361 -2580
rect 1235 -2627 1265 -2596
rect 1331 -2627 1361 -2596
rect 1427 -2546 1553 -2530
rect 1427 -2580 1437 -2546
rect 1542 -2580 1553 -2546
rect 1427 -2596 1553 -2580
rect 1427 -2627 1457 -2596
rect 1523 -2627 1553 -2596
rect 1619 -2546 1745 -2530
rect 1619 -2580 1630 -2546
rect 1735 -2580 1745 -2546
rect 1619 -2596 1745 -2580
rect 1619 -2627 1649 -2596
rect 1715 -2627 1745 -2596
rect 1811 -2546 1937 -2530
rect 1811 -2580 1822 -2546
rect 1927 -2580 1937 -2546
rect 1811 -2596 1937 -2580
rect 1811 -2627 1841 -2596
rect 1907 -2627 1937 -2596
rect 2003 -2546 2129 -2530
rect 2003 -2580 2014 -2546
rect 2119 -2580 2129 -2546
rect 2003 -2596 2129 -2580
rect 2003 -2627 2033 -2596
rect 2099 -2627 2129 -2596
rect 2195 -2546 2321 -2530
rect 2195 -2580 2206 -2546
rect 2311 -2580 2321 -2546
rect 2195 -2596 2321 -2580
rect 2195 -2627 2225 -2596
rect 2291 -2627 2321 -2596
rect 2387 -2546 2513 -2530
rect 2387 -2580 2398 -2546
rect 2503 -2580 2513 -2546
rect 2387 -2596 2513 -2580
rect 2387 -2627 2417 -2596
rect 2483 -2627 2513 -2596
rect 2579 -2546 2705 -2530
rect 2579 -2580 2590 -2546
rect 2695 -2580 2705 -2546
rect 2579 -2596 2705 -2580
rect 2579 -2627 2609 -2596
rect 2675 -2627 2705 -2596
rect 2771 -2546 2897 -2530
rect 2771 -2580 2782 -2546
rect 2887 -2580 2897 -2546
rect 2771 -2596 2897 -2580
rect 2771 -2627 2801 -2596
rect 2867 -2627 2897 -2596
rect 2963 -2546 3089 -2530
rect 2963 -2580 2973 -2546
rect 3079 -2580 3089 -2546
rect 2963 -2596 3089 -2580
rect 2963 -2627 2993 -2596
rect 3059 -2627 3089 -2596
rect 3155 -2546 3281 -2530
rect 3155 -2580 3165 -2546
rect 3270 -2580 3281 -2546
rect 3155 -2596 3281 -2580
rect 3155 -2627 3185 -2596
rect 3251 -2627 3281 -2596
rect 3347 -2546 3473 -2530
rect 3347 -2580 3357 -2546
rect 3462 -2580 3473 -2546
rect 3347 -2596 3473 -2580
rect 3347 -2627 3377 -2596
rect 3443 -2627 3473 -2596
rect 3539 -2546 3665 -2530
rect 3539 -2580 3549 -2546
rect 3654 -2580 3665 -2546
rect 3539 -2596 3665 -2580
rect 3539 -2627 3569 -2596
rect 3635 -2627 3665 -2596
rect 3731 -2546 3857 -2530
rect 3731 -2580 3741 -2546
rect 3846 -2580 3857 -2546
rect 3731 -2596 3857 -2580
rect 3731 -2627 3761 -2596
rect 3827 -2627 3857 -2596
rect 3923 -2546 4049 -2530
rect 3923 -2580 3933 -2546
rect 4038 -2580 4049 -2546
rect 3923 -2596 4049 -2580
rect 3923 -2627 3953 -2596
rect 4019 -2627 4049 -2596
rect 4115 -2546 4241 -2530
rect 4115 -2580 4125 -2546
rect 4230 -2580 4241 -2546
rect 4115 -2596 4241 -2580
rect 4115 -2627 4145 -2596
rect 4211 -2627 4241 -2596
rect 4307 -2546 4433 -2530
rect 4307 -2580 4317 -2546
rect 4422 -2580 4433 -2546
rect 4307 -2596 4433 -2580
rect 4307 -2627 4337 -2596
rect 4403 -2627 4433 -2596
rect 4499 -2546 4625 -2530
rect 4499 -2580 4510 -2546
rect 4615 -2580 4625 -2546
rect 4499 -2596 4625 -2580
rect 4499 -2627 4529 -2596
rect 4595 -2627 4625 -2596
rect 4691 -2546 4817 -2530
rect 4691 -2580 4702 -2546
rect 4807 -2580 4817 -2546
rect 4691 -2596 4817 -2580
rect 4691 -2627 4721 -2596
rect 4787 -2627 4817 -2596
rect 4883 -2546 5009 -2530
rect 4883 -2580 4894 -2546
rect 4999 -2580 5009 -2546
rect 4883 -2596 5009 -2580
rect 4883 -2627 4913 -2596
rect 4979 -2627 5009 -2596
rect 5075 -2546 5201 -2530
rect 5075 -2580 5086 -2546
rect 5191 -2580 5201 -2546
rect 5075 -2596 5201 -2580
rect 5075 -2627 5105 -2596
rect 5171 -2627 5201 -2596
rect 5267 -2546 5393 -2530
rect 5267 -2580 5278 -2546
rect 5383 -2580 5393 -2546
rect 5267 -2596 5393 -2580
rect 5267 -2627 5297 -2596
rect 5363 -2627 5393 -2596
rect 5459 -2546 5585 -2530
rect 5459 -2580 5470 -2546
rect 5575 -2580 5585 -2546
rect 5459 -2596 5585 -2580
rect 5459 -2627 5489 -2596
rect 5555 -2627 5585 -2596
rect 5651 -2546 5777 -2530
rect 5651 -2580 5662 -2546
rect 5767 -2580 5777 -2546
rect 5651 -2596 5777 -2580
rect 5651 -2627 5681 -2596
rect 5747 -2627 5777 -2596
rect 5843 -2546 5969 -2530
rect 5843 -2580 5854 -2546
rect 5959 -2580 5969 -2546
rect 5843 -2596 5969 -2580
rect 5843 -2627 5873 -2596
rect 5939 -2627 5969 -2596
rect 83 -3378 113 -3347
rect 179 -3378 209 -3347
rect 275 -3378 305 -3347
rect 371 -3378 401 -3347
rect 467 -3378 497 -3347
rect 563 -3378 593 -3347
rect 659 -3378 689 -3347
rect 755 -3378 785 -3347
rect 851 -3378 881 -3347
rect 947 -3378 977 -3347
rect 1043 -3378 1073 -3347
rect 1139 -3378 1169 -3347
rect 1235 -3378 1265 -3347
rect 1331 -3378 1361 -3347
rect 1427 -3378 1457 -3347
rect 1523 -3378 1553 -3347
rect 1619 -3378 1649 -3347
rect 1715 -3378 1745 -3347
rect 1811 -3378 1841 -3347
rect 1907 -3378 1937 -3347
rect 2003 -3378 2033 -3347
rect 2099 -3378 2129 -3347
rect 2195 -3378 2225 -3347
rect 2291 -3378 2321 -3347
rect 2387 -3378 2417 -3347
rect 2483 -3378 2513 -3347
rect 2579 -3378 2609 -3347
rect 2675 -3378 2705 -3347
rect 2771 -3378 2801 -3347
rect 2867 -3378 2897 -3347
rect 2963 -3378 2993 -3347
rect 3059 -3378 3089 -3347
rect 3155 -3378 3185 -3347
rect 3251 -3378 3281 -3347
rect 3347 -3378 3377 -3347
rect 3443 -3378 3473 -3347
rect 3539 -3378 3569 -3347
rect 3635 -3378 3665 -3347
rect 3731 -3378 3761 -3347
rect 3827 -3378 3857 -3347
rect 3923 -3378 3953 -3347
rect 4019 -3378 4049 -3347
rect 4115 -3378 4145 -3347
rect 4211 -3378 4241 -3347
rect 4307 -3378 4337 -3347
rect 4403 -3378 4433 -3347
rect 4499 -3378 4529 -3347
rect 4595 -3378 4625 -3347
rect 4691 -3378 4721 -3347
rect 4787 -3378 4817 -3347
rect 4883 -3378 4913 -3347
rect 4979 -3378 5009 -3347
rect 5075 -3378 5105 -3347
rect 5171 -3378 5201 -3347
rect 5267 -3378 5297 -3347
rect 5363 -3378 5393 -3347
rect 5459 -3378 5489 -3347
rect 5555 -3378 5585 -3347
rect 5651 -3378 5681 -3347
rect 5747 -3378 5777 -3347
rect 5843 -3378 5873 -3347
rect 5939 -3378 5969 -3347
<< polycont >>
rect 93 1126 198 1160
rect 285 1126 390 1160
rect 477 1126 582 1160
rect 669 1126 774 1160
rect 861 1126 966 1160
rect 1053 1126 1158 1160
rect 1245 1126 1350 1160
rect 1437 1126 1542 1160
rect 1630 1126 1735 1160
rect 1822 1126 1927 1160
rect 2014 1126 2119 1160
rect 2206 1126 2311 1160
rect 2398 1126 2503 1160
rect 2590 1126 2695 1160
rect 2782 1126 2887 1160
rect 2973 1126 3079 1160
rect 3165 1126 3270 1160
rect 3357 1126 3462 1160
rect 3549 1126 3654 1160
rect 3741 1126 3846 1160
rect 3933 1126 4038 1160
rect 4125 1126 4230 1160
rect 4317 1126 4422 1160
rect 4510 1126 4615 1160
rect 4702 1126 4807 1160
rect 4894 1126 4999 1160
rect 5086 1126 5191 1160
rect 5278 1126 5383 1160
rect 5470 1126 5575 1160
rect 5662 1126 5767 1160
rect 5854 1126 5959 1160
rect 93 890 198 924
rect 368 896 402 930
rect 477 890 582 924
rect 669 890 774 924
rect 861 890 966 924
rect 1053 890 1158 924
rect 1245 890 1350 924
rect 1437 890 1542 924
rect 1630 890 1735 924
rect 1822 890 1927 924
rect 2014 890 2119 924
rect 2206 890 2311 924
rect 2398 890 2503 924
rect 2590 890 2695 924
rect 2770 896 2804 930
rect 2973 890 3079 924
rect 3248 896 3282 930
rect 3357 890 3462 924
rect 3549 890 3654 924
rect 3741 890 3846 924
rect 3933 890 4038 924
rect 4125 890 4230 924
rect 4317 890 4422 924
rect 4510 890 4615 924
rect 4702 890 4807 924
rect 4894 890 4999 924
rect 5086 890 5191 924
rect 5278 890 5383 924
rect 5470 890 5575 924
rect 5650 896 5684 930
rect 5854 890 5959 924
rect 93 -2344 198 -2310
rect 368 -2350 402 -2316
rect 477 -2344 582 -2310
rect 669 -2344 774 -2310
rect 861 -2344 966 -2310
rect 1053 -2344 1158 -2310
rect 1245 -2344 1350 -2310
rect 1437 -2344 1542 -2310
rect 1630 -2344 1735 -2310
rect 1822 -2344 1927 -2310
rect 2014 -2344 2119 -2310
rect 2206 -2344 2311 -2310
rect 2398 -2344 2503 -2310
rect 2590 -2344 2695 -2310
rect 2770 -2350 2804 -2316
rect 2973 -2344 3079 -2310
rect 3248 -2350 3282 -2316
rect 3357 -2344 3462 -2310
rect 3549 -2344 3654 -2310
rect 3741 -2344 3846 -2310
rect 3933 -2344 4038 -2310
rect 4125 -2344 4230 -2310
rect 4317 -2344 4422 -2310
rect 4510 -2344 4615 -2310
rect 4702 -2344 4807 -2310
rect 4894 -2344 4999 -2310
rect 5086 -2344 5191 -2310
rect 5278 -2344 5383 -2310
rect 5470 -2344 5575 -2310
rect 5650 -2350 5684 -2316
rect 5854 -2344 5959 -2310
rect 93 -2580 198 -2546
rect 285 -2580 390 -2546
rect 477 -2580 582 -2546
rect 669 -2580 774 -2546
rect 861 -2580 966 -2546
rect 1053 -2580 1158 -2546
rect 1245 -2580 1350 -2546
rect 1437 -2580 1542 -2546
rect 1630 -2580 1735 -2546
rect 1822 -2580 1927 -2546
rect 2014 -2580 2119 -2546
rect 2206 -2580 2311 -2546
rect 2398 -2580 2503 -2546
rect 2590 -2580 2695 -2546
rect 2782 -2580 2887 -2546
rect 2973 -2580 3079 -2546
rect 3165 -2580 3270 -2546
rect 3357 -2580 3462 -2546
rect 3549 -2580 3654 -2546
rect 3741 -2580 3846 -2546
rect 3933 -2580 4038 -2546
rect 4125 -2580 4230 -2546
rect 4317 -2580 4422 -2546
rect 4510 -2580 4615 -2546
rect 4702 -2580 4807 -2546
rect 4894 -2580 4999 -2546
rect 5086 -2580 5191 -2546
rect 5278 -2580 5383 -2546
rect 5470 -2580 5575 -2546
rect 5662 -2580 5767 -2546
rect 5854 -2580 5959 -2546
<< locali >>
rect 26 2024 126 2058
rect 5926 2024 6026 2058
rect 33 1915 67 1931
rect 33 1203 67 1219
rect 129 1915 163 1931
rect 129 1203 163 1219
rect 225 1915 259 1931
rect 225 1203 259 1219
rect 321 1915 355 1931
rect 321 1203 355 1219
rect 417 1915 451 1931
rect 417 1203 451 1219
rect 513 1915 547 1931
rect 513 1203 547 1219
rect 609 1915 643 1931
rect 609 1203 643 1219
rect 705 1915 739 1931
rect 705 1203 739 1219
rect 801 1915 835 1931
rect 801 1203 835 1219
rect 897 1915 931 1931
rect 897 1203 931 1219
rect 993 1915 1027 1931
rect 993 1203 1027 1219
rect 1089 1915 1123 1931
rect 1089 1203 1123 1219
rect 1185 1915 1219 1931
rect 1185 1203 1219 1219
rect 1281 1915 1315 1931
rect 1281 1203 1315 1219
rect 1377 1915 1411 1931
rect 1377 1203 1411 1219
rect 1473 1915 1507 1931
rect 1473 1203 1507 1219
rect 1569 1915 1603 1931
rect 1569 1203 1603 1219
rect 1665 1915 1699 1931
rect 1665 1203 1699 1219
rect 1761 1915 1795 1931
rect 1761 1203 1795 1219
rect 1857 1915 1891 1931
rect 1857 1203 1891 1219
rect 1953 1915 1987 1931
rect 1953 1203 1987 1219
rect 2049 1915 2083 1931
rect 2049 1203 2083 1219
rect 2145 1915 2179 1931
rect 2145 1203 2179 1219
rect 2241 1915 2275 1931
rect 2241 1203 2275 1219
rect 2337 1915 2371 1931
rect 2337 1203 2371 1219
rect 2433 1915 2467 1931
rect 2433 1203 2467 1219
rect 2529 1915 2563 1931
rect 2529 1203 2563 1219
rect 2625 1915 2659 1931
rect 2625 1203 2659 1219
rect 2721 1915 2755 1931
rect 2721 1203 2755 1219
rect 2817 1915 2851 1931
rect 2817 1203 2851 1219
rect 2913 1915 2947 1931
rect 2913 1203 2947 1219
rect 3009 1915 3043 1931
rect 3009 1203 3043 1219
rect 3105 1915 3139 1931
rect 3105 1203 3139 1219
rect 3201 1915 3235 1931
rect 3201 1203 3235 1219
rect 3297 1915 3331 1931
rect 3297 1203 3331 1219
rect 3393 1915 3427 1931
rect 3393 1203 3427 1219
rect 3489 1915 3523 1931
rect 3489 1203 3523 1219
rect 3585 1915 3619 1931
rect 3585 1203 3619 1219
rect 3681 1915 3715 1931
rect 3681 1203 3715 1219
rect 3777 1915 3811 1931
rect 3777 1203 3811 1219
rect 3873 1915 3907 1931
rect 3873 1203 3907 1219
rect 3969 1915 4003 1931
rect 3969 1203 4003 1219
rect 4065 1915 4099 1931
rect 4065 1203 4099 1219
rect 4161 1915 4195 1931
rect 4161 1203 4195 1219
rect 4257 1915 4291 1931
rect 4257 1203 4291 1219
rect 4353 1915 4387 1931
rect 4353 1203 4387 1219
rect 4449 1915 4483 1931
rect 4449 1203 4483 1219
rect 4545 1915 4579 1931
rect 4545 1203 4579 1219
rect 4641 1915 4675 1931
rect 4641 1203 4675 1219
rect 4737 1915 4771 1931
rect 4737 1203 4771 1219
rect 4833 1915 4867 1931
rect 4833 1203 4867 1219
rect 4929 1915 4963 1931
rect 4929 1203 4963 1219
rect 5025 1915 5059 1931
rect 5025 1203 5059 1219
rect 5121 1915 5155 1931
rect 5121 1203 5155 1219
rect 5217 1915 5251 1931
rect 5217 1203 5251 1219
rect 5313 1915 5347 1931
rect 5313 1203 5347 1219
rect 5409 1915 5443 1931
rect 5409 1203 5443 1219
rect 5505 1915 5539 1931
rect 5505 1203 5539 1219
rect 5601 1915 5635 1931
rect 5601 1203 5635 1219
rect 5697 1915 5731 1931
rect 5697 1203 5731 1219
rect 5793 1915 5827 1931
rect 5793 1203 5827 1219
rect 5889 1915 5923 1931
rect 5889 1203 5923 1219
rect 5985 1915 6019 1931
rect 5985 1203 6019 1219
rect 77 1126 93 1160
rect 198 1126 214 1160
rect 269 1126 285 1160
rect 390 1126 406 1160
rect 461 1126 477 1160
rect 582 1126 598 1160
rect 653 1126 669 1160
rect 774 1126 790 1160
rect 845 1126 861 1160
rect 966 1126 982 1160
rect 1037 1126 1053 1160
rect 1158 1126 1174 1160
rect 1229 1126 1245 1160
rect 1350 1126 1366 1160
rect 1421 1126 1437 1160
rect 1542 1126 1558 1160
rect 1614 1126 1630 1160
rect 1735 1126 1751 1160
rect 1806 1126 1822 1160
rect 1927 1126 1943 1160
rect 1998 1126 2014 1160
rect 2119 1126 2135 1160
rect 2190 1126 2206 1160
rect 2311 1126 2327 1160
rect 2382 1126 2398 1160
rect 2503 1126 2519 1160
rect 2574 1126 2590 1160
rect 2695 1126 2711 1160
rect 2766 1126 2782 1160
rect 2887 1126 2903 1160
rect 2957 1126 2973 1160
rect 3079 1126 3095 1160
rect 3149 1126 3165 1160
rect 3270 1126 3286 1160
rect 3341 1126 3357 1160
rect 3462 1126 3478 1160
rect 3533 1126 3549 1160
rect 3654 1126 3670 1160
rect 3725 1126 3741 1160
rect 3846 1126 3862 1160
rect 3917 1126 3933 1160
rect 4038 1126 4054 1160
rect 4109 1126 4125 1160
rect 4230 1126 4246 1160
rect 4301 1126 4317 1160
rect 4422 1126 4438 1160
rect 4494 1126 4510 1160
rect 4615 1126 4631 1160
rect 4686 1126 4702 1160
rect 4807 1126 4823 1160
rect 4878 1126 4894 1160
rect 4999 1126 5015 1160
rect 5070 1126 5086 1160
rect 5191 1126 5207 1160
rect 5262 1126 5278 1160
rect 5383 1126 5399 1160
rect 5454 1126 5470 1160
rect 5575 1126 5591 1160
rect 5646 1126 5662 1160
rect 5767 1126 5783 1160
rect 5838 1126 5854 1160
rect 5959 1126 5975 1160
rect 116 1120 128 1126
rect 162 1120 174 1126
rect 116 1110 174 1120
rect 308 1120 320 1126
rect 354 1120 366 1126
rect 308 1110 366 1120
rect 500 1120 512 1126
rect 546 1120 558 1126
rect 500 1082 558 1120
rect 500 1048 512 1082
rect 546 1048 558 1082
rect 500 1042 558 1048
rect 692 1120 704 1126
rect 738 1120 750 1126
rect 692 1082 750 1120
rect 692 1048 704 1082
rect 738 1048 750 1082
rect 692 1042 750 1048
rect 884 1120 896 1126
rect 930 1120 942 1126
rect 884 1082 942 1120
rect 884 1048 896 1082
rect 930 1048 942 1082
rect 884 1042 942 1048
rect 1076 1120 1088 1126
rect 1122 1120 1134 1126
rect 1076 1082 1134 1120
rect 1076 1048 1088 1082
rect 1122 1048 1134 1082
rect 1076 1042 1134 1048
rect 1268 1120 1280 1126
rect 1314 1120 1326 1126
rect 1268 1082 1326 1120
rect 1268 1048 1280 1082
rect 1314 1048 1326 1082
rect 1268 1042 1326 1048
rect 1460 1120 1472 1126
rect 1506 1120 1518 1126
rect 1460 1082 1518 1120
rect 1460 1048 1472 1082
rect 1506 1048 1518 1082
rect 1460 1042 1518 1048
rect 1654 1120 1666 1126
rect 1700 1120 1712 1126
rect 1654 1082 1712 1120
rect 1654 1048 1666 1082
rect 1700 1048 1712 1082
rect 1654 1042 1712 1048
rect 1846 1120 1858 1126
rect 1892 1120 1904 1126
rect 1846 1082 1904 1120
rect 1846 1048 1858 1082
rect 1892 1048 1904 1082
rect 1846 1042 1904 1048
rect 2038 1120 2050 1126
rect 2084 1120 2096 1126
rect 2038 1082 2096 1120
rect 2038 1048 2050 1082
rect 2084 1048 2096 1082
rect 2038 1042 2096 1048
rect 2230 1120 2242 1126
rect 2276 1120 2288 1126
rect 2230 1082 2288 1120
rect 2230 1048 2242 1082
rect 2276 1048 2288 1082
rect 2230 1042 2288 1048
rect 2422 1120 2434 1126
rect 2468 1120 2480 1126
rect 2422 1082 2480 1120
rect 2422 1048 2434 1082
rect 2468 1048 2480 1082
rect 2422 1042 2480 1048
rect 2614 1120 2626 1126
rect 2660 1120 2672 1126
rect 2614 1082 2672 1120
rect 2806 1120 2818 1126
rect 2852 1120 2864 1126
rect 2806 1110 2864 1120
rect 2996 1120 3008 1126
rect 3044 1120 3056 1126
rect 2996 1110 3056 1120
rect 3188 1120 3200 1126
rect 3234 1120 3246 1126
rect 3188 1110 3246 1120
rect 3380 1120 3392 1126
rect 3426 1120 3438 1126
rect 2614 1048 2626 1082
rect 2660 1048 2672 1082
rect 2614 1042 2672 1048
rect 3380 1082 3438 1120
rect 3380 1048 3392 1082
rect 3426 1048 3438 1082
rect 3380 1042 3438 1048
rect 3572 1120 3584 1126
rect 3618 1120 3630 1126
rect 3572 1082 3630 1120
rect 3572 1048 3584 1082
rect 3618 1048 3630 1082
rect 3572 1042 3630 1048
rect 3764 1120 3776 1126
rect 3810 1120 3822 1126
rect 3764 1082 3822 1120
rect 3764 1048 3776 1082
rect 3810 1048 3822 1082
rect 3764 1042 3822 1048
rect 3956 1120 3968 1126
rect 4002 1120 4014 1126
rect 3956 1082 4014 1120
rect 3956 1048 3968 1082
rect 4002 1048 4014 1082
rect 3956 1042 4014 1048
rect 4148 1120 4160 1126
rect 4194 1120 4206 1126
rect 4148 1082 4206 1120
rect 4148 1048 4160 1082
rect 4194 1048 4206 1082
rect 4148 1042 4206 1048
rect 4340 1120 4352 1126
rect 4386 1120 4398 1126
rect 4340 1082 4398 1120
rect 4340 1048 4352 1082
rect 4386 1048 4398 1082
rect 4340 1042 4398 1048
rect 4534 1120 4546 1126
rect 4580 1120 4592 1126
rect 4534 1082 4592 1120
rect 4534 1048 4546 1082
rect 4580 1048 4592 1082
rect 4534 1042 4592 1048
rect 4726 1120 4738 1126
rect 4772 1120 4784 1126
rect 4726 1082 4784 1120
rect 4726 1048 4738 1082
rect 4772 1048 4784 1082
rect 4726 1042 4784 1048
rect 4918 1120 4930 1126
rect 4964 1120 4976 1126
rect 4918 1082 4976 1120
rect 4918 1048 4930 1082
rect 4964 1048 4976 1082
rect 4918 1042 4976 1048
rect 5110 1120 5122 1126
rect 5156 1120 5168 1126
rect 5110 1082 5168 1120
rect 5110 1048 5122 1082
rect 5156 1048 5168 1082
rect 5110 1042 5168 1048
rect 5302 1120 5314 1126
rect 5348 1120 5360 1126
rect 5302 1082 5360 1120
rect 5302 1048 5314 1082
rect 5348 1048 5360 1082
rect 5302 1042 5360 1048
rect 5494 1120 5506 1126
rect 5540 1120 5552 1126
rect 5494 1082 5552 1120
rect 5686 1120 5698 1126
rect 5732 1120 5744 1126
rect 5686 1110 5744 1120
rect 5878 1120 5890 1126
rect 5924 1120 5936 1126
rect 5878 1110 5936 1120
rect 5494 1048 5506 1082
rect 5540 1048 5552 1082
rect 5494 1042 5552 1048
rect 350 1002 422 1008
rect 350 968 368 1002
rect 402 968 422 1002
rect 116 930 174 940
rect 116 924 128 930
rect 162 924 174 930
rect 350 930 422 968
rect 77 890 93 924
rect 198 890 214 924
rect 350 896 368 930
rect 402 896 422 930
rect 500 1002 558 1008
rect 500 968 512 1002
rect 546 968 558 1002
rect 500 930 558 968
rect 500 924 512 930
rect 546 924 558 930
rect 692 1002 750 1008
rect 692 968 704 1002
rect 738 968 750 1002
rect 692 930 750 968
rect 692 924 704 930
rect 738 924 750 930
rect 884 1002 942 1008
rect 884 968 896 1002
rect 930 968 942 1002
rect 884 930 942 968
rect 884 924 896 930
rect 930 924 942 930
rect 1076 1002 1134 1008
rect 1076 968 1088 1002
rect 1122 968 1134 1002
rect 1076 930 1134 968
rect 1076 924 1088 930
rect 1122 924 1134 930
rect 1268 1002 1326 1008
rect 1268 968 1280 1002
rect 1314 968 1326 1002
rect 1268 930 1326 968
rect 1268 924 1280 930
rect 1314 924 1326 930
rect 1460 1002 1518 1008
rect 1460 968 1472 1002
rect 1506 968 1518 1002
rect 1460 930 1518 968
rect 1460 924 1472 930
rect 1506 924 1518 930
rect 1654 1002 1712 1008
rect 1654 968 1666 1002
rect 1700 968 1712 1002
rect 1654 930 1712 968
rect 1654 924 1666 930
rect 1700 924 1712 930
rect 1846 1002 1904 1008
rect 1846 968 1858 1002
rect 1892 968 1904 1002
rect 1846 930 1904 968
rect 1846 924 1858 930
rect 1892 924 1904 930
rect 2038 1002 2096 1008
rect 2038 968 2050 1002
rect 2084 968 2096 1002
rect 2038 930 2096 968
rect 2038 924 2050 930
rect 2084 924 2096 930
rect 2230 1002 2288 1008
rect 2230 968 2242 1002
rect 2276 968 2288 1002
rect 2230 930 2288 968
rect 2230 924 2242 930
rect 2276 924 2288 930
rect 2422 1002 2480 1008
rect 2422 968 2434 1002
rect 2468 968 2480 1002
rect 2422 930 2480 968
rect 2422 924 2434 930
rect 2468 924 2480 930
rect 2614 1002 2672 1008
rect 2614 968 2626 1002
rect 2660 968 2672 1002
rect 2614 930 2672 968
rect 2614 924 2626 930
rect 2660 924 2672 930
rect 2750 1002 2822 1008
rect 2750 968 2770 1002
rect 2804 968 2822 1002
rect 2750 930 2822 968
rect 3230 1002 3302 1008
rect 3230 968 3248 1002
rect 3282 968 3302 1002
rect 350 890 422 896
rect 461 890 477 924
rect 582 890 598 924
rect 653 890 669 924
rect 774 890 790 924
rect 845 890 861 924
rect 966 890 982 924
rect 1037 890 1053 924
rect 1158 890 1174 924
rect 1229 890 1245 924
rect 1350 890 1366 924
rect 1421 890 1437 924
rect 1542 890 1558 924
rect 1614 890 1630 924
rect 1735 890 1751 924
rect 1806 890 1822 924
rect 1927 890 1943 924
rect 1998 890 2014 924
rect 2119 890 2135 924
rect 2190 890 2206 924
rect 2311 890 2327 924
rect 2382 890 2398 924
rect 2503 890 2519 924
rect 2574 890 2590 924
rect 2695 890 2711 924
rect 2750 896 2770 930
rect 2804 896 2822 930
rect 2996 930 3056 940
rect 2996 924 3008 930
rect 3044 924 3056 930
rect 3230 930 3302 968
rect 2750 890 2822 896
rect 2957 890 2973 924
rect 3079 890 3095 924
rect 3230 896 3248 930
rect 3282 896 3302 930
rect 3380 1002 3438 1008
rect 3380 968 3392 1002
rect 3426 968 3438 1002
rect 3380 930 3438 968
rect 3380 924 3392 930
rect 3426 924 3438 930
rect 3572 1002 3630 1008
rect 3572 968 3584 1002
rect 3618 968 3630 1002
rect 3572 930 3630 968
rect 3572 924 3584 930
rect 3618 924 3630 930
rect 3764 1002 3822 1008
rect 3764 968 3776 1002
rect 3810 968 3822 1002
rect 3764 930 3822 968
rect 3764 924 3776 930
rect 3810 924 3822 930
rect 3956 1002 4014 1008
rect 3956 968 3968 1002
rect 4002 968 4014 1002
rect 3956 930 4014 968
rect 3956 924 3968 930
rect 4002 924 4014 930
rect 4148 1002 4206 1008
rect 4148 968 4160 1002
rect 4194 968 4206 1002
rect 4148 930 4206 968
rect 4148 924 4160 930
rect 4194 924 4206 930
rect 4340 1002 4398 1008
rect 4340 968 4352 1002
rect 4386 968 4398 1002
rect 4340 930 4398 968
rect 4340 924 4352 930
rect 4386 924 4398 930
rect 4534 1002 4592 1008
rect 4534 968 4546 1002
rect 4580 968 4592 1002
rect 4534 930 4592 968
rect 4534 924 4546 930
rect 4580 924 4592 930
rect 4726 1002 4784 1008
rect 4726 968 4738 1002
rect 4772 968 4784 1002
rect 4726 930 4784 968
rect 4726 924 4738 930
rect 4772 924 4784 930
rect 4918 1002 4976 1008
rect 4918 968 4930 1002
rect 4964 968 4976 1002
rect 4918 930 4976 968
rect 4918 924 4930 930
rect 4964 924 4976 930
rect 5110 1002 5168 1008
rect 5110 968 5122 1002
rect 5156 968 5168 1002
rect 5110 930 5168 968
rect 5110 924 5122 930
rect 5156 924 5168 930
rect 5302 1002 5360 1008
rect 5302 968 5314 1002
rect 5348 968 5360 1002
rect 5302 930 5360 968
rect 5302 924 5314 930
rect 5348 924 5360 930
rect 5494 1002 5552 1008
rect 5494 968 5506 1002
rect 5540 968 5552 1002
rect 5494 930 5552 968
rect 5494 924 5506 930
rect 5540 924 5552 930
rect 5630 1002 5702 1008
rect 5630 968 5650 1002
rect 5684 968 5702 1002
rect 5630 930 5702 968
rect 3230 890 3302 896
rect 3341 890 3357 924
rect 3462 890 3478 924
rect 3533 890 3549 924
rect 3654 890 3670 924
rect 3725 890 3741 924
rect 3846 890 3862 924
rect 3917 890 3933 924
rect 4038 890 4054 924
rect 4109 890 4125 924
rect 4230 890 4246 924
rect 4301 890 4317 924
rect 4422 890 4438 924
rect 4494 890 4510 924
rect 4615 890 4631 924
rect 4686 890 4702 924
rect 4807 890 4823 924
rect 4878 890 4894 924
rect 4999 890 5015 924
rect 5070 890 5086 924
rect 5191 890 5207 924
rect 5262 890 5278 924
rect 5383 890 5399 924
rect 5454 890 5470 924
rect 5575 890 5591 924
rect 5630 896 5650 930
rect 5684 896 5702 930
rect 5878 930 5936 940
rect 5878 924 5890 930
rect 5924 924 5936 930
rect 5630 890 5702 896
rect 5838 890 5854 924
rect 5959 890 5975 924
rect 33 840 67 856
rect 33 448 67 464
rect 129 840 163 856
rect 129 448 163 464
rect 225 840 259 856
rect 225 448 259 464
rect 321 840 355 856
rect 321 448 355 464
rect 417 840 451 856
rect 417 448 451 464
rect 513 840 547 856
rect 513 448 547 464
rect 609 840 643 856
rect 609 448 643 464
rect 705 840 739 856
rect 705 448 739 464
rect 801 840 835 856
rect 801 448 835 464
rect 897 840 931 856
rect 897 448 931 464
rect 993 840 1027 856
rect 993 448 1027 464
rect 1089 840 1123 856
rect 1089 448 1123 464
rect 1185 840 1219 856
rect 1185 448 1219 464
rect 1281 840 1315 856
rect 1281 448 1315 464
rect 1377 840 1411 856
rect 1377 448 1411 464
rect 1473 840 1507 856
rect 1473 448 1507 464
rect 1569 840 1603 856
rect 1569 448 1603 464
rect 1665 840 1699 856
rect 1665 448 1699 464
rect 1761 840 1795 856
rect 1761 448 1795 464
rect 1857 840 1891 856
rect 1857 448 1891 464
rect 1953 840 1987 856
rect 1953 448 1987 464
rect 2049 840 2083 856
rect 2049 448 2083 464
rect 2145 840 2179 856
rect 2145 448 2179 464
rect 2241 840 2275 856
rect 2241 448 2275 464
rect 2337 840 2371 856
rect 2337 448 2371 464
rect 2433 840 2467 856
rect 2433 448 2467 464
rect 2529 840 2563 856
rect 2529 448 2563 464
rect 2625 840 2659 856
rect 2625 448 2659 464
rect 2721 840 2755 856
rect 2721 448 2755 464
rect 2817 840 2851 856
rect 2817 448 2851 464
rect 2913 840 2947 856
rect 2913 448 2947 464
rect 3009 840 3043 856
rect 3009 448 3043 464
rect 3105 840 3139 856
rect 3105 448 3139 464
rect 3201 840 3235 856
rect 3201 448 3235 464
rect 3297 840 3331 856
rect 3297 448 3331 464
rect 3393 840 3427 856
rect 3393 448 3427 464
rect 3489 840 3523 856
rect 3489 448 3523 464
rect 3585 840 3619 856
rect 3585 448 3619 464
rect 3681 840 3715 856
rect 3681 448 3715 464
rect 3777 840 3811 856
rect 3777 448 3811 464
rect 3873 840 3907 856
rect 3873 448 3907 464
rect 3969 840 4003 856
rect 3969 448 4003 464
rect 4065 840 4099 856
rect 4065 448 4099 464
rect 4161 840 4195 856
rect 4161 448 4195 464
rect 4257 840 4291 856
rect 4257 448 4291 464
rect 4353 840 4387 856
rect 4353 448 4387 464
rect 4449 840 4483 856
rect 4449 448 4483 464
rect 4545 840 4579 856
rect 4545 448 4579 464
rect 4641 840 4675 856
rect 4641 448 4675 464
rect 4737 840 4771 856
rect 4737 448 4771 464
rect 4833 840 4867 856
rect 4833 448 4867 464
rect 4929 840 4963 856
rect 4929 448 4963 464
rect 5025 840 5059 856
rect 5025 448 5059 464
rect 5121 840 5155 856
rect 5121 448 5155 464
rect 5217 840 5251 856
rect 5217 448 5251 464
rect 5313 840 5347 856
rect 5313 448 5347 464
rect 5409 840 5443 856
rect 5409 448 5443 464
rect 5505 840 5539 856
rect 5505 448 5539 464
rect 5601 840 5635 856
rect 5601 448 5635 464
rect 5697 840 5731 856
rect 5697 448 5731 464
rect 5793 840 5827 856
rect 5793 448 5827 464
rect 5889 840 5923 856
rect 5889 448 5923 464
rect 5985 840 6019 856
rect 5985 448 6019 464
rect 26 322 126 356
rect 5926 322 6026 356
rect 26 -1776 126 -1742
rect 5926 -1776 6026 -1742
rect 33 -1884 67 -1868
rect 33 -2276 67 -2260
rect 129 -1884 163 -1868
rect 129 -2276 163 -2260
rect 225 -1884 259 -1868
rect 225 -2276 259 -2260
rect 321 -1884 355 -1868
rect 321 -2276 355 -2260
rect 417 -1884 451 -1868
rect 417 -2276 451 -2260
rect 513 -1884 547 -1868
rect 513 -2276 547 -2260
rect 609 -1884 643 -1868
rect 609 -2276 643 -2260
rect 705 -1884 739 -1868
rect 705 -2276 739 -2260
rect 801 -1884 835 -1868
rect 801 -2276 835 -2260
rect 897 -1884 931 -1868
rect 897 -2276 931 -2260
rect 993 -1884 1027 -1868
rect 993 -2276 1027 -2260
rect 1089 -1884 1123 -1868
rect 1089 -2276 1123 -2260
rect 1185 -1884 1219 -1868
rect 1185 -2276 1219 -2260
rect 1281 -1884 1315 -1868
rect 1281 -2276 1315 -2260
rect 1377 -1884 1411 -1868
rect 1377 -2276 1411 -2260
rect 1473 -1884 1507 -1868
rect 1473 -2276 1507 -2260
rect 1569 -1884 1603 -1868
rect 1569 -2276 1603 -2260
rect 1665 -1884 1699 -1868
rect 1665 -2276 1699 -2260
rect 1761 -1884 1795 -1868
rect 1761 -2276 1795 -2260
rect 1857 -1884 1891 -1868
rect 1857 -2276 1891 -2260
rect 1953 -1884 1987 -1868
rect 1953 -2276 1987 -2260
rect 2049 -1884 2083 -1868
rect 2049 -2276 2083 -2260
rect 2145 -1884 2179 -1868
rect 2145 -2276 2179 -2260
rect 2241 -1884 2275 -1868
rect 2241 -2276 2275 -2260
rect 2337 -1884 2371 -1868
rect 2337 -2276 2371 -2260
rect 2433 -1884 2467 -1868
rect 2433 -2276 2467 -2260
rect 2529 -1884 2563 -1868
rect 2529 -2276 2563 -2260
rect 2625 -1884 2659 -1868
rect 2625 -2276 2659 -2260
rect 2721 -1884 2755 -1868
rect 2721 -2276 2755 -2260
rect 2817 -1884 2851 -1868
rect 2817 -2276 2851 -2260
rect 2913 -1884 2947 -1868
rect 2913 -2276 2947 -2260
rect 3009 -1884 3043 -1868
rect 3009 -2276 3043 -2260
rect 3105 -1884 3139 -1868
rect 3105 -2276 3139 -2260
rect 3201 -1884 3235 -1868
rect 3201 -2276 3235 -2260
rect 3297 -1884 3331 -1868
rect 3297 -2276 3331 -2260
rect 3393 -1884 3427 -1868
rect 3393 -2276 3427 -2260
rect 3489 -1884 3523 -1868
rect 3489 -2276 3523 -2260
rect 3585 -1884 3619 -1868
rect 3585 -2276 3619 -2260
rect 3681 -1884 3715 -1868
rect 3681 -2276 3715 -2260
rect 3777 -1884 3811 -1868
rect 3777 -2276 3811 -2260
rect 3873 -1884 3907 -1868
rect 3873 -2276 3907 -2260
rect 3969 -1884 4003 -1868
rect 3969 -2276 4003 -2260
rect 4065 -1884 4099 -1868
rect 4065 -2276 4099 -2260
rect 4161 -1884 4195 -1868
rect 4161 -2276 4195 -2260
rect 4257 -1884 4291 -1868
rect 4257 -2276 4291 -2260
rect 4353 -1884 4387 -1868
rect 4353 -2276 4387 -2260
rect 4449 -1884 4483 -1868
rect 4449 -2276 4483 -2260
rect 4545 -1884 4579 -1868
rect 4545 -2276 4579 -2260
rect 4641 -1884 4675 -1868
rect 4641 -2276 4675 -2260
rect 4737 -1884 4771 -1868
rect 4737 -2276 4771 -2260
rect 4833 -1884 4867 -1868
rect 4833 -2276 4867 -2260
rect 4929 -1884 4963 -1868
rect 4929 -2276 4963 -2260
rect 5025 -1884 5059 -1868
rect 5025 -2276 5059 -2260
rect 5121 -1884 5155 -1868
rect 5121 -2276 5155 -2260
rect 5217 -1884 5251 -1868
rect 5217 -2276 5251 -2260
rect 5313 -1884 5347 -1868
rect 5313 -2276 5347 -2260
rect 5409 -1884 5443 -1868
rect 5409 -2276 5443 -2260
rect 5505 -1884 5539 -1868
rect 5505 -2276 5539 -2260
rect 5601 -1884 5635 -1868
rect 5601 -2276 5635 -2260
rect 5697 -1884 5731 -1868
rect 5697 -2276 5731 -2260
rect 5793 -1884 5827 -1868
rect 5793 -2276 5827 -2260
rect 5889 -1884 5923 -1868
rect 5889 -2276 5923 -2260
rect 5985 -1884 6019 -1868
rect 5985 -2276 6019 -2260
rect 77 -2344 93 -2310
rect 198 -2344 214 -2310
rect 350 -2316 422 -2310
rect 116 -2350 128 -2344
rect 162 -2350 174 -2344
rect 116 -2360 174 -2350
rect 350 -2350 368 -2316
rect 402 -2350 422 -2316
rect 461 -2344 477 -2310
rect 582 -2344 598 -2310
rect 653 -2344 669 -2310
rect 774 -2344 790 -2310
rect 845 -2344 861 -2310
rect 966 -2344 982 -2310
rect 1037 -2344 1053 -2310
rect 1158 -2344 1174 -2310
rect 1229 -2344 1245 -2310
rect 1350 -2344 1366 -2310
rect 1421 -2344 1437 -2310
rect 1542 -2344 1558 -2310
rect 1614 -2344 1630 -2310
rect 1735 -2344 1751 -2310
rect 1806 -2344 1822 -2310
rect 1927 -2344 1943 -2310
rect 1998 -2344 2014 -2310
rect 2119 -2344 2135 -2310
rect 2190 -2344 2206 -2310
rect 2311 -2344 2327 -2310
rect 2382 -2344 2398 -2310
rect 2503 -2344 2519 -2310
rect 2574 -2344 2590 -2310
rect 2695 -2344 2711 -2310
rect 2750 -2316 2822 -2310
rect 350 -2388 422 -2350
rect 350 -2422 368 -2388
rect 402 -2422 422 -2388
rect 350 -2428 422 -2422
rect 500 -2350 512 -2344
rect 546 -2350 558 -2344
rect 500 -2388 558 -2350
rect 500 -2422 512 -2388
rect 546 -2422 558 -2388
rect 500 -2428 558 -2422
rect 692 -2350 704 -2344
rect 738 -2350 750 -2344
rect 692 -2388 750 -2350
rect 692 -2422 704 -2388
rect 738 -2422 750 -2388
rect 692 -2428 750 -2422
rect 884 -2350 896 -2344
rect 930 -2350 942 -2344
rect 884 -2388 942 -2350
rect 884 -2422 896 -2388
rect 930 -2422 942 -2388
rect 884 -2428 942 -2422
rect 1076 -2350 1088 -2344
rect 1122 -2350 1134 -2344
rect 1076 -2388 1134 -2350
rect 1076 -2422 1088 -2388
rect 1122 -2422 1134 -2388
rect 1076 -2428 1134 -2422
rect 1268 -2350 1280 -2344
rect 1314 -2350 1326 -2344
rect 1268 -2388 1326 -2350
rect 1268 -2422 1280 -2388
rect 1314 -2422 1326 -2388
rect 1268 -2428 1326 -2422
rect 1460 -2350 1472 -2344
rect 1506 -2350 1518 -2344
rect 1460 -2388 1518 -2350
rect 1460 -2422 1472 -2388
rect 1506 -2422 1518 -2388
rect 1460 -2428 1518 -2422
rect 1654 -2350 1666 -2344
rect 1700 -2350 1712 -2344
rect 1654 -2388 1712 -2350
rect 1654 -2422 1666 -2388
rect 1700 -2422 1712 -2388
rect 1654 -2428 1712 -2422
rect 1846 -2350 1858 -2344
rect 1892 -2350 1904 -2344
rect 1846 -2388 1904 -2350
rect 1846 -2422 1858 -2388
rect 1892 -2422 1904 -2388
rect 1846 -2428 1904 -2422
rect 2038 -2350 2050 -2344
rect 2084 -2350 2096 -2344
rect 2038 -2388 2096 -2350
rect 2038 -2422 2050 -2388
rect 2084 -2422 2096 -2388
rect 2038 -2428 2096 -2422
rect 2230 -2350 2242 -2344
rect 2276 -2350 2288 -2344
rect 2230 -2388 2288 -2350
rect 2230 -2422 2242 -2388
rect 2276 -2422 2288 -2388
rect 2230 -2428 2288 -2422
rect 2422 -2350 2434 -2344
rect 2468 -2350 2480 -2344
rect 2422 -2388 2480 -2350
rect 2422 -2422 2434 -2388
rect 2468 -2422 2480 -2388
rect 2422 -2428 2480 -2422
rect 2614 -2350 2626 -2344
rect 2660 -2350 2672 -2344
rect 2614 -2388 2672 -2350
rect 2614 -2422 2626 -2388
rect 2660 -2422 2672 -2388
rect 2614 -2428 2672 -2422
rect 2750 -2350 2770 -2316
rect 2804 -2350 2822 -2316
rect 2957 -2344 2973 -2310
rect 3079 -2344 3095 -2310
rect 3230 -2316 3302 -2310
rect 2750 -2388 2822 -2350
rect 2996 -2350 3008 -2344
rect 3044 -2350 3056 -2344
rect 2996 -2360 3056 -2350
rect 3230 -2350 3248 -2316
rect 3282 -2350 3302 -2316
rect 3341 -2344 3357 -2310
rect 3462 -2344 3478 -2310
rect 3533 -2344 3549 -2310
rect 3654 -2344 3670 -2310
rect 3725 -2344 3741 -2310
rect 3846 -2344 3862 -2310
rect 3917 -2344 3933 -2310
rect 4038 -2344 4054 -2310
rect 4109 -2344 4125 -2310
rect 4230 -2344 4246 -2310
rect 4301 -2344 4317 -2310
rect 4422 -2344 4438 -2310
rect 4494 -2344 4510 -2310
rect 4615 -2344 4631 -2310
rect 4686 -2344 4702 -2310
rect 4807 -2344 4823 -2310
rect 4878 -2344 4894 -2310
rect 4999 -2344 5015 -2310
rect 5070 -2344 5086 -2310
rect 5191 -2344 5207 -2310
rect 5262 -2344 5278 -2310
rect 5383 -2344 5399 -2310
rect 5454 -2344 5470 -2310
rect 5575 -2344 5591 -2310
rect 5630 -2316 5702 -2310
rect 2750 -2422 2770 -2388
rect 2804 -2422 2822 -2388
rect 2750 -2428 2822 -2422
rect 3230 -2388 3302 -2350
rect 3230 -2422 3248 -2388
rect 3282 -2422 3302 -2388
rect 3230 -2428 3302 -2422
rect 3380 -2350 3392 -2344
rect 3426 -2350 3438 -2344
rect 3380 -2388 3438 -2350
rect 3380 -2422 3392 -2388
rect 3426 -2422 3438 -2388
rect 3380 -2428 3438 -2422
rect 3572 -2350 3584 -2344
rect 3618 -2350 3630 -2344
rect 3572 -2388 3630 -2350
rect 3572 -2422 3584 -2388
rect 3618 -2422 3630 -2388
rect 3572 -2428 3630 -2422
rect 3764 -2350 3776 -2344
rect 3810 -2350 3822 -2344
rect 3764 -2388 3822 -2350
rect 3764 -2422 3776 -2388
rect 3810 -2422 3822 -2388
rect 3764 -2428 3822 -2422
rect 3956 -2350 3968 -2344
rect 4002 -2350 4014 -2344
rect 3956 -2388 4014 -2350
rect 3956 -2422 3968 -2388
rect 4002 -2422 4014 -2388
rect 3956 -2428 4014 -2422
rect 4148 -2350 4160 -2344
rect 4194 -2350 4206 -2344
rect 4148 -2388 4206 -2350
rect 4148 -2422 4160 -2388
rect 4194 -2422 4206 -2388
rect 4148 -2428 4206 -2422
rect 4340 -2350 4352 -2344
rect 4386 -2350 4398 -2344
rect 4340 -2388 4398 -2350
rect 4340 -2422 4352 -2388
rect 4386 -2422 4398 -2388
rect 4340 -2428 4398 -2422
rect 4534 -2350 4546 -2344
rect 4580 -2350 4592 -2344
rect 4534 -2388 4592 -2350
rect 4534 -2422 4546 -2388
rect 4580 -2422 4592 -2388
rect 4534 -2428 4592 -2422
rect 4726 -2350 4738 -2344
rect 4772 -2350 4784 -2344
rect 4726 -2388 4784 -2350
rect 4726 -2422 4738 -2388
rect 4772 -2422 4784 -2388
rect 4726 -2428 4784 -2422
rect 4918 -2350 4930 -2344
rect 4964 -2350 4976 -2344
rect 4918 -2388 4976 -2350
rect 4918 -2422 4930 -2388
rect 4964 -2422 4976 -2388
rect 4918 -2428 4976 -2422
rect 5110 -2350 5122 -2344
rect 5156 -2350 5168 -2344
rect 5110 -2388 5168 -2350
rect 5110 -2422 5122 -2388
rect 5156 -2422 5168 -2388
rect 5110 -2428 5168 -2422
rect 5302 -2350 5314 -2344
rect 5348 -2350 5360 -2344
rect 5302 -2388 5360 -2350
rect 5302 -2422 5314 -2388
rect 5348 -2422 5360 -2388
rect 5302 -2428 5360 -2422
rect 5494 -2350 5506 -2344
rect 5540 -2350 5552 -2344
rect 5494 -2388 5552 -2350
rect 5494 -2422 5506 -2388
rect 5540 -2422 5552 -2388
rect 5494 -2428 5552 -2422
rect 5630 -2350 5650 -2316
rect 5684 -2350 5702 -2316
rect 5838 -2344 5854 -2310
rect 5959 -2344 5975 -2310
rect 5630 -2388 5702 -2350
rect 5878 -2350 5890 -2344
rect 5924 -2350 5936 -2344
rect 5878 -2360 5936 -2350
rect 5630 -2422 5650 -2388
rect 5684 -2422 5702 -2388
rect 5630 -2428 5702 -2422
rect 500 -2468 558 -2462
rect 500 -2502 512 -2468
rect 546 -2502 558 -2468
rect 116 -2540 174 -2530
rect 116 -2546 128 -2540
rect 162 -2546 174 -2540
rect 308 -2540 366 -2530
rect 308 -2546 320 -2540
rect 354 -2546 366 -2540
rect 500 -2540 558 -2502
rect 500 -2546 512 -2540
rect 546 -2546 558 -2540
rect 692 -2468 750 -2462
rect 692 -2502 704 -2468
rect 738 -2502 750 -2468
rect 692 -2540 750 -2502
rect 692 -2546 704 -2540
rect 738 -2546 750 -2540
rect 884 -2468 942 -2462
rect 884 -2502 896 -2468
rect 930 -2502 942 -2468
rect 884 -2540 942 -2502
rect 884 -2546 896 -2540
rect 930 -2546 942 -2540
rect 1076 -2468 1134 -2462
rect 1076 -2502 1088 -2468
rect 1122 -2502 1134 -2468
rect 1076 -2540 1134 -2502
rect 1076 -2546 1088 -2540
rect 1122 -2546 1134 -2540
rect 1268 -2468 1326 -2462
rect 1268 -2502 1280 -2468
rect 1314 -2502 1326 -2468
rect 1268 -2540 1326 -2502
rect 1268 -2546 1280 -2540
rect 1314 -2546 1326 -2540
rect 1460 -2468 1518 -2462
rect 1460 -2502 1472 -2468
rect 1506 -2502 1518 -2468
rect 1460 -2540 1518 -2502
rect 1460 -2546 1472 -2540
rect 1506 -2546 1518 -2540
rect 1654 -2468 1712 -2462
rect 1654 -2502 1666 -2468
rect 1700 -2502 1712 -2468
rect 1654 -2540 1712 -2502
rect 1654 -2546 1666 -2540
rect 1700 -2546 1712 -2540
rect 1846 -2468 1904 -2462
rect 1846 -2502 1858 -2468
rect 1892 -2502 1904 -2468
rect 1846 -2540 1904 -2502
rect 1846 -2546 1858 -2540
rect 1892 -2546 1904 -2540
rect 2038 -2468 2096 -2462
rect 2038 -2502 2050 -2468
rect 2084 -2502 2096 -2468
rect 2038 -2540 2096 -2502
rect 2038 -2546 2050 -2540
rect 2084 -2546 2096 -2540
rect 2230 -2468 2288 -2462
rect 2230 -2502 2242 -2468
rect 2276 -2502 2288 -2468
rect 2230 -2540 2288 -2502
rect 2230 -2546 2242 -2540
rect 2276 -2546 2288 -2540
rect 2422 -2468 2480 -2462
rect 2422 -2502 2434 -2468
rect 2468 -2502 2480 -2468
rect 2422 -2540 2480 -2502
rect 2422 -2546 2434 -2540
rect 2468 -2546 2480 -2540
rect 2614 -2468 2672 -2462
rect 2614 -2502 2626 -2468
rect 2660 -2502 2672 -2468
rect 2614 -2540 2672 -2502
rect 3380 -2468 3438 -2462
rect 3380 -2502 3392 -2468
rect 3426 -2502 3438 -2468
rect 2614 -2546 2626 -2540
rect 2660 -2546 2672 -2540
rect 2806 -2540 2864 -2530
rect 2806 -2546 2818 -2540
rect 2852 -2546 2864 -2540
rect 2996 -2540 3056 -2530
rect 2996 -2546 3008 -2540
rect 3044 -2546 3056 -2540
rect 3188 -2540 3246 -2530
rect 3188 -2546 3200 -2540
rect 3234 -2546 3246 -2540
rect 3380 -2540 3438 -2502
rect 3380 -2546 3392 -2540
rect 3426 -2546 3438 -2540
rect 3572 -2468 3630 -2462
rect 3572 -2502 3584 -2468
rect 3618 -2502 3630 -2468
rect 3572 -2540 3630 -2502
rect 3572 -2546 3584 -2540
rect 3618 -2546 3630 -2540
rect 3764 -2468 3822 -2462
rect 3764 -2502 3776 -2468
rect 3810 -2502 3822 -2468
rect 3764 -2540 3822 -2502
rect 3764 -2546 3776 -2540
rect 3810 -2546 3822 -2540
rect 3956 -2468 4014 -2462
rect 3956 -2502 3968 -2468
rect 4002 -2502 4014 -2468
rect 3956 -2540 4014 -2502
rect 3956 -2546 3968 -2540
rect 4002 -2546 4014 -2540
rect 4148 -2468 4206 -2462
rect 4148 -2502 4160 -2468
rect 4194 -2502 4206 -2468
rect 4148 -2540 4206 -2502
rect 4148 -2546 4160 -2540
rect 4194 -2546 4206 -2540
rect 4340 -2468 4398 -2462
rect 4340 -2502 4352 -2468
rect 4386 -2502 4398 -2468
rect 4340 -2540 4398 -2502
rect 4340 -2546 4352 -2540
rect 4386 -2546 4398 -2540
rect 4534 -2468 4592 -2462
rect 4534 -2502 4546 -2468
rect 4580 -2502 4592 -2468
rect 4534 -2540 4592 -2502
rect 4534 -2546 4546 -2540
rect 4580 -2546 4592 -2540
rect 4726 -2468 4784 -2462
rect 4726 -2502 4738 -2468
rect 4772 -2502 4784 -2468
rect 4726 -2540 4784 -2502
rect 4726 -2546 4738 -2540
rect 4772 -2546 4784 -2540
rect 4918 -2468 4976 -2462
rect 4918 -2502 4930 -2468
rect 4964 -2502 4976 -2468
rect 4918 -2540 4976 -2502
rect 4918 -2546 4930 -2540
rect 4964 -2546 4976 -2540
rect 5110 -2468 5168 -2462
rect 5110 -2502 5122 -2468
rect 5156 -2502 5168 -2468
rect 5110 -2540 5168 -2502
rect 5110 -2546 5122 -2540
rect 5156 -2546 5168 -2540
rect 5302 -2468 5360 -2462
rect 5302 -2502 5314 -2468
rect 5348 -2502 5360 -2468
rect 5302 -2540 5360 -2502
rect 5302 -2546 5314 -2540
rect 5348 -2546 5360 -2540
rect 5494 -2468 5552 -2462
rect 5494 -2502 5506 -2468
rect 5540 -2502 5552 -2468
rect 5494 -2540 5552 -2502
rect 5494 -2546 5506 -2540
rect 5540 -2546 5552 -2540
rect 5686 -2540 5744 -2530
rect 5686 -2546 5698 -2540
rect 5732 -2546 5744 -2540
rect 5878 -2540 5936 -2530
rect 5878 -2546 5890 -2540
rect 5924 -2546 5936 -2540
rect 77 -2580 93 -2546
rect 198 -2580 214 -2546
rect 269 -2580 285 -2546
rect 390 -2580 406 -2546
rect 461 -2580 477 -2546
rect 582 -2580 598 -2546
rect 653 -2580 669 -2546
rect 774 -2580 790 -2546
rect 845 -2580 861 -2546
rect 966 -2580 982 -2546
rect 1037 -2580 1053 -2546
rect 1158 -2580 1174 -2546
rect 1229 -2580 1245 -2546
rect 1350 -2580 1366 -2546
rect 1421 -2580 1437 -2546
rect 1542 -2580 1558 -2546
rect 1614 -2580 1630 -2546
rect 1735 -2580 1751 -2546
rect 1806 -2580 1822 -2546
rect 1927 -2580 1943 -2546
rect 1998 -2580 2014 -2546
rect 2119 -2580 2135 -2546
rect 2190 -2580 2206 -2546
rect 2311 -2580 2327 -2546
rect 2382 -2580 2398 -2546
rect 2503 -2580 2519 -2546
rect 2574 -2580 2590 -2546
rect 2695 -2580 2711 -2546
rect 2766 -2580 2782 -2546
rect 2887 -2580 2903 -2546
rect 2957 -2580 2973 -2546
rect 3079 -2580 3095 -2546
rect 3149 -2580 3165 -2546
rect 3270 -2580 3286 -2546
rect 3341 -2580 3357 -2546
rect 3462 -2580 3478 -2546
rect 3533 -2580 3549 -2546
rect 3654 -2580 3670 -2546
rect 3725 -2580 3741 -2546
rect 3846 -2580 3862 -2546
rect 3917 -2580 3933 -2546
rect 4038 -2580 4054 -2546
rect 4109 -2580 4125 -2546
rect 4230 -2580 4246 -2546
rect 4301 -2580 4317 -2546
rect 4422 -2580 4438 -2546
rect 4494 -2580 4510 -2546
rect 4615 -2580 4631 -2546
rect 4686 -2580 4702 -2546
rect 4807 -2580 4823 -2546
rect 4878 -2580 4894 -2546
rect 4999 -2580 5015 -2546
rect 5070 -2580 5086 -2546
rect 5191 -2580 5207 -2546
rect 5262 -2580 5278 -2546
rect 5383 -2580 5399 -2546
rect 5454 -2580 5470 -2546
rect 5575 -2580 5591 -2546
rect 5646 -2580 5662 -2546
rect 5767 -2580 5783 -2546
rect 5838 -2580 5854 -2546
rect 5959 -2580 5975 -2546
rect 33 -2639 67 -2623
rect 33 -3351 67 -3335
rect 129 -2639 163 -2623
rect 129 -3351 163 -3335
rect 225 -2639 259 -2623
rect 225 -3351 259 -3335
rect 321 -2639 355 -2623
rect 321 -3351 355 -3335
rect 417 -2639 451 -2623
rect 417 -3351 451 -3335
rect 513 -2639 547 -2623
rect 513 -3351 547 -3335
rect 609 -2639 643 -2623
rect 609 -3351 643 -3335
rect 705 -2639 739 -2623
rect 705 -3351 739 -3335
rect 801 -2639 835 -2623
rect 801 -3351 835 -3335
rect 897 -2639 931 -2623
rect 897 -3351 931 -3335
rect 993 -2639 1027 -2623
rect 993 -3351 1027 -3335
rect 1089 -2639 1123 -2623
rect 1089 -3351 1123 -3335
rect 1185 -2639 1219 -2623
rect 1185 -3351 1219 -3335
rect 1281 -2639 1315 -2623
rect 1281 -3351 1315 -3335
rect 1377 -2639 1411 -2623
rect 1377 -3351 1411 -3335
rect 1473 -2639 1507 -2623
rect 1473 -3351 1507 -3335
rect 1569 -2639 1603 -2623
rect 1569 -3351 1603 -3335
rect 1665 -2639 1699 -2623
rect 1665 -3351 1699 -3335
rect 1761 -2639 1795 -2623
rect 1761 -3351 1795 -3335
rect 1857 -2639 1891 -2623
rect 1857 -3351 1891 -3335
rect 1953 -2639 1987 -2623
rect 1953 -3351 1987 -3335
rect 2049 -2639 2083 -2623
rect 2049 -3351 2083 -3335
rect 2145 -2639 2179 -2623
rect 2145 -3351 2179 -3335
rect 2241 -2639 2275 -2623
rect 2241 -3351 2275 -3335
rect 2337 -2639 2371 -2623
rect 2337 -3351 2371 -3335
rect 2433 -2639 2467 -2623
rect 2433 -3351 2467 -3335
rect 2529 -2639 2563 -2623
rect 2529 -3351 2563 -3335
rect 2625 -2639 2659 -2623
rect 2625 -3351 2659 -3335
rect 2721 -2639 2755 -2623
rect 2721 -3351 2755 -3335
rect 2817 -2639 2851 -2623
rect 2817 -3351 2851 -3335
rect 2913 -2639 2947 -2623
rect 2913 -3351 2947 -3335
rect 3009 -2639 3043 -2623
rect 3009 -3351 3043 -3335
rect 3105 -2639 3139 -2623
rect 3105 -3351 3139 -3335
rect 3201 -2639 3235 -2623
rect 3201 -3351 3235 -3335
rect 3297 -2639 3331 -2623
rect 3297 -3351 3331 -3335
rect 3393 -2639 3427 -2623
rect 3393 -3351 3427 -3335
rect 3489 -2639 3523 -2623
rect 3489 -3351 3523 -3335
rect 3585 -2639 3619 -2623
rect 3585 -3351 3619 -3335
rect 3681 -2639 3715 -2623
rect 3681 -3351 3715 -3335
rect 3777 -2639 3811 -2623
rect 3777 -3351 3811 -3335
rect 3873 -2639 3907 -2623
rect 3873 -3351 3907 -3335
rect 3969 -2639 4003 -2623
rect 3969 -3351 4003 -3335
rect 4065 -2639 4099 -2623
rect 4065 -3351 4099 -3335
rect 4161 -2639 4195 -2623
rect 4161 -3351 4195 -3335
rect 4257 -2639 4291 -2623
rect 4257 -3351 4291 -3335
rect 4353 -2639 4387 -2623
rect 4353 -3351 4387 -3335
rect 4449 -2639 4483 -2623
rect 4449 -3351 4483 -3335
rect 4545 -2639 4579 -2623
rect 4545 -3351 4579 -3335
rect 4641 -2639 4675 -2623
rect 4641 -3351 4675 -3335
rect 4737 -2639 4771 -2623
rect 4737 -3351 4771 -3335
rect 4833 -2639 4867 -2623
rect 4833 -3351 4867 -3335
rect 4929 -2639 4963 -2623
rect 4929 -3351 4963 -3335
rect 5025 -2639 5059 -2623
rect 5025 -3351 5059 -3335
rect 5121 -2639 5155 -2623
rect 5121 -3351 5155 -3335
rect 5217 -2639 5251 -2623
rect 5217 -3351 5251 -3335
rect 5313 -2639 5347 -2623
rect 5313 -3351 5347 -3335
rect 5409 -2639 5443 -2623
rect 5409 -3351 5443 -3335
rect 5505 -2639 5539 -2623
rect 5505 -3351 5539 -3335
rect 5601 -2639 5635 -2623
rect 5601 -3351 5635 -3335
rect 5697 -2639 5731 -2623
rect 5697 -3351 5731 -3335
rect 5793 -2639 5827 -2623
rect 5793 -3351 5827 -3335
rect 5889 -2639 5923 -2623
rect 5889 -3351 5923 -3335
rect 5985 -2639 6019 -2623
rect 5985 -3351 6019 -3335
rect 26 -3478 126 -3444
rect 5926 -3478 6026 -3444
<< viali >>
rect 126 2024 5926 2058
rect 33 1219 67 1915
rect 129 1219 163 1915
rect 225 1219 259 1915
rect 321 1219 355 1915
rect 417 1219 451 1915
rect 513 1219 547 1915
rect 609 1219 643 1915
rect 705 1219 739 1915
rect 801 1219 835 1915
rect 897 1219 931 1915
rect 993 1219 1027 1915
rect 1089 1219 1123 1915
rect 1185 1219 1219 1915
rect 1281 1219 1315 1915
rect 1377 1219 1411 1915
rect 1473 1219 1507 1915
rect 1569 1219 1603 1915
rect 1665 1219 1699 1915
rect 1761 1219 1795 1915
rect 1857 1219 1891 1915
rect 1953 1219 1987 1915
rect 2049 1219 2083 1915
rect 2145 1219 2179 1915
rect 2241 1219 2275 1915
rect 2337 1219 2371 1915
rect 2433 1219 2467 1915
rect 2529 1219 2563 1915
rect 2625 1219 2659 1915
rect 2721 1219 2755 1915
rect 2817 1219 2851 1915
rect 2913 1219 2947 1915
rect 3009 1219 3043 1915
rect 3105 1219 3139 1915
rect 3201 1219 3235 1915
rect 3297 1219 3331 1915
rect 3393 1219 3427 1915
rect 3489 1219 3523 1915
rect 3585 1219 3619 1915
rect 3681 1219 3715 1915
rect 3777 1219 3811 1915
rect 3873 1219 3907 1915
rect 3969 1219 4003 1915
rect 4065 1219 4099 1915
rect 4161 1219 4195 1915
rect 4257 1219 4291 1915
rect 4353 1219 4387 1915
rect 4449 1219 4483 1915
rect 4545 1219 4579 1915
rect 4641 1219 4675 1915
rect 4737 1219 4771 1915
rect 4833 1219 4867 1915
rect 4929 1219 4963 1915
rect 5025 1219 5059 1915
rect 5121 1219 5155 1915
rect 5217 1219 5251 1915
rect 5313 1219 5347 1915
rect 5409 1219 5443 1915
rect 5505 1219 5539 1915
rect 5601 1219 5635 1915
rect 5697 1219 5731 1915
rect 5793 1219 5827 1915
rect 5889 1219 5923 1915
rect 5985 1219 6019 1915
rect 128 1126 162 1154
rect 320 1126 354 1154
rect 512 1126 546 1154
rect 704 1126 738 1154
rect 896 1126 930 1154
rect 1088 1126 1122 1154
rect 1280 1126 1314 1154
rect 1472 1126 1506 1154
rect 1666 1126 1700 1154
rect 1858 1126 1892 1154
rect 2050 1126 2084 1154
rect 2242 1126 2276 1154
rect 2434 1126 2468 1154
rect 2626 1126 2660 1154
rect 2818 1126 2852 1154
rect 3008 1126 3044 1154
rect 3200 1126 3234 1154
rect 3392 1126 3426 1154
rect 3584 1126 3618 1154
rect 3776 1126 3810 1154
rect 3968 1126 4002 1154
rect 4160 1126 4194 1154
rect 4352 1126 4386 1154
rect 4546 1126 4580 1154
rect 4738 1126 4772 1154
rect 4930 1126 4964 1154
rect 5122 1126 5156 1154
rect 5314 1126 5348 1154
rect 5506 1126 5540 1154
rect 5698 1126 5732 1154
rect 5890 1126 5924 1154
rect 128 1120 162 1126
rect 320 1120 354 1126
rect 512 1120 546 1126
rect 512 1048 546 1082
rect 704 1120 738 1126
rect 704 1048 738 1082
rect 896 1120 930 1126
rect 896 1048 930 1082
rect 1088 1120 1122 1126
rect 1088 1048 1122 1082
rect 1280 1120 1314 1126
rect 1280 1048 1314 1082
rect 1472 1120 1506 1126
rect 1472 1048 1506 1082
rect 1666 1120 1700 1126
rect 1666 1048 1700 1082
rect 1858 1120 1892 1126
rect 1858 1048 1892 1082
rect 2050 1120 2084 1126
rect 2050 1048 2084 1082
rect 2242 1120 2276 1126
rect 2242 1048 2276 1082
rect 2434 1120 2468 1126
rect 2434 1048 2468 1082
rect 2626 1120 2660 1126
rect 2818 1120 2852 1126
rect 3008 1120 3044 1126
rect 3200 1120 3234 1126
rect 3392 1120 3426 1126
rect 2626 1048 2660 1082
rect 3392 1048 3426 1082
rect 3584 1120 3618 1126
rect 3584 1048 3618 1082
rect 3776 1120 3810 1126
rect 3776 1048 3810 1082
rect 3968 1120 4002 1126
rect 3968 1048 4002 1082
rect 4160 1120 4194 1126
rect 4160 1048 4194 1082
rect 4352 1120 4386 1126
rect 4352 1048 4386 1082
rect 4546 1120 4580 1126
rect 4546 1048 4580 1082
rect 4738 1120 4772 1126
rect 4738 1048 4772 1082
rect 4930 1120 4964 1126
rect 4930 1048 4964 1082
rect 5122 1120 5156 1126
rect 5122 1048 5156 1082
rect 5314 1120 5348 1126
rect 5314 1048 5348 1082
rect 5506 1120 5540 1126
rect 5698 1120 5732 1126
rect 5890 1120 5924 1126
rect 5506 1048 5540 1082
rect 368 968 402 1002
rect 128 924 162 930
rect 128 896 162 924
rect 368 896 402 930
rect 512 968 546 1002
rect 512 924 546 930
rect 704 968 738 1002
rect 704 924 738 930
rect 896 968 930 1002
rect 896 924 930 930
rect 1088 968 1122 1002
rect 1088 924 1122 930
rect 1280 968 1314 1002
rect 1280 924 1314 930
rect 1472 968 1506 1002
rect 1472 924 1506 930
rect 1666 968 1700 1002
rect 1666 924 1700 930
rect 1858 968 1892 1002
rect 1858 924 1892 930
rect 2050 968 2084 1002
rect 2050 924 2084 930
rect 2242 968 2276 1002
rect 2242 924 2276 930
rect 2434 968 2468 1002
rect 2434 924 2468 930
rect 2626 968 2660 1002
rect 2626 924 2660 930
rect 2770 968 2804 1002
rect 3248 968 3282 1002
rect 512 896 546 924
rect 704 896 738 924
rect 896 896 930 924
rect 1088 896 1122 924
rect 1280 896 1314 924
rect 1472 896 1506 924
rect 1666 896 1700 924
rect 1858 896 1892 924
rect 2050 896 2084 924
rect 2242 896 2276 924
rect 2434 896 2468 924
rect 2626 896 2660 924
rect 2770 896 2804 930
rect 3008 924 3044 930
rect 3008 896 3044 924
rect 3248 896 3282 930
rect 3392 968 3426 1002
rect 3392 924 3426 930
rect 3584 968 3618 1002
rect 3584 924 3618 930
rect 3776 968 3810 1002
rect 3776 924 3810 930
rect 3968 968 4002 1002
rect 3968 924 4002 930
rect 4160 968 4194 1002
rect 4160 924 4194 930
rect 4352 968 4386 1002
rect 4352 924 4386 930
rect 4546 968 4580 1002
rect 4546 924 4580 930
rect 4738 968 4772 1002
rect 4738 924 4772 930
rect 4930 968 4964 1002
rect 4930 924 4964 930
rect 5122 968 5156 1002
rect 5122 924 5156 930
rect 5314 968 5348 1002
rect 5314 924 5348 930
rect 5506 968 5540 1002
rect 5506 924 5540 930
rect 5650 968 5684 1002
rect 3392 896 3426 924
rect 3584 896 3618 924
rect 3776 896 3810 924
rect 3968 896 4002 924
rect 4160 896 4194 924
rect 4352 896 4386 924
rect 4546 896 4580 924
rect 4738 896 4772 924
rect 4930 896 4964 924
rect 5122 896 5156 924
rect 5314 896 5348 924
rect 5506 896 5540 924
rect 5650 896 5684 930
rect 5890 924 5924 930
rect 5890 896 5924 924
rect 33 464 67 840
rect 129 464 163 840
rect 225 464 259 840
rect 321 464 355 840
rect 417 464 451 840
rect 513 464 547 840
rect 609 464 643 840
rect 705 464 739 840
rect 801 464 835 840
rect 897 464 931 840
rect 993 464 1027 840
rect 1089 464 1123 840
rect 1185 464 1219 840
rect 1281 464 1315 840
rect 1377 464 1411 840
rect 1473 464 1507 840
rect 1569 464 1603 840
rect 1665 464 1699 840
rect 1761 464 1795 840
rect 1857 464 1891 840
rect 1953 464 1987 840
rect 2049 464 2083 840
rect 2145 464 2179 840
rect 2241 464 2275 840
rect 2337 464 2371 840
rect 2433 464 2467 840
rect 2529 464 2563 840
rect 2625 464 2659 840
rect 2721 464 2755 840
rect 2817 464 2851 840
rect 2913 464 2947 840
rect 3009 464 3043 840
rect 3105 464 3139 840
rect 3201 464 3235 840
rect 3297 464 3331 840
rect 3393 464 3427 840
rect 3489 464 3523 840
rect 3585 464 3619 840
rect 3681 464 3715 840
rect 3777 464 3811 840
rect 3873 464 3907 840
rect 3969 464 4003 840
rect 4065 464 4099 840
rect 4161 464 4195 840
rect 4257 464 4291 840
rect 4353 464 4387 840
rect 4449 464 4483 840
rect 4545 464 4579 840
rect 4641 464 4675 840
rect 4737 464 4771 840
rect 4833 464 4867 840
rect 4929 464 4963 840
rect 5025 464 5059 840
rect 5121 464 5155 840
rect 5217 464 5251 840
rect 5313 464 5347 840
rect 5409 464 5443 840
rect 5505 464 5539 840
rect 5601 464 5635 840
rect 5697 464 5731 840
rect 5793 464 5827 840
rect 5889 464 5923 840
rect 5985 464 6019 840
rect 126 322 5926 356
rect 126 -1776 5926 -1742
rect 33 -2260 67 -1884
rect 129 -2260 163 -1884
rect 225 -2260 259 -1884
rect 321 -2260 355 -1884
rect 417 -2260 451 -1884
rect 513 -2260 547 -1884
rect 609 -2260 643 -1884
rect 705 -2260 739 -1884
rect 801 -2260 835 -1884
rect 897 -2260 931 -1884
rect 993 -2260 1027 -1884
rect 1089 -2260 1123 -1884
rect 1185 -2260 1219 -1884
rect 1281 -2260 1315 -1884
rect 1377 -2260 1411 -1884
rect 1473 -2260 1507 -1884
rect 1569 -2260 1603 -1884
rect 1665 -2260 1699 -1884
rect 1761 -2260 1795 -1884
rect 1857 -2260 1891 -1884
rect 1953 -2260 1987 -1884
rect 2049 -2260 2083 -1884
rect 2145 -2260 2179 -1884
rect 2241 -2260 2275 -1884
rect 2337 -2260 2371 -1884
rect 2433 -2260 2467 -1884
rect 2529 -2260 2563 -1884
rect 2625 -2260 2659 -1884
rect 2721 -2260 2755 -1884
rect 2817 -2260 2851 -1884
rect 2913 -2260 2947 -1884
rect 3009 -2260 3043 -1884
rect 3105 -2260 3139 -1884
rect 3201 -2260 3235 -1884
rect 3297 -2260 3331 -1884
rect 3393 -2260 3427 -1884
rect 3489 -2260 3523 -1884
rect 3585 -2260 3619 -1884
rect 3681 -2260 3715 -1884
rect 3777 -2260 3811 -1884
rect 3873 -2260 3907 -1884
rect 3969 -2260 4003 -1884
rect 4065 -2260 4099 -1884
rect 4161 -2260 4195 -1884
rect 4257 -2260 4291 -1884
rect 4353 -2260 4387 -1884
rect 4449 -2260 4483 -1884
rect 4545 -2260 4579 -1884
rect 4641 -2260 4675 -1884
rect 4737 -2260 4771 -1884
rect 4833 -2260 4867 -1884
rect 4929 -2260 4963 -1884
rect 5025 -2260 5059 -1884
rect 5121 -2260 5155 -1884
rect 5217 -2260 5251 -1884
rect 5313 -2260 5347 -1884
rect 5409 -2260 5443 -1884
rect 5505 -2260 5539 -1884
rect 5601 -2260 5635 -1884
rect 5697 -2260 5731 -1884
rect 5793 -2260 5827 -1884
rect 5889 -2260 5923 -1884
rect 5985 -2260 6019 -1884
rect 128 -2344 162 -2316
rect 128 -2350 162 -2344
rect 368 -2350 402 -2316
rect 512 -2344 546 -2316
rect 704 -2344 738 -2316
rect 896 -2344 930 -2316
rect 1088 -2344 1122 -2316
rect 1280 -2344 1314 -2316
rect 1472 -2344 1506 -2316
rect 1666 -2344 1700 -2316
rect 1858 -2344 1892 -2316
rect 2050 -2344 2084 -2316
rect 2242 -2344 2276 -2316
rect 2434 -2344 2468 -2316
rect 2626 -2344 2660 -2316
rect 368 -2422 402 -2388
rect 512 -2350 546 -2344
rect 512 -2422 546 -2388
rect 704 -2350 738 -2344
rect 704 -2422 738 -2388
rect 896 -2350 930 -2344
rect 896 -2422 930 -2388
rect 1088 -2350 1122 -2344
rect 1088 -2422 1122 -2388
rect 1280 -2350 1314 -2344
rect 1280 -2422 1314 -2388
rect 1472 -2350 1506 -2344
rect 1472 -2422 1506 -2388
rect 1666 -2350 1700 -2344
rect 1666 -2422 1700 -2388
rect 1858 -2350 1892 -2344
rect 1858 -2422 1892 -2388
rect 2050 -2350 2084 -2344
rect 2050 -2422 2084 -2388
rect 2242 -2350 2276 -2344
rect 2242 -2422 2276 -2388
rect 2434 -2350 2468 -2344
rect 2434 -2422 2468 -2388
rect 2626 -2350 2660 -2344
rect 2626 -2422 2660 -2388
rect 2770 -2350 2804 -2316
rect 3008 -2344 3044 -2316
rect 3008 -2350 3044 -2344
rect 3248 -2350 3282 -2316
rect 3392 -2344 3426 -2316
rect 3584 -2344 3618 -2316
rect 3776 -2344 3810 -2316
rect 3968 -2344 4002 -2316
rect 4160 -2344 4194 -2316
rect 4352 -2344 4386 -2316
rect 4546 -2344 4580 -2316
rect 4738 -2344 4772 -2316
rect 4930 -2344 4964 -2316
rect 5122 -2344 5156 -2316
rect 5314 -2344 5348 -2316
rect 5506 -2344 5540 -2316
rect 2770 -2422 2804 -2388
rect 3248 -2422 3282 -2388
rect 3392 -2350 3426 -2344
rect 3392 -2422 3426 -2388
rect 3584 -2350 3618 -2344
rect 3584 -2422 3618 -2388
rect 3776 -2350 3810 -2344
rect 3776 -2422 3810 -2388
rect 3968 -2350 4002 -2344
rect 3968 -2422 4002 -2388
rect 4160 -2350 4194 -2344
rect 4160 -2422 4194 -2388
rect 4352 -2350 4386 -2344
rect 4352 -2422 4386 -2388
rect 4546 -2350 4580 -2344
rect 4546 -2422 4580 -2388
rect 4738 -2350 4772 -2344
rect 4738 -2422 4772 -2388
rect 4930 -2350 4964 -2344
rect 4930 -2422 4964 -2388
rect 5122 -2350 5156 -2344
rect 5122 -2422 5156 -2388
rect 5314 -2350 5348 -2344
rect 5314 -2422 5348 -2388
rect 5506 -2350 5540 -2344
rect 5506 -2422 5540 -2388
rect 5650 -2350 5684 -2316
rect 5890 -2344 5924 -2316
rect 5890 -2350 5924 -2344
rect 5650 -2422 5684 -2388
rect 512 -2502 546 -2468
rect 128 -2546 162 -2540
rect 320 -2546 354 -2540
rect 512 -2546 546 -2540
rect 704 -2502 738 -2468
rect 704 -2546 738 -2540
rect 896 -2502 930 -2468
rect 896 -2546 930 -2540
rect 1088 -2502 1122 -2468
rect 1088 -2546 1122 -2540
rect 1280 -2502 1314 -2468
rect 1280 -2546 1314 -2540
rect 1472 -2502 1506 -2468
rect 1472 -2546 1506 -2540
rect 1666 -2502 1700 -2468
rect 1666 -2546 1700 -2540
rect 1858 -2502 1892 -2468
rect 1858 -2546 1892 -2540
rect 2050 -2502 2084 -2468
rect 2050 -2546 2084 -2540
rect 2242 -2502 2276 -2468
rect 2242 -2546 2276 -2540
rect 2434 -2502 2468 -2468
rect 2434 -2546 2468 -2540
rect 2626 -2502 2660 -2468
rect 3392 -2502 3426 -2468
rect 2626 -2546 2660 -2540
rect 2818 -2546 2852 -2540
rect 3008 -2546 3044 -2540
rect 3200 -2546 3234 -2540
rect 3392 -2546 3426 -2540
rect 3584 -2502 3618 -2468
rect 3584 -2546 3618 -2540
rect 3776 -2502 3810 -2468
rect 3776 -2546 3810 -2540
rect 3968 -2502 4002 -2468
rect 3968 -2546 4002 -2540
rect 4160 -2502 4194 -2468
rect 4160 -2546 4194 -2540
rect 4352 -2502 4386 -2468
rect 4352 -2546 4386 -2540
rect 4546 -2502 4580 -2468
rect 4546 -2546 4580 -2540
rect 4738 -2502 4772 -2468
rect 4738 -2546 4772 -2540
rect 4930 -2502 4964 -2468
rect 4930 -2546 4964 -2540
rect 5122 -2502 5156 -2468
rect 5122 -2546 5156 -2540
rect 5314 -2502 5348 -2468
rect 5314 -2546 5348 -2540
rect 5506 -2502 5540 -2468
rect 5506 -2546 5540 -2540
rect 5698 -2546 5732 -2540
rect 5890 -2546 5924 -2540
rect 128 -2574 162 -2546
rect 320 -2574 354 -2546
rect 512 -2574 546 -2546
rect 704 -2574 738 -2546
rect 896 -2574 930 -2546
rect 1088 -2574 1122 -2546
rect 1280 -2574 1314 -2546
rect 1472 -2574 1506 -2546
rect 1666 -2574 1700 -2546
rect 1858 -2574 1892 -2546
rect 2050 -2574 2084 -2546
rect 2242 -2574 2276 -2546
rect 2434 -2574 2468 -2546
rect 2626 -2574 2660 -2546
rect 2818 -2574 2852 -2546
rect 3008 -2574 3044 -2546
rect 3200 -2574 3234 -2546
rect 3392 -2574 3426 -2546
rect 3584 -2574 3618 -2546
rect 3776 -2574 3810 -2546
rect 3968 -2574 4002 -2546
rect 4160 -2574 4194 -2546
rect 4352 -2574 4386 -2546
rect 4546 -2574 4580 -2546
rect 4738 -2574 4772 -2546
rect 4930 -2574 4964 -2546
rect 5122 -2574 5156 -2546
rect 5314 -2574 5348 -2546
rect 5506 -2574 5540 -2546
rect 5698 -2574 5732 -2546
rect 5890 -2574 5924 -2546
rect 33 -3335 67 -2639
rect 129 -3335 163 -2639
rect 225 -3335 259 -2639
rect 321 -3335 355 -2639
rect 417 -3335 451 -2639
rect 513 -3335 547 -2639
rect 609 -3335 643 -2639
rect 705 -3335 739 -2639
rect 801 -3335 835 -2639
rect 897 -3335 931 -2639
rect 993 -3335 1027 -2639
rect 1089 -3335 1123 -2639
rect 1185 -3335 1219 -2639
rect 1281 -3335 1315 -2639
rect 1377 -3335 1411 -2639
rect 1473 -3335 1507 -2639
rect 1569 -3335 1603 -2639
rect 1665 -3335 1699 -2639
rect 1761 -3335 1795 -2639
rect 1857 -3335 1891 -2639
rect 1953 -3335 1987 -2639
rect 2049 -3335 2083 -2639
rect 2145 -3335 2179 -2639
rect 2241 -3335 2275 -2639
rect 2337 -3335 2371 -2639
rect 2433 -3335 2467 -2639
rect 2529 -3335 2563 -2639
rect 2625 -3335 2659 -2639
rect 2721 -3335 2755 -2639
rect 2817 -3335 2851 -2639
rect 2913 -3335 2947 -2639
rect 3009 -3335 3043 -2639
rect 3105 -3335 3139 -2639
rect 3201 -3335 3235 -2639
rect 3297 -3335 3331 -2639
rect 3393 -3335 3427 -2639
rect 3489 -3335 3523 -2639
rect 3585 -3335 3619 -2639
rect 3681 -3335 3715 -2639
rect 3777 -3335 3811 -2639
rect 3873 -3335 3907 -2639
rect 3969 -3335 4003 -2639
rect 4065 -3335 4099 -2639
rect 4161 -3335 4195 -2639
rect 4257 -3335 4291 -2639
rect 4353 -3335 4387 -2639
rect 4449 -3335 4483 -2639
rect 4545 -3335 4579 -2639
rect 4641 -3335 4675 -2639
rect 4737 -3335 4771 -2639
rect 4833 -3335 4867 -2639
rect 4929 -3335 4963 -2639
rect 5025 -3335 5059 -2639
rect 5121 -3335 5155 -2639
rect 5217 -3335 5251 -2639
rect 5313 -3335 5347 -2639
rect 5409 -3335 5443 -2639
rect 5505 -3335 5539 -2639
rect 5601 -3335 5635 -2639
rect 5697 -3335 5731 -2639
rect 5793 -3335 5827 -2639
rect 5889 -3335 5923 -2639
rect 5985 -3335 6019 -2639
rect 126 -3478 5926 -3444
<< metal1 >>
rect 26 2058 6026 2094
rect 26 2024 126 2058
rect 5926 2024 6026 2058
rect 26 1994 6026 2024
rect 26 1915 74 1994
rect 122 1932 170 1994
rect 26 1219 33 1915
rect 67 1219 74 1915
rect 26 1176 74 1219
rect 120 1916 172 1932
rect 120 1204 172 1218
rect 218 1915 266 1994
rect 314 1932 362 1994
rect 218 1219 225 1915
rect 259 1219 266 1915
rect 218 1176 266 1219
rect 312 1916 364 1932
rect 312 1204 364 1218
rect 410 1915 458 1994
rect 410 1219 417 1915
rect 451 1219 458 1915
rect 410 1176 458 1219
rect 504 1916 556 1932
rect 504 1204 556 1218
rect 602 1915 650 1994
rect 602 1219 609 1915
rect 643 1219 650 1915
rect 602 1206 650 1219
rect 696 1916 748 1932
rect 696 1204 748 1218
rect 794 1915 842 1994
rect 794 1219 801 1915
rect 835 1219 842 1915
rect 794 1206 842 1219
rect 888 1916 940 1932
rect 888 1204 940 1218
rect 986 1915 1034 1994
rect 986 1219 993 1915
rect 1027 1219 1034 1915
rect 986 1206 1034 1219
rect 1080 1916 1132 1932
rect 1080 1204 1132 1218
rect 1178 1915 1226 1994
rect 1178 1219 1185 1915
rect 1219 1219 1226 1915
rect 1178 1206 1226 1219
rect 1272 1916 1324 1932
rect 1272 1204 1324 1218
rect 1370 1915 1418 1994
rect 1370 1219 1377 1915
rect 1411 1219 1418 1915
rect 1370 1206 1418 1219
rect 1464 1916 1516 1932
rect 1464 1204 1516 1218
rect 1562 1915 1610 1994
rect 1562 1219 1569 1915
rect 1603 1219 1610 1915
rect 1562 1206 1610 1219
rect 1656 1915 1708 1931
rect 1656 1203 1708 1217
rect 1754 1915 1802 1994
rect 1754 1219 1761 1915
rect 1795 1219 1802 1915
rect 1754 1206 1802 1219
rect 1848 1915 1900 1931
rect 1848 1203 1900 1217
rect 1946 1915 1994 1994
rect 1946 1219 1953 1915
rect 1987 1219 1994 1915
rect 1946 1206 1994 1219
rect 2040 1915 2092 1931
rect 2040 1203 2092 1217
rect 2138 1915 2186 1994
rect 2138 1219 2145 1915
rect 2179 1219 2186 1915
rect 2138 1206 2186 1219
rect 2232 1915 2284 1931
rect 2232 1203 2284 1217
rect 2330 1915 2378 1994
rect 2330 1219 2337 1915
rect 2371 1219 2378 1915
rect 2330 1206 2378 1219
rect 2424 1915 2476 1931
rect 2424 1203 2476 1217
rect 2522 1915 2570 1994
rect 2522 1219 2529 1915
rect 2563 1219 2570 1915
rect 2522 1206 2570 1219
rect 2616 1915 2668 1931
rect 2616 1203 2668 1217
rect 2714 1915 2762 1994
rect 2810 1932 2858 1994
rect 2714 1219 2721 1915
rect 2755 1219 2762 1915
rect 26 1154 458 1176
rect 2714 1176 2762 1219
rect 2808 1916 2860 1932
rect 2808 1204 2860 1218
rect 2906 1915 2954 1994
rect 3002 1932 3050 1994
rect 2906 1219 2913 1915
rect 2947 1219 2954 1915
rect 2906 1176 2954 1219
rect 3000 1916 3052 1932
rect 3000 1204 3052 1218
rect 3098 1915 3146 1994
rect 3194 1932 3242 1994
rect 3098 1219 3105 1915
rect 3139 1219 3146 1915
rect 3098 1176 3146 1219
rect 3192 1916 3244 1932
rect 3192 1204 3244 1218
rect 3290 1915 3338 1994
rect 3290 1219 3297 1915
rect 3331 1219 3338 1915
rect 3290 1176 3338 1219
rect 3384 1916 3436 1932
rect 3384 1204 3436 1218
rect 3482 1915 3530 1994
rect 3482 1219 3489 1915
rect 3523 1219 3530 1915
rect 3482 1206 3530 1219
rect 3576 1916 3628 1932
rect 3576 1204 3628 1218
rect 3674 1915 3722 1994
rect 3674 1219 3681 1915
rect 3715 1219 3722 1915
rect 3674 1206 3722 1219
rect 3768 1916 3820 1932
rect 3768 1204 3820 1218
rect 3866 1915 3914 1994
rect 3866 1219 3873 1915
rect 3907 1219 3914 1915
rect 3866 1206 3914 1219
rect 3960 1916 4012 1932
rect 3960 1204 4012 1218
rect 4058 1915 4106 1994
rect 4058 1219 4065 1915
rect 4099 1219 4106 1915
rect 4058 1206 4106 1219
rect 4152 1916 4204 1932
rect 4152 1204 4204 1218
rect 4250 1915 4298 1994
rect 4250 1219 4257 1915
rect 4291 1219 4298 1915
rect 4250 1206 4298 1219
rect 4344 1916 4396 1932
rect 4344 1204 4396 1218
rect 4442 1915 4490 1994
rect 4442 1219 4449 1915
rect 4483 1219 4490 1915
rect 4442 1206 4490 1219
rect 4536 1915 4588 1931
rect 4536 1203 4588 1217
rect 4634 1915 4682 1994
rect 4634 1219 4641 1915
rect 4675 1219 4682 1915
rect 4634 1206 4682 1219
rect 4728 1915 4780 1931
rect 4728 1203 4780 1217
rect 4826 1915 4874 1994
rect 4826 1219 4833 1915
rect 4867 1219 4874 1915
rect 4826 1206 4874 1219
rect 4920 1915 4972 1931
rect 4920 1203 4972 1217
rect 5018 1915 5066 1994
rect 5018 1219 5025 1915
rect 5059 1219 5066 1915
rect 5018 1206 5066 1219
rect 5112 1915 5164 1931
rect 5112 1203 5164 1217
rect 5210 1915 5258 1994
rect 5210 1219 5217 1915
rect 5251 1219 5258 1915
rect 5210 1206 5258 1219
rect 5304 1915 5356 1931
rect 5304 1203 5356 1217
rect 5402 1915 5450 1994
rect 5402 1219 5409 1915
rect 5443 1219 5450 1915
rect 5402 1206 5450 1219
rect 5496 1915 5548 1931
rect 5496 1203 5548 1217
rect 5594 1915 5642 1994
rect 5690 1932 5738 1994
rect 5594 1219 5601 1915
rect 5635 1219 5642 1915
rect 26 1120 128 1154
rect 162 1120 320 1154
rect 354 1120 458 1154
rect 26 1110 458 1120
rect 500 1154 558 1160
rect 500 1120 512 1154
rect 546 1120 558 1154
rect 500 1082 558 1120
rect 692 1154 750 1160
rect 692 1120 704 1154
rect 738 1120 750 1154
rect 692 1082 750 1120
rect 884 1154 942 1160
rect 884 1120 896 1154
rect 930 1120 942 1154
rect 884 1082 942 1120
rect 1076 1154 1134 1160
rect 1076 1120 1088 1154
rect 1122 1120 1134 1154
rect 1076 1082 1134 1120
rect 1268 1154 1326 1160
rect 1268 1120 1280 1154
rect 1314 1120 1326 1154
rect 1268 1082 1326 1120
rect 1460 1154 1518 1160
rect 1460 1120 1472 1154
rect 1506 1120 1518 1154
rect 1460 1082 1518 1120
rect 500 1048 512 1082
rect 546 1048 704 1082
rect 738 1048 896 1082
rect 930 1048 1088 1082
rect 1122 1048 1134 1082
rect 350 1028 422 1034
rect 350 976 358 1028
rect 410 976 422 1028
rect 350 968 368 976
rect 402 968 422 976
rect 350 948 422 968
rect 26 930 266 940
rect 26 896 128 930
rect 162 896 266 930
rect 26 890 266 896
rect 350 896 358 948
rect 410 896 422 948
rect 350 890 422 896
rect 500 1002 1134 1048
rect 500 968 512 1002
rect 546 968 704 1002
rect 738 968 896 1002
rect 930 968 1088 1002
rect 1122 968 1134 1002
rect 1170 1076 1280 1082
rect 1170 1006 1176 1076
rect 1250 1048 1280 1076
rect 1314 1048 1472 1082
rect 1506 1048 1518 1082
rect 1250 1006 1518 1048
rect 1170 1002 1518 1006
rect 1170 1000 1280 1002
rect 500 930 558 968
rect 500 896 512 930
rect 546 896 558 930
rect 500 890 558 896
rect 692 930 750 968
rect 692 896 704 930
rect 738 896 750 930
rect 692 890 750 896
rect 884 930 942 968
rect 884 896 896 930
rect 930 896 942 930
rect 884 890 942 896
rect 1076 962 1134 968
rect 1268 968 1280 1000
rect 1314 968 1472 1002
rect 1506 968 1518 1002
rect 1076 956 1234 962
rect 1076 930 1170 956
rect 1076 896 1088 930
rect 1122 896 1170 930
rect 1076 894 1170 896
rect 1076 890 1234 894
rect 1268 930 1326 968
rect 1268 896 1280 930
rect 1314 896 1326 930
rect 1268 890 1326 896
rect 1460 930 1518 968
rect 1460 896 1472 930
rect 1506 896 1518 930
rect 1460 890 1518 896
rect 1654 1154 1712 1160
rect 1654 1120 1666 1154
rect 1700 1120 1712 1154
rect 1654 1082 1712 1120
rect 1846 1154 1904 1160
rect 1846 1120 1858 1154
rect 1892 1120 1904 1154
rect 1846 1082 1904 1120
rect 2038 1154 2096 1160
rect 2038 1120 2050 1154
rect 2084 1120 2096 1154
rect 2038 1082 2096 1120
rect 2230 1154 2288 1160
rect 2230 1120 2242 1154
rect 2276 1120 2288 1154
rect 2230 1082 2288 1120
rect 2422 1154 2480 1160
rect 2422 1120 2434 1154
rect 2468 1120 2480 1154
rect 2422 1082 2480 1120
rect 2614 1154 2672 1160
rect 2614 1120 2626 1154
rect 2660 1120 2672 1154
rect 2614 1082 2672 1120
rect 2714 1154 3338 1176
rect 5594 1176 5642 1219
rect 5688 1916 5740 1932
rect 5688 1204 5740 1218
rect 5786 1915 5834 1994
rect 5882 1932 5930 1994
rect 5786 1219 5793 1915
rect 5827 1219 5834 1915
rect 5786 1176 5834 1219
rect 5880 1916 5932 1932
rect 5880 1204 5932 1218
rect 5978 1915 6026 1994
rect 5978 1219 5985 1915
rect 6019 1219 6026 1915
rect 5978 1176 6026 1219
rect 2714 1120 2818 1154
rect 2852 1120 3008 1154
rect 3044 1120 3200 1154
rect 3234 1120 3338 1154
rect 2714 1110 3338 1120
rect 3380 1154 3438 1160
rect 3380 1120 3392 1154
rect 3426 1120 3438 1154
rect 1654 1048 1666 1082
rect 1700 1048 1858 1082
rect 1892 1076 2002 1082
rect 1892 1048 1922 1076
rect 1654 1006 1922 1048
rect 1996 1006 2002 1076
rect 1654 1002 2002 1006
rect 1654 968 1666 1002
rect 1700 968 1858 1002
rect 1892 1000 2002 1002
rect 2038 1048 2050 1082
rect 2084 1048 2242 1082
rect 2276 1048 2434 1082
rect 2468 1048 2626 1082
rect 2660 1048 2672 1082
rect 2038 1002 2672 1048
rect 3380 1082 3438 1120
rect 3572 1154 3630 1160
rect 3572 1120 3584 1154
rect 3618 1120 3630 1154
rect 3572 1082 3630 1120
rect 3764 1154 3822 1160
rect 3764 1120 3776 1154
rect 3810 1120 3822 1154
rect 3764 1082 3822 1120
rect 3956 1154 4014 1160
rect 3956 1120 3968 1154
rect 4002 1120 4014 1154
rect 3956 1082 4014 1120
rect 4148 1154 4206 1160
rect 4148 1120 4160 1154
rect 4194 1120 4206 1154
rect 4148 1082 4206 1120
rect 4340 1154 4398 1160
rect 4340 1120 4352 1154
rect 4386 1120 4398 1154
rect 4340 1082 4398 1120
rect 3380 1048 3392 1082
rect 3426 1048 3584 1082
rect 3618 1048 3776 1082
rect 3810 1048 3968 1082
rect 4002 1048 4014 1082
rect 1892 968 1904 1000
rect 1654 930 1712 968
rect 1654 896 1666 930
rect 1700 896 1712 930
rect 1654 890 1712 896
rect 1846 930 1904 968
rect 2038 968 2050 1002
rect 2084 968 2242 1002
rect 2276 968 2434 1002
rect 2468 968 2626 1002
rect 2660 968 2672 1002
rect 2038 962 2096 968
rect 1846 896 1858 930
rect 1892 896 1904 930
rect 1846 890 1904 896
rect 1938 956 2096 962
rect 2002 930 2096 956
rect 2002 896 2050 930
rect 2084 896 2096 930
rect 2002 894 2096 896
rect 1938 890 2096 894
rect 2230 930 2288 968
rect 2230 896 2242 930
rect 2276 896 2288 930
rect 2230 890 2288 896
rect 2422 930 2480 968
rect 2422 896 2434 930
rect 2468 896 2480 930
rect 2422 890 2480 896
rect 2614 930 2672 968
rect 2614 896 2626 930
rect 2660 896 2672 930
rect 2614 890 2672 896
rect 2750 1028 2822 1034
rect 2750 976 2762 1028
rect 2814 976 2822 1028
rect 2750 968 2770 976
rect 2804 968 2822 976
rect 2750 948 2822 968
rect 2750 896 2762 948
rect 2814 896 2822 948
rect 3230 1028 3302 1034
rect 3230 976 3238 1028
rect 3290 976 3302 1028
rect 3230 968 3248 976
rect 3282 968 3302 976
rect 3230 948 3302 968
rect 2750 890 2822 896
rect 2906 930 3146 940
rect 2906 896 3008 930
rect 3044 896 3146 930
rect 2906 890 3146 896
rect 3230 896 3238 948
rect 3290 896 3302 948
rect 3230 890 3302 896
rect 3380 1002 4014 1048
rect 3380 968 3392 1002
rect 3426 968 3584 1002
rect 3618 968 3776 1002
rect 3810 968 3968 1002
rect 4002 968 4014 1002
rect 4050 1076 4160 1082
rect 4050 1006 4056 1076
rect 4130 1048 4160 1076
rect 4194 1048 4352 1082
rect 4386 1048 4398 1082
rect 4130 1006 4398 1048
rect 4050 1002 4398 1006
rect 4050 1000 4160 1002
rect 3380 930 3438 968
rect 3380 896 3392 930
rect 3426 896 3438 930
rect 3380 890 3438 896
rect 3572 930 3630 968
rect 3572 896 3584 930
rect 3618 896 3630 930
rect 3572 890 3630 896
rect 3764 930 3822 968
rect 3764 896 3776 930
rect 3810 896 3822 930
rect 3764 890 3822 896
rect 3956 962 4014 968
rect 4148 968 4160 1000
rect 4194 968 4352 1002
rect 4386 968 4398 1002
rect 3956 956 4114 962
rect 3956 930 4050 956
rect 3956 896 3968 930
rect 4002 896 4050 930
rect 3956 894 4050 896
rect 3956 890 4114 894
rect 4148 930 4206 968
rect 4148 896 4160 930
rect 4194 896 4206 930
rect 4148 890 4206 896
rect 4340 930 4398 968
rect 4340 896 4352 930
rect 4386 896 4398 930
rect 4340 890 4398 896
rect 4534 1154 4592 1160
rect 4534 1120 4546 1154
rect 4580 1120 4592 1154
rect 4534 1082 4592 1120
rect 4726 1154 4784 1160
rect 4726 1120 4738 1154
rect 4772 1120 4784 1154
rect 4726 1082 4784 1120
rect 4918 1154 4976 1160
rect 4918 1120 4930 1154
rect 4964 1120 4976 1154
rect 4918 1082 4976 1120
rect 5110 1154 5168 1160
rect 5110 1120 5122 1154
rect 5156 1120 5168 1154
rect 5110 1082 5168 1120
rect 5302 1154 5360 1160
rect 5302 1120 5314 1154
rect 5348 1120 5360 1154
rect 5302 1082 5360 1120
rect 5494 1154 5552 1160
rect 5494 1120 5506 1154
rect 5540 1120 5552 1154
rect 5494 1082 5552 1120
rect 5594 1154 6026 1176
rect 5594 1120 5698 1154
rect 5732 1120 5890 1154
rect 5924 1120 6026 1154
rect 5594 1110 6026 1120
rect 4534 1048 4546 1082
rect 4580 1048 4738 1082
rect 4772 1076 4882 1082
rect 4772 1048 4802 1076
rect 4534 1006 4802 1048
rect 4876 1006 4882 1076
rect 4534 1002 4882 1006
rect 4534 968 4546 1002
rect 4580 968 4738 1002
rect 4772 1000 4882 1002
rect 4918 1048 4930 1082
rect 4964 1048 5122 1082
rect 5156 1048 5314 1082
rect 5348 1048 5506 1082
rect 5540 1048 5552 1082
rect 4918 1002 5552 1048
rect 4772 968 4784 1000
rect 4534 930 4592 968
rect 4534 896 4546 930
rect 4580 896 4592 930
rect 4534 890 4592 896
rect 4726 930 4784 968
rect 4918 968 4930 1002
rect 4964 968 5122 1002
rect 5156 968 5314 1002
rect 5348 968 5506 1002
rect 5540 968 5552 1002
rect 4918 962 4976 968
rect 4726 896 4738 930
rect 4772 896 4784 930
rect 4726 890 4784 896
rect 4818 956 4976 962
rect 4882 930 4976 956
rect 4882 896 4930 930
rect 4964 896 4976 930
rect 4882 894 4976 896
rect 4818 890 4976 894
rect 5110 930 5168 968
rect 5110 896 5122 930
rect 5156 896 5168 930
rect 5110 890 5168 896
rect 5302 930 5360 968
rect 5302 896 5314 930
rect 5348 896 5360 930
rect 5302 890 5360 896
rect 5494 930 5552 968
rect 5494 896 5506 930
rect 5540 896 5552 930
rect 5494 890 5552 896
rect 5630 1028 5702 1034
rect 5630 976 5642 1028
rect 5694 976 5702 1028
rect 5630 968 5650 976
rect 5684 968 5702 976
rect 5630 948 5702 968
rect 5630 896 5642 948
rect 5694 896 5702 948
rect 5630 890 5702 896
rect 5786 930 6026 940
rect 5786 896 5890 930
rect 5924 896 6026 930
rect 5786 890 6026 896
rect 26 840 74 890
rect 26 464 33 840
rect 67 464 74 840
rect 26 386 74 464
rect 120 840 172 856
rect 120 448 172 462
rect 218 840 266 890
rect 1170 880 1234 890
rect 1938 888 2038 890
rect 218 464 225 840
rect 259 464 266 840
rect 122 386 170 448
rect 218 386 266 464
rect 312 840 364 856
rect 312 448 364 462
rect 410 840 458 852
rect 410 464 417 840
rect 451 464 458 840
rect 410 386 458 464
rect 504 840 556 856
rect 504 448 556 462
rect 602 840 650 852
rect 602 464 609 840
rect 643 464 650 840
rect 602 386 650 464
rect 696 840 748 856
rect 696 448 748 462
rect 794 840 842 852
rect 794 464 801 840
rect 835 464 842 840
rect 794 386 842 464
rect 888 840 940 856
rect 888 448 940 462
rect 986 840 1034 852
rect 986 464 993 840
rect 1027 464 1034 840
rect 986 386 1034 464
rect 1080 840 1132 856
rect 1080 448 1132 462
rect 1178 840 1226 852
rect 1178 464 1185 840
rect 1219 464 1226 840
rect 1178 386 1226 464
rect 1272 840 1324 856
rect 1272 448 1324 462
rect 1370 840 1418 852
rect 1370 464 1377 840
rect 1411 464 1418 840
rect 1370 386 1418 464
rect 1464 840 1516 856
rect 1464 448 1516 462
rect 1562 840 1610 852
rect 1562 464 1569 840
rect 1603 464 1610 840
rect 1562 386 1610 464
rect 1656 840 1708 856
rect 1656 448 1708 462
rect 1754 840 1802 852
rect 1754 464 1761 840
rect 1795 464 1802 840
rect 1754 386 1802 464
rect 1848 840 1900 856
rect 1848 448 1900 462
rect 1946 840 1994 852
rect 1946 464 1953 840
rect 1987 464 1994 840
rect 1946 386 1994 464
rect 2040 840 2092 856
rect 2040 448 2092 462
rect 2138 840 2186 852
rect 2138 464 2145 840
rect 2179 464 2186 840
rect 2138 386 2186 464
rect 2232 840 2284 856
rect 2232 448 2284 462
rect 2330 840 2378 852
rect 2330 464 2337 840
rect 2371 464 2378 840
rect 2330 386 2378 464
rect 2424 840 2476 856
rect 2424 448 2476 462
rect 2522 840 2570 852
rect 2522 464 2529 840
rect 2563 464 2570 840
rect 2522 386 2570 464
rect 2616 840 2668 856
rect 2616 448 2668 462
rect 2714 840 2762 852
rect 2714 464 2721 840
rect 2755 464 2762 840
rect 2714 386 2762 464
rect 2808 840 2860 856
rect 2808 448 2860 462
rect 2906 840 2954 890
rect 2906 464 2913 840
rect 2947 464 2954 840
rect 2906 386 2954 464
rect 3000 840 3052 856
rect 3000 448 3052 462
rect 3098 840 3146 890
rect 4050 880 4114 890
rect 4818 888 4918 890
rect 3098 464 3105 840
rect 3139 464 3146 840
rect 3002 386 3050 448
rect 3098 386 3146 464
rect 3192 840 3244 856
rect 3192 448 3244 462
rect 3290 840 3338 852
rect 3290 464 3297 840
rect 3331 464 3338 840
rect 3290 386 3338 464
rect 3384 840 3436 856
rect 3384 448 3436 462
rect 3482 840 3530 852
rect 3482 464 3489 840
rect 3523 464 3530 840
rect 3482 386 3530 464
rect 3576 840 3628 856
rect 3576 448 3628 462
rect 3674 840 3722 852
rect 3674 464 3681 840
rect 3715 464 3722 840
rect 3674 386 3722 464
rect 3768 840 3820 856
rect 3768 448 3820 462
rect 3866 840 3914 852
rect 3866 464 3873 840
rect 3907 464 3914 840
rect 3866 386 3914 464
rect 3960 840 4012 856
rect 3960 448 4012 462
rect 4058 840 4106 852
rect 4058 464 4065 840
rect 4099 464 4106 840
rect 4058 386 4106 464
rect 4152 840 4204 856
rect 4152 448 4204 462
rect 4250 840 4298 852
rect 4250 464 4257 840
rect 4291 464 4298 840
rect 4250 386 4298 464
rect 4344 840 4396 856
rect 4344 448 4396 462
rect 4442 840 4490 852
rect 4442 464 4449 840
rect 4483 464 4490 840
rect 4442 386 4490 464
rect 4536 840 4588 856
rect 4536 448 4588 462
rect 4634 840 4682 852
rect 4634 464 4641 840
rect 4675 464 4682 840
rect 4634 386 4682 464
rect 4728 840 4780 856
rect 4728 448 4780 462
rect 4826 840 4874 852
rect 4826 464 4833 840
rect 4867 464 4874 840
rect 4826 386 4874 464
rect 4920 840 4972 856
rect 4920 448 4972 462
rect 5018 840 5066 852
rect 5018 464 5025 840
rect 5059 464 5066 840
rect 5018 386 5066 464
rect 5112 840 5164 856
rect 5112 448 5164 462
rect 5210 840 5258 852
rect 5210 464 5217 840
rect 5251 464 5258 840
rect 5210 386 5258 464
rect 5304 840 5356 856
rect 5304 448 5356 462
rect 5402 840 5450 852
rect 5402 464 5409 840
rect 5443 464 5450 840
rect 5402 386 5450 464
rect 5496 840 5548 856
rect 5496 448 5548 462
rect 5594 840 5642 852
rect 5594 464 5601 840
rect 5635 464 5642 840
rect 5594 386 5642 464
rect 5688 840 5740 856
rect 5688 448 5740 462
rect 5786 840 5834 890
rect 5786 464 5793 840
rect 5827 464 5834 840
rect 5786 386 5834 464
rect 5880 840 5932 856
rect 5880 448 5932 462
rect 5978 840 6026 890
rect 5978 464 5985 840
rect 6019 464 6026 840
rect 5882 386 5930 448
rect 5978 386 6026 464
rect 26 356 6026 386
rect 26 322 126 356
rect 5926 322 6026 356
rect 26 306 6026 322
rect 26 -1742 6026 -1726
rect 26 -1776 126 -1742
rect 5926 -1776 6026 -1742
rect 26 -1806 6026 -1776
rect 26 -1884 74 -1806
rect 122 -1868 170 -1806
rect 26 -2260 33 -1884
rect 67 -2260 74 -1884
rect 26 -2310 74 -2260
rect 120 -1882 172 -1868
rect 120 -2276 172 -2260
rect 218 -1884 266 -1806
rect 218 -2260 225 -1884
rect 259 -2260 266 -1884
rect 218 -2310 266 -2260
rect 312 -1882 364 -1868
rect 312 -2276 364 -2260
rect 410 -1884 458 -1806
rect 410 -2260 417 -1884
rect 451 -2260 458 -1884
rect 410 -2272 458 -2260
rect 504 -1882 556 -1868
rect 504 -2276 556 -2260
rect 602 -1884 650 -1806
rect 602 -2260 609 -1884
rect 643 -2260 650 -1884
rect 602 -2272 650 -2260
rect 696 -1882 748 -1868
rect 696 -2276 748 -2260
rect 794 -1884 842 -1806
rect 794 -2260 801 -1884
rect 835 -2260 842 -1884
rect 794 -2272 842 -2260
rect 888 -1882 940 -1868
rect 888 -2276 940 -2260
rect 986 -1884 1034 -1806
rect 986 -2260 993 -1884
rect 1027 -2260 1034 -1884
rect 986 -2272 1034 -2260
rect 1080 -1882 1132 -1868
rect 1080 -2276 1132 -2260
rect 1178 -1884 1226 -1806
rect 1178 -2260 1185 -1884
rect 1219 -2260 1226 -1884
rect 1178 -2272 1226 -2260
rect 1272 -1882 1324 -1868
rect 1272 -2276 1324 -2260
rect 1370 -1884 1418 -1806
rect 1370 -2260 1377 -1884
rect 1411 -2260 1418 -1884
rect 1370 -2272 1418 -2260
rect 1464 -1882 1516 -1868
rect 1464 -2276 1516 -2260
rect 1562 -1884 1610 -1806
rect 1562 -2260 1569 -1884
rect 1603 -2260 1610 -1884
rect 1562 -2272 1610 -2260
rect 1656 -1882 1708 -1868
rect 1656 -2276 1708 -2260
rect 1754 -1884 1802 -1806
rect 1754 -2260 1761 -1884
rect 1795 -2260 1802 -1884
rect 1754 -2272 1802 -2260
rect 1848 -1882 1900 -1868
rect 1848 -2276 1900 -2260
rect 1946 -1884 1994 -1806
rect 1946 -2260 1953 -1884
rect 1987 -2260 1994 -1884
rect 1946 -2272 1994 -2260
rect 2040 -1882 2092 -1868
rect 2040 -2276 2092 -2260
rect 2138 -1884 2186 -1806
rect 2138 -2260 2145 -1884
rect 2179 -2260 2186 -1884
rect 2138 -2272 2186 -2260
rect 2232 -1882 2284 -1868
rect 2232 -2276 2284 -2260
rect 2330 -1884 2378 -1806
rect 2330 -2260 2337 -1884
rect 2371 -2260 2378 -1884
rect 2330 -2272 2378 -2260
rect 2424 -1882 2476 -1868
rect 2424 -2276 2476 -2260
rect 2522 -1884 2570 -1806
rect 2522 -2260 2529 -1884
rect 2563 -2260 2570 -1884
rect 2522 -2272 2570 -2260
rect 2616 -1882 2668 -1868
rect 2616 -2276 2668 -2260
rect 2714 -1884 2762 -1806
rect 2714 -2260 2721 -1884
rect 2755 -2260 2762 -1884
rect 2714 -2272 2762 -2260
rect 2808 -1882 2860 -1868
rect 2808 -2276 2860 -2260
rect 2906 -1884 2954 -1806
rect 3002 -1868 3050 -1806
rect 2906 -2260 2913 -1884
rect 2947 -2260 2954 -1884
rect 1170 -2310 1234 -2300
rect 1938 -2310 2038 -2308
rect 2906 -2310 2954 -2260
rect 3000 -1882 3052 -1868
rect 3000 -2276 3052 -2260
rect 3098 -1884 3146 -1806
rect 3098 -2260 3105 -1884
rect 3139 -2260 3146 -1884
rect 3098 -2310 3146 -2260
rect 3192 -1882 3244 -1868
rect 3192 -2276 3244 -2260
rect 3290 -1884 3338 -1806
rect 3290 -2260 3297 -1884
rect 3331 -2260 3338 -1884
rect 3290 -2272 3338 -2260
rect 3384 -1882 3436 -1868
rect 3384 -2276 3436 -2260
rect 3482 -1884 3530 -1806
rect 3482 -2260 3489 -1884
rect 3523 -2260 3530 -1884
rect 3482 -2272 3530 -2260
rect 3576 -1882 3628 -1868
rect 3576 -2276 3628 -2260
rect 3674 -1884 3722 -1806
rect 3674 -2260 3681 -1884
rect 3715 -2260 3722 -1884
rect 3674 -2272 3722 -2260
rect 3768 -1882 3820 -1868
rect 3768 -2276 3820 -2260
rect 3866 -1884 3914 -1806
rect 3866 -2260 3873 -1884
rect 3907 -2260 3914 -1884
rect 3866 -2272 3914 -2260
rect 3960 -1882 4012 -1868
rect 3960 -2276 4012 -2260
rect 4058 -1884 4106 -1806
rect 4058 -2260 4065 -1884
rect 4099 -2260 4106 -1884
rect 4058 -2272 4106 -2260
rect 4152 -1882 4204 -1868
rect 4152 -2276 4204 -2260
rect 4250 -1884 4298 -1806
rect 4250 -2260 4257 -1884
rect 4291 -2260 4298 -1884
rect 4250 -2272 4298 -2260
rect 4344 -1882 4396 -1868
rect 4344 -2276 4396 -2260
rect 4442 -1884 4490 -1806
rect 4442 -2260 4449 -1884
rect 4483 -2260 4490 -1884
rect 4442 -2272 4490 -2260
rect 4536 -1882 4588 -1868
rect 4536 -2276 4588 -2260
rect 4634 -1884 4682 -1806
rect 4634 -2260 4641 -1884
rect 4675 -2260 4682 -1884
rect 4634 -2272 4682 -2260
rect 4728 -1882 4780 -1868
rect 4728 -2276 4780 -2260
rect 4826 -1884 4874 -1806
rect 4826 -2260 4833 -1884
rect 4867 -2260 4874 -1884
rect 4826 -2272 4874 -2260
rect 4920 -1882 4972 -1868
rect 4920 -2276 4972 -2260
rect 5018 -1884 5066 -1806
rect 5018 -2260 5025 -1884
rect 5059 -2260 5066 -1884
rect 5018 -2272 5066 -2260
rect 5112 -1882 5164 -1868
rect 5112 -2276 5164 -2260
rect 5210 -1884 5258 -1806
rect 5210 -2260 5217 -1884
rect 5251 -2260 5258 -1884
rect 5210 -2272 5258 -2260
rect 5304 -1882 5356 -1868
rect 5304 -2276 5356 -2260
rect 5402 -1884 5450 -1806
rect 5402 -2260 5409 -1884
rect 5443 -2260 5450 -1884
rect 5402 -2272 5450 -2260
rect 5496 -1882 5548 -1868
rect 5496 -2276 5548 -2260
rect 5594 -1884 5642 -1806
rect 5594 -2260 5601 -1884
rect 5635 -2260 5642 -1884
rect 5594 -2272 5642 -2260
rect 5688 -1882 5740 -1868
rect 5688 -2276 5740 -2260
rect 5786 -1884 5834 -1806
rect 5882 -1868 5930 -1806
rect 5786 -2260 5793 -1884
rect 5827 -2260 5834 -1884
rect 4050 -2310 4114 -2300
rect 4818 -2310 4918 -2308
rect 5786 -2310 5834 -2260
rect 5880 -1882 5932 -1868
rect 5880 -2276 5932 -2260
rect 5978 -1884 6026 -1806
rect 5978 -2260 5985 -1884
rect 6019 -2260 6026 -1884
rect 5978 -2310 6026 -2260
rect 26 -2316 266 -2310
rect 26 -2350 128 -2316
rect 162 -2350 266 -2316
rect 26 -2360 266 -2350
rect 350 -2316 422 -2310
rect 350 -2368 358 -2316
rect 410 -2368 422 -2316
rect 350 -2388 422 -2368
rect 350 -2396 368 -2388
rect 402 -2396 422 -2388
rect 350 -2448 358 -2396
rect 410 -2448 422 -2396
rect 350 -2454 422 -2448
rect 500 -2316 558 -2310
rect 500 -2350 512 -2316
rect 546 -2350 558 -2316
rect 500 -2388 558 -2350
rect 692 -2316 750 -2310
rect 692 -2350 704 -2316
rect 738 -2350 750 -2316
rect 692 -2388 750 -2350
rect 884 -2316 942 -2310
rect 884 -2350 896 -2316
rect 930 -2350 942 -2316
rect 884 -2388 942 -2350
rect 1076 -2314 1234 -2310
rect 1076 -2316 1170 -2314
rect 1076 -2350 1088 -2316
rect 1122 -2350 1170 -2316
rect 1076 -2376 1170 -2350
rect 1076 -2382 1234 -2376
rect 1268 -2316 1326 -2310
rect 1268 -2350 1280 -2316
rect 1314 -2350 1326 -2316
rect 1076 -2388 1134 -2382
rect 500 -2422 512 -2388
rect 546 -2422 704 -2388
rect 738 -2422 896 -2388
rect 930 -2422 1088 -2388
rect 1122 -2422 1134 -2388
rect 1268 -2388 1326 -2350
rect 1460 -2316 1518 -2310
rect 1460 -2350 1472 -2316
rect 1506 -2350 1518 -2316
rect 1460 -2388 1518 -2350
rect 1268 -2420 1280 -2388
rect 500 -2468 1134 -2422
rect 500 -2502 512 -2468
rect 546 -2502 704 -2468
rect 738 -2502 896 -2468
rect 930 -2502 1088 -2468
rect 1122 -2502 1134 -2468
rect 1170 -2422 1280 -2420
rect 1314 -2422 1472 -2388
rect 1506 -2422 1518 -2388
rect 1170 -2426 1518 -2422
rect 1170 -2496 1176 -2426
rect 1250 -2468 1518 -2426
rect 1250 -2496 1280 -2468
rect 1170 -2502 1280 -2496
rect 1314 -2502 1472 -2468
rect 1506 -2502 1518 -2468
rect 26 -2540 458 -2530
rect 26 -2574 128 -2540
rect 162 -2574 320 -2540
rect 354 -2574 458 -2540
rect 26 -2596 458 -2574
rect 500 -2540 558 -2502
rect 500 -2574 512 -2540
rect 546 -2574 558 -2540
rect 500 -2580 558 -2574
rect 692 -2540 750 -2502
rect 692 -2574 704 -2540
rect 738 -2574 750 -2540
rect 692 -2580 750 -2574
rect 884 -2540 942 -2502
rect 884 -2574 896 -2540
rect 930 -2574 942 -2540
rect 884 -2580 942 -2574
rect 1076 -2540 1134 -2502
rect 1076 -2574 1088 -2540
rect 1122 -2574 1134 -2540
rect 1076 -2580 1134 -2574
rect 1268 -2540 1326 -2502
rect 1268 -2574 1280 -2540
rect 1314 -2574 1326 -2540
rect 1268 -2580 1326 -2574
rect 1460 -2540 1518 -2502
rect 1460 -2574 1472 -2540
rect 1506 -2574 1518 -2540
rect 1460 -2580 1518 -2574
rect 1654 -2316 1712 -2310
rect 1654 -2350 1666 -2316
rect 1700 -2350 1712 -2316
rect 1654 -2388 1712 -2350
rect 1846 -2316 1904 -2310
rect 1846 -2350 1858 -2316
rect 1892 -2350 1904 -2316
rect 1846 -2388 1904 -2350
rect 1938 -2314 2096 -2310
rect 2002 -2316 2096 -2314
rect 2002 -2350 2050 -2316
rect 2084 -2350 2096 -2316
rect 2002 -2376 2096 -2350
rect 1938 -2382 2096 -2376
rect 1654 -2422 1666 -2388
rect 1700 -2422 1858 -2388
rect 1892 -2420 1904 -2388
rect 2038 -2388 2096 -2382
rect 2230 -2316 2288 -2310
rect 2230 -2350 2242 -2316
rect 2276 -2350 2288 -2316
rect 2230 -2388 2288 -2350
rect 2422 -2316 2480 -2310
rect 2422 -2350 2434 -2316
rect 2468 -2350 2480 -2316
rect 2422 -2388 2480 -2350
rect 2614 -2316 2672 -2310
rect 2614 -2350 2626 -2316
rect 2660 -2350 2672 -2316
rect 2614 -2388 2672 -2350
rect 1892 -2422 2002 -2420
rect 1654 -2426 2002 -2422
rect 1654 -2468 1922 -2426
rect 1654 -2502 1666 -2468
rect 1700 -2502 1858 -2468
rect 1892 -2496 1922 -2468
rect 1996 -2496 2002 -2426
rect 1892 -2502 2002 -2496
rect 2038 -2422 2050 -2388
rect 2084 -2422 2242 -2388
rect 2276 -2422 2434 -2388
rect 2468 -2422 2626 -2388
rect 2660 -2422 2672 -2388
rect 2038 -2468 2672 -2422
rect 2750 -2316 2822 -2310
rect 2750 -2368 2762 -2316
rect 2814 -2368 2822 -2316
rect 2906 -2316 3146 -2310
rect 2906 -2350 3008 -2316
rect 3044 -2350 3146 -2316
rect 2906 -2360 3146 -2350
rect 3230 -2316 3302 -2310
rect 2750 -2388 2822 -2368
rect 2750 -2396 2770 -2388
rect 2804 -2396 2822 -2388
rect 2750 -2448 2762 -2396
rect 2814 -2448 2822 -2396
rect 2750 -2454 2822 -2448
rect 3230 -2368 3238 -2316
rect 3290 -2368 3302 -2316
rect 3230 -2388 3302 -2368
rect 3230 -2396 3248 -2388
rect 3282 -2396 3302 -2388
rect 3230 -2448 3238 -2396
rect 3290 -2448 3302 -2396
rect 3230 -2454 3302 -2448
rect 3380 -2316 3438 -2310
rect 3380 -2350 3392 -2316
rect 3426 -2350 3438 -2316
rect 3380 -2388 3438 -2350
rect 3572 -2316 3630 -2310
rect 3572 -2350 3584 -2316
rect 3618 -2350 3630 -2316
rect 3572 -2388 3630 -2350
rect 3764 -2316 3822 -2310
rect 3764 -2350 3776 -2316
rect 3810 -2350 3822 -2316
rect 3764 -2388 3822 -2350
rect 3956 -2314 4114 -2310
rect 3956 -2316 4050 -2314
rect 3956 -2350 3968 -2316
rect 4002 -2350 4050 -2316
rect 3956 -2376 4050 -2350
rect 3956 -2382 4114 -2376
rect 4148 -2316 4206 -2310
rect 4148 -2350 4160 -2316
rect 4194 -2350 4206 -2316
rect 3956 -2388 4014 -2382
rect 3380 -2422 3392 -2388
rect 3426 -2422 3584 -2388
rect 3618 -2422 3776 -2388
rect 3810 -2422 3968 -2388
rect 4002 -2422 4014 -2388
rect 4148 -2388 4206 -2350
rect 4340 -2316 4398 -2310
rect 4340 -2350 4352 -2316
rect 4386 -2350 4398 -2316
rect 4340 -2388 4398 -2350
rect 4148 -2420 4160 -2388
rect 2038 -2502 2050 -2468
rect 2084 -2502 2242 -2468
rect 2276 -2502 2434 -2468
rect 2468 -2502 2626 -2468
rect 2660 -2502 2672 -2468
rect 1654 -2540 1712 -2502
rect 1654 -2574 1666 -2540
rect 1700 -2574 1712 -2540
rect 1654 -2580 1712 -2574
rect 1846 -2540 1904 -2502
rect 1846 -2574 1858 -2540
rect 1892 -2574 1904 -2540
rect 1846 -2580 1904 -2574
rect 2038 -2540 2096 -2502
rect 2038 -2574 2050 -2540
rect 2084 -2574 2096 -2540
rect 2038 -2580 2096 -2574
rect 2230 -2540 2288 -2502
rect 2230 -2574 2242 -2540
rect 2276 -2574 2288 -2540
rect 2230 -2580 2288 -2574
rect 2422 -2540 2480 -2502
rect 2422 -2574 2434 -2540
rect 2468 -2574 2480 -2540
rect 2422 -2580 2480 -2574
rect 2614 -2540 2672 -2502
rect 3380 -2468 4014 -2422
rect 3380 -2502 3392 -2468
rect 3426 -2502 3584 -2468
rect 3618 -2502 3776 -2468
rect 3810 -2502 3968 -2468
rect 4002 -2502 4014 -2468
rect 4050 -2422 4160 -2420
rect 4194 -2422 4352 -2388
rect 4386 -2422 4398 -2388
rect 4050 -2426 4398 -2422
rect 4050 -2496 4056 -2426
rect 4130 -2468 4398 -2426
rect 4130 -2496 4160 -2468
rect 4050 -2502 4160 -2496
rect 4194 -2502 4352 -2468
rect 4386 -2502 4398 -2468
rect 2614 -2574 2626 -2540
rect 2660 -2574 2672 -2540
rect 2614 -2580 2672 -2574
rect 2714 -2540 3338 -2530
rect 2714 -2574 2818 -2540
rect 2852 -2574 3008 -2540
rect 3044 -2574 3200 -2540
rect 3234 -2574 3338 -2540
rect 26 -2639 74 -2596
rect 26 -3335 33 -2639
rect 67 -3335 74 -2639
rect 26 -3414 74 -3335
rect 120 -2638 172 -2624
rect 120 -3352 172 -3336
rect 218 -2639 266 -2596
rect 218 -3335 225 -2639
rect 259 -3335 266 -2639
rect 122 -3414 170 -3352
rect 218 -3414 266 -3335
rect 312 -2638 364 -2624
rect 312 -3352 364 -3336
rect 410 -2639 458 -2596
rect 2714 -2596 3338 -2574
rect 3380 -2540 3438 -2502
rect 3380 -2574 3392 -2540
rect 3426 -2574 3438 -2540
rect 3380 -2580 3438 -2574
rect 3572 -2540 3630 -2502
rect 3572 -2574 3584 -2540
rect 3618 -2574 3630 -2540
rect 3572 -2580 3630 -2574
rect 3764 -2540 3822 -2502
rect 3764 -2574 3776 -2540
rect 3810 -2574 3822 -2540
rect 3764 -2580 3822 -2574
rect 3956 -2540 4014 -2502
rect 3956 -2574 3968 -2540
rect 4002 -2574 4014 -2540
rect 3956 -2580 4014 -2574
rect 4148 -2540 4206 -2502
rect 4148 -2574 4160 -2540
rect 4194 -2574 4206 -2540
rect 4148 -2580 4206 -2574
rect 4340 -2540 4398 -2502
rect 4340 -2574 4352 -2540
rect 4386 -2574 4398 -2540
rect 4340 -2580 4398 -2574
rect 4534 -2316 4592 -2310
rect 4534 -2350 4546 -2316
rect 4580 -2350 4592 -2316
rect 4534 -2388 4592 -2350
rect 4726 -2316 4784 -2310
rect 4726 -2350 4738 -2316
rect 4772 -2350 4784 -2316
rect 4726 -2388 4784 -2350
rect 4818 -2314 4976 -2310
rect 4882 -2316 4976 -2314
rect 4882 -2350 4930 -2316
rect 4964 -2350 4976 -2316
rect 4882 -2376 4976 -2350
rect 4818 -2382 4976 -2376
rect 4534 -2422 4546 -2388
rect 4580 -2422 4738 -2388
rect 4772 -2420 4784 -2388
rect 4918 -2388 4976 -2382
rect 5110 -2316 5168 -2310
rect 5110 -2350 5122 -2316
rect 5156 -2350 5168 -2316
rect 5110 -2388 5168 -2350
rect 5302 -2316 5360 -2310
rect 5302 -2350 5314 -2316
rect 5348 -2350 5360 -2316
rect 5302 -2388 5360 -2350
rect 5494 -2316 5552 -2310
rect 5494 -2350 5506 -2316
rect 5540 -2350 5552 -2316
rect 5494 -2388 5552 -2350
rect 4772 -2422 4882 -2420
rect 4534 -2426 4882 -2422
rect 4534 -2468 4802 -2426
rect 4534 -2502 4546 -2468
rect 4580 -2502 4738 -2468
rect 4772 -2496 4802 -2468
rect 4876 -2496 4882 -2426
rect 4772 -2502 4882 -2496
rect 4918 -2422 4930 -2388
rect 4964 -2422 5122 -2388
rect 5156 -2422 5314 -2388
rect 5348 -2422 5506 -2388
rect 5540 -2422 5552 -2388
rect 4918 -2468 5552 -2422
rect 5630 -2316 5702 -2310
rect 5630 -2368 5642 -2316
rect 5694 -2368 5702 -2316
rect 5786 -2316 6026 -2310
rect 5786 -2350 5890 -2316
rect 5924 -2350 6026 -2316
rect 5786 -2360 6026 -2350
rect 5630 -2388 5702 -2368
rect 5630 -2396 5650 -2388
rect 5684 -2396 5702 -2388
rect 5630 -2448 5642 -2396
rect 5694 -2448 5702 -2396
rect 5630 -2454 5702 -2448
rect 4918 -2502 4930 -2468
rect 4964 -2502 5122 -2468
rect 5156 -2502 5314 -2468
rect 5348 -2502 5506 -2468
rect 5540 -2502 5552 -2468
rect 4534 -2540 4592 -2502
rect 4534 -2574 4546 -2540
rect 4580 -2574 4592 -2540
rect 4534 -2580 4592 -2574
rect 4726 -2540 4784 -2502
rect 4726 -2574 4738 -2540
rect 4772 -2574 4784 -2540
rect 4726 -2580 4784 -2574
rect 4918 -2540 4976 -2502
rect 4918 -2574 4930 -2540
rect 4964 -2574 4976 -2540
rect 4918 -2580 4976 -2574
rect 5110 -2540 5168 -2502
rect 5110 -2574 5122 -2540
rect 5156 -2574 5168 -2540
rect 5110 -2580 5168 -2574
rect 5302 -2540 5360 -2502
rect 5302 -2574 5314 -2540
rect 5348 -2574 5360 -2540
rect 5302 -2580 5360 -2574
rect 5494 -2540 5552 -2502
rect 5494 -2574 5506 -2540
rect 5540 -2574 5552 -2540
rect 5494 -2580 5552 -2574
rect 5594 -2540 6026 -2530
rect 5594 -2574 5698 -2540
rect 5732 -2574 5890 -2540
rect 5924 -2574 6026 -2540
rect 410 -3335 417 -2639
rect 451 -3335 458 -2639
rect 314 -3414 362 -3352
rect 410 -3414 458 -3335
rect 504 -2638 556 -2624
rect 504 -3352 556 -3336
rect 602 -2639 650 -2626
rect 602 -3335 609 -2639
rect 643 -3335 650 -2639
rect 602 -3414 650 -3335
rect 696 -2638 748 -2624
rect 696 -3352 748 -3336
rect 794 -2639 842 -2626
rect 794 -3335 801 -2639
rect 835 -3335 842 -2639
rect 794 -3414 842 -3335
rect 888 -2638 940 -2624
rect 888 -3352 940 -3336
rect 986 -2639 1034 -2626
rect 986 -3335 993 -2639
rect 1027 -3335 1034 -2639
rect 986 -3414 1034 -3335
rect 1080 -2638 1132 -2624
rect 1080 -3352 1132 -3336
rect 1178 -2639 1226 -2626
rect 1178 -3335 1185 -2639
rect 1219 -3335 1226 -2639
rect 1178 -3414 1226 -3335
rect 1272 -2638 1324 -2624
rect 1272 -3352 1324 -3336
rect 1370 -2639 1418 -2626
rect 1370 -3335 1377 -2639
rect 1411 -3335 1418 -2639
rect 1370 -3414 1418 -3335
rect 1464 -2638 1516 -2624
rect 1464 -3352 1516 -3336
rect 1562 -2639 1610 -2626
rect 1562 -3335 1569 -2639
rect 1603 -3335 1610 -2639
rect 1562 -3414 1610 -3335
rect 1656 -2637 1708 -2623
rect 1656 -3351 1708 -3335
rect 1754 -2639 1802 -2626
rect 1754 -3335 1761 -2639
rect 1795 -3335 1802 -2639
rect 1754 -3414 1802 -3335
rect 1848 -2637 1900 -2623
rect 1848 -3351 1900 -3335
rect 1946 -2639 1994 -2626
rect 1946 -3335 1953 -2639
rect 1987 -3335 1994 -2639
rect 1946 -3414 1994 -3335
rect 2040 -2637 2092 -2623
rect 2040 -3351 2092 -3335
rect 2138 -2639 2186 -2626
rect 2138 -3335 2145 -2639
rect 2179 -3335 2186 -2639
rect 2138 -3414 2186 -3335
rect 2232 -2637 2284 -2623
rect 2232 -3351 2284 -3335
rect 2330 -2639 2378 -2626
rect 2330 -3335 2337 -2639
rect 2371 -3335 2378 -2639
rect 2330 -3414 2378 -3335
rect 2424 -2637 2476 -2623
rect 2424 -3351 2476 -3335
rect 2522 -2639 2570 -2626
rect 2522 -3335 2529 -2639
rect 2563 -3335 2570 -2639
rect 2522 -3414 2570 -3335
rect 2616 -2637 2668 -2623
rect 2616 -3351 2668 -3335
rect 2714 -2639 2762 -2596
rect 2714 -3335 2721 -2639
rect 2755 -3335 2762 -2639
rect 2714 -3414 2762 -3335
rect 2808 -2638 2860 -2624
rect 2808 -3352 2860 -3336
rect 2906 -2639 2954 -2596
rect 2906 -3335 2913 -2639
rect 2947 -3335 2954 -2639
rect 2810 -3414 2858 -3352
rect 2906 -3414 2954 -3335
rect 3000 -2638 3052 -2624
rect 3000 -3352 3052 -3336
rect 3098 -2639 3146 -2596
rect 3098 -3335 3105 -2639
rect 3139 -3335 3146 -2639
rect 3002 -3414 3050 -3352
rect 3098 -3414 3146 -3335
rect 3192 -2638 3244 -2624
rect 3192 -3352 3244 -3336
rect 3290 -2639 3338 -2596
rect 5594 -2596 6026 -2574
rect 3290 -3335 3297 -2639
rect 3331 -3335 3338 -2639
rect 3194 -3414 3242 -3352
rect 3290 -3414 3338 -3335
rect 3384 -2638 3436 -2624
rect 3384 -3352 3436 -3336
rect 3482 -2639 3530 -2626
rect 3482 -3335 3489 -2639
rect 3523 -3335 3530 -2639
rect 3482 -3414 3530 -3335
rect 3576 -2638 3628 -2624
rect 3576 -3352 3628 -3336
rect 3674 -2639 3722 -2626
rect 3674 -3335 3681 -2639
rect 3715 -3335 3722 -2639
rect 3674 -3414 3722 -3335
rect 3768 -2638 3820 -2624
rect 3768 -3352 3820 -3336
rect 3866 -2639 3914 -2626
rect 3866 -3335 3873 -2639
rect 3907 -3335 3914 -2639
rect 3866 -3414 3914 -3335
rect 3960 -2638 4012 -2624
rect 3960 -3352 4012 -3336
rect 4058 -2639 4106 -2626
rect 4058 -3335 4065 -2639
rect 4099 -3335 4106 -2639
rect 4058 -3414 4106 -3335
rect 4152 -2638 4204 -2624
rect 4152 -3352 4204 -3336
rect 4250 -2639 4298 -2626
rect 4250 -3335 4257 -2639
rect 4291 -3335 4298 -2639
rect 4250 -3414 4298 -3335
rect 4344 -2638 4396 -2624
rect 4344 -3352 4396 -3336
rect 4442 -2639 4490 -2626
rect 4442 -3335 4449 -2639
rect 4483 -3335 4490 -2639
rect 4442 -3414 4490 -3335
rect 4536 -2637 4588 -2623
rect 4536 -3351 4588 -3335
rect 4634 -2639 4682 -2626
rect 4634 -3335 4641 -2639
rect 4675 -3335 4682 -2639
rect 4634 -3414 4682 -3335
rect 4728 -2637 4780 -2623
rect 4728 -3351 4780 -3335
rect 4826 -2639 4874 -2626
rect 4826 -3335 4833 -2639
rect 4867 -3335 4874 -2639
rect 4826 -3414 4874 -3335
rect 4920 -2637 4972 -2623
rect 4920 -3351 4972 -3335
rect 5018 -2639 5066 -2626
rect 5018 -3335 5025 -2639
rect 5059 -3335 5066 -2639
rect 5018 -3414 5066 -3335
rect 5112 -2637 5164 -2623
rect 5112 -3351 5164 -3335
rect 5210 -2639 5258 -2626
rect 5210 -3335 5217 -2639
rect 5251 -3335 5258 -2639
rect 5210 -3414 5258 -3335
rect 5304 -2637 5356 -2623
rect 5304 -3351 5356 -3335
rect 5402 -2639 5450 -2626
rect 5402 -3335 5409 -2639
rect 5443 -3335 5450 -2639
rect 5402 -3414 5450 -3335
rect 5496 -2637 5548 -2623
rect 5496 -3351 5548 -3335
rect 5594 -2639 5642 -2596
rect 5594 -3335 5601 -2639
rect 5635 -3335 5642 -2639
rect 5594 -3414 5642 -3335
rect 5688 -2638 5740 -2624
rect 5688 -3352 5740 -3336
rect 5786 -2639 5834 -2596
rect 5786 -3335 5793 -2639
rect 5827 -3335 5834 -2639
rect 5690 -3414 5738 -3352
rect 5786 -3414 5834 -3335
rect 5880 -2638 5932 -2624
rect 5880 -3352 5932 -3336
rect 5978 -2639 6026 -2596
rect 5978 -3335 5985 -2639
rect 6019 -3335 6026 -2639
rect 5882 -3414 5930 -3352
rect 5978 -3414 6026 -3335
rect 26 -3444 6026 -3414
rect 26 -3478 126 -3444
rect 5926 -3478 6026 -3444
rect 26 -3514 6026 -3478
<< via1 >>
rect 120 1915 172 1916
rect 120 1219 129 1915
rect 129 1219 163 1915
rect 163 1219 172 1915
rect 120 1218 172 1219
rect 312 1915 364 1916
rect 312 1219 321 1915
rect 321 1219 355 1915
rect 355 1219 364 1915
rect 312 1218 364 1219
rect 504 1915 556 1916
rect 504 1219 513 1915
rect 513 1219 547 1915
rect 547 1219 556 1915
rect 504 1218 556 1219
rect 696 1915 748 1916
rect 696 1219 705 1915
rect 705 1219 739 1915
rect 739 1219 748 1915
rect 696 1218 748 1219
rect 888 1915 940 1916
rect 888 1219 897 1915
rect 897 1219 931 1915
rect 931 1219 940 1915
rect 888 1218 940 1219
rect 1080 1915 1132 1916
rect 1080 1219 1089 1915
rect 1089 1219 1123 1915
rect 1123 1219 1132 1915
rect 1080 1218 1132 1219
rect 1272 1915 1324 1916
rect 1272 1219 1281 1915
rect 1281 1219 1315 1915
rect 1315 1219 1324 1915
rect 1272 1218 1324 1219
rect 1464 1915 1516 1916
rect 1464 1219 1473 1915
rect 1473 1219 1507 1915
rect 1507 1219 1516 1915
rect 1464 1218 1516 1219
rect 1656 1219 1665 1915
rect 1665 1219 1699 1915
rect 1699 1219 1708 1915
rect 1656 1217 1708 1219
rect 1848 1219 1857 1915
rect 1857 1219 1891 1915
rect 1891 1219 1900 1915
rect 1848 1217 1900 1219
rect 2040 1219 2049 1915
rect 2049 1219 2083 1915
rect 2083 1219 2092 1915
rect 2040 1217 2092 1219
rect 2232 1219 2241 1915
rect 2241 1219 2275 1915
rect 2275 1219 2284 1915
rect 2232 1217 2284 1219
rect 2424 1219 2433 1915
rect 2433 1219 2467 1915
rect 2467 1219 2476 1915
rect 2424 1217 2476 1219
rect 2616 1219 2625 1915
rect 2625 1219 2659 1915
rect 2659 1219 2668 1915
rect 2616 1217 2668 1219
rect 2808 1915 2860 1916
rect 2808 1219 2817 1915
rect 2817 1219 2851 1915
rect 2851 1219 2860 1915
rect 2808 1218 2860 1219
rect 3000 1915 3052 1916
rect 3000 1219 3009 1915
rect 3009 1219 3043 1915
rect 3043 1219 3052 1915
rect 3000 1218 3052 1219
rect 3192 1915 3244 1916
rect 3192 1219 3201 1915
rect 3201 1219 3235 1915
rect 3235 1219 3244 1915
rect 3192 1218 3244 1219
rect 3384 1915 3436 1916
rect 3384 1219 3393 1915
rect 3393 1219 3427 1915
rect 3427 1219 3436 1915
rect 3384 1218 3436 1219
rect 3576 1915 3628 1916
rect 3576 1219 3585 1915
rect 3585 1219 3619 1915
rect 3619 1219 3628 1915
rect 3576 1218 3628 1219
rect 3768 1915 3820 1916
rect 3768 1219 3777 1915
rect 3777 1219 3811 1915
rect 3811 1219 3820 1915
rect 3768 1218 3820 1219
rect 3960 1915 4012 1916
rect 3960 1219 3969 1915
rect 3969 1219 4003 1915
rect 4003 1219 4012 1915
rect 3960 1218 4012 1219
rect 4152 1915 4204 1916
rect 4152 1219 4161 1915
rect 4161 1219 4195 1915
rect 4195 1219 4204 1915
rect 4152 1218 4204 1219
rect 4344 1915 4396 1916
rect 4344 1219 4353 1915
rect 4353 1219 4387 1915
rect 4387 1219 4396 1915
rect 4344 1218 4396 1219
rect 4536 1219 4545 1915
rect 4545 1219 4579 1915
rect 4579 1219 4588 1915
rect 4536 1217 4588 1219
rect 4728 1219 4737 1915
rect 4737 1219 4771 1915
rect 4771 1219 4780 1915
rect 4728 1217 4780 1219
rect 4920 1219 4929 1915
rect 4929 1219 4963 1915
rect 4963 1219 4972 1915
rect 4920 1217 4972 1219
rect 5112 1219 5121 1915
rect 5121 1219 5155 1915
rect 5155 1219 5164 1915
rect 5112 1217 5164 1219
rect 5304 1219 5313 1915
rect 5313 1219 5347 1915
rect 5347 1219 5356 1915
rect 5304 1217 5356 1219
rect 5496 1219 5505 1915
rect 5505 1219 5539 1915
rect 5539 1219 5548 1915
rect 5496 1217 5548 1219
rect 358 1002 410 1028
rect 358 976 368 1002
rect 368 976 402 1002
rect 402 976 410 1002
rect 358 930 410 948
rect 358 896 368 930
rect 368 896 402 930
rect 402 896 410 930
rect 1176 1006 1250 1076
rect 1170 894 1234 956
rect 5688 1915 5740 1916
rect 5688 1219 5697 1915
rect 5697 1219 5731 1915
rect 5731 1219 5740 1915
rect 5688 1218 5740 1219
rect 5880 1915 5932 1916
rect 5880 1219 5889 1915
rect 5889 1219 5923 1915
rect 5923 1219 5932 1915
rect 5880 1218 5932 1219
rect 1922 1006 1996 1076
rect 1938 894 2002 956
rect 2762 1002 2814 1028
rect 2762 976 2770 1002
rect 2770 976 2804 1002
rect 2804 976 2814 1002
rect 2762 930 2814 948
rect 2762 896 2770 930
rect 2770 896 2804 930
rect 2804 896 2814 930
rect 3238 1002 3290 1028
rect 3238 976 3248 1002
rect 3248 976 3282 1002
rect 3282 976 3290 1002
rect 3238 930 3290 948
rect 3238 896 3248 930
rect 3248 896 3282 930
rect 3282 896 3290 930
rect 4056 1006 4130 1076
rect 4050 894 4114 956
rect 4802 1006 4876 1076
rect 4818 894 4882 956
rect 5642 1002 5694 1028
rect 5642 976 5650 1002
rect 5650 976 5684 1002
rect 5684 976 5694 1002
rect 5642 930 5694 948
rect 5642 896 5650 930
rect 5650 896 5684 930
rect 5684 896 5694 930
rect 120 464 129 840
rect 129 464 163 840
rect 163 464 172 840
rect 120 462 172 464
rect 312 464 321 840
rect 321 464 355 840
rect 355 464 364 840
rect 312 462 364 464
rect 504 464 513 840
rect 513 464 547 840
rect 547 464 556 840
rect 504 462 556 464
rect 696 464 705 840
rect 705 464 739 840
rect 739 464 748 840
rect 696 462 748 464
rect 888 464 897 840
rect 897 464 931 840
rect 931 464 940 840
rect 888 462 940 464
rect 1080 464 1089 840
rect 1089 464 1123 840
rect 1123 464 1132 840
rect 1080 462 1132 464
rect 1272 464 1281 840
rect 1281 464 1315 840
rect 1315 464 1324 840
rect 1272 462 1324 464
rect 1464 464 1473 840
rect 1473 464 1507 840
rect 1507 464 1516 840
rect 1464 462 1516 464
rect 1656 464 1665 840
rect 1665 464 1699 840
rect 1699 464 1708 840
rect 1656 462 1708 464
rect 1848 464 1857 840
rect 1857 464 1891 840
rect 1891 464 1900 840
rect 1848 462 1900 464
rect 2040 464 2049 840
rect 2049 464 2083 840
rect 2083 464 2092 840
rect 2040 462 2092 464
rect 2232 464 2241 840
rect 2241 464 2275 840
rect 2275 464 2284 840
rect 2232 462 2284 464
rect 2424 464 2433 840
rect 2433 464 2467 840
rect 2467 464 2476 840
rect 2424 462 2476 464
rect 2616 464 2625 840
rect 2625 464 2659 840
rect 2659 464 2668 840
rect 2616 462 2668 464
rect 2808 464 2817 840
rect 2817 464 2851 840
rect 2851 464 2860 840
rect 2808 462 2860 464
rect 3000 464 3009 840
rect 3009 464 3043 840
rect 3043 464 3052 840
rect 3000 462 3052 464
rect 3192 464 3201 840
rect 3201 464 3235 840
rect 3235 464 3244 840
rect 3192 462 3244 464
rect 3384 464 3393 840
rect 3393 464 3427 840
rect 3427 464 3436 840
rect 3384 462 3436 464
rect 3576 464 3585 840
rect 3585 464 3619 840
rect 3619 464 3628 840
rect 3576 462 3628 464
rect 3768 464 3777 840
rect 3777 464 3811 840
rect 3811 464 3820 840
rect 3768 462 3820 464
rect 3960 464 3969 840
rect 3969 464 4003 840
rect 4003 464 4012 840
rect 3960 462 4012 464
rect 4152 464 4161 840
rect 4161 464 4195 840
rect 4195 464 4204 840
rect 4152 462 4204 464
rect 4344 464 4353 840
rect 4353 464 4387 840
rect 4387 464 4396 840
rect 4344 462 4396 464
rect 4536 464 4545 840
rect 4545 464 4579 840
rect 4579 464 4588 840
rect 4536 462 4588 464
rect 4728 464 4737 840
rect 4737 464 4771 840
rect 4771 464 4780 840
rect 4728 462 4780 464
rect 4920 464 4929 840
rect 4929 464 4963 840
rect 4963 464 4972 840
rect 4920 462 4972 464
rect 5112 464 5121 840
rect 5121 464 5155 840
rect 5155 464 5164 840
rect 5112 462 5164 464
rect 5304 464 5313 840
rect 5313 464 5347 840
rect 5347 464 5356 840
rect 5304 462 5356 464
rect 5496 464 5505 840
rect 5505 464 5539 840
rect 5539 464 5548 840
rect 5496 462 5548 464
rect 5688 464 5697 840
rect 5697 464 5731 840
rect 5731 464 5740 840
rect 5688 462 5740 464
rect 5880 464 5889 840
rect 5889 464 5923 840
rect 5923 464 5932 840
rect 5880 462 5932 464
rect 120 -1884 172 -1882
rect 120 -2260 129 -1884
rect 129 -2260 163 -1884
rect 163 -2260 172 -1884
rect 312 -1884 364 -1882
rect 312 -2260 321 -1884
rect 321 -2260 355 -1884
rect 355 -2260 364 -1884
rect 504 -1884 556 -1882
rect 504 -2260 513 -1884
rect 513 -2260 547 -1884
rect 547 -2260 556 -1884
rect 696 -1884 748 -1882
rect 696 -2260 705 -1884
rect 705 -2260 739 -1884
rect 739 -2260 748 -1884
rect 888 -1884 940 -1882
rect 888 -2260 897 -1884
rect 897 -2260 931 -1884
rect 931 -2260 940 -1884
rect 1080 -1884 1132 -1882
rect 1080 -2260 1089 -1884
rect 1089 -2260 1123 -1884
rect 1123 -2260 1132 -1884
rect 1272 -1884 1324 -1882
rect 1272 -2260 1281 -1884
rect 1281 -2260 1315 -1884
rect 1315 -2260 1324 -1884
rect 1464 -1884 1516 -1882
rect 1464 -2260 1473 -1884
rect 1473 -2260 1507 -1884
rect 1507 -2260 1516 -1884
rect 1656 -1884 1708 -1882
rect 1656 -2260 1665 -1884
rect 1665 -2260 1699 -1884
rect 1699 -2260 1708 -1884
rect 1848 -1884 1900 -1882
rect 1848 -2260 1857 -1884
rect 1857 -2260 1891 -1884
rect 1891 -2260 1900 -1884
rect 2040 -1884 2092 -1882
rect 2040 -2260 2049 -1884
rect 2049 -2260 2083 -1884
rect 2083 -2260 2092 -1884
rect 2232 -1884 2284 -1882
rect 2232 -2260 2241 -1884
rect 2241 -2260 2275 -1884
rect 2275 -2260 2284 -1884
rect 2424 -1884 2476 -1882
rect 2424 -2260 2433 -1884
rect 2433 -2260 2467 -1884
rect 2467 -2260 2476 -1884
rect 2616 -1884 2668 -1882
rect 2616 -2260 2625 -1884
rect 2625 -2260 2659 -1884
rect 2659 -2260 2668 -1884
rect 2808 -1884 2860 -1882
rect 2808 -2260 2817 -1884
rect 2817 -2260 2851 -1884
rect 2851 -2260 2860 -1884
rect 3000 -1884 3052 -1882
rect 3000 -2260 3009 -1884
rect 3009 -2260 3043 -1884
rect 3043 -2260 3052 -1884
rect 3192 -1884 3244 -1882
rect 3192 -2260 3201 -1884
rect 3201 -2260 3235 -1884
rect 3235 -2260 3244 -1884
rect 3384 -1884 3436 -1882
rect 3384 -2260 3393 -1884
rect 3393 -2260 3427 -1884
rect 3427 -2260 3436 -1884
rect 3576 -1884 3628 -1882
rect 3576 -2260 3585 -1884
rect 3585 -2260 3619 -1884
rect 3619 -2260 3628 -1884
rect 3768 -1884 3820 -1882
rect 3768 -2260 3777 -1884
rect 3777 -2260 3811 -1884
rect 3811 -2260 3820 -1884
rect 3960 -1884 4012 -1882
rect 3960 -2260 3969 -1884
rect 3969 -2260 4003 -1884
rect 4003 -2260 4012 -1884
rect 4152 -1884 4204 -1882
rect 4152 -2260 4161 -1884
rect 4161 -2260 4195 -1884
rect 4195 -2260 4204 -1884
rect 4344 -1884 4396 -1882
rect 4344 -2260 4353 -1884
rect 4353 -2260 4387 -1884
rect 4387 -2260 4396 -1884
rect 4536 -1884 4588 -1882
rect 4536 -2260 4545 -1884
rect 4545 -2260 4579 -1884
rect 4579 -2260 4588 -1884
rect 4728 -1884 4780 -1882
rect 4728 -2260 4737 -1884
rect 4737 -2260 4771 -1884
rect 4771 -2260 4780 -1884
rect 4920 -1884 4972 -1882
rect 4920 -2260 4929 -1884
rect 4929 -2260 4963 -1884
rect 4963 -2260 4972 -1884
rect 5112 -1884 5164 -1882
rect 5112 -2260 5121 -1884
rect 5121 -2260 5155 -1884
rect 5155 -2260 5164 -1884
rect 5304 -1884 5356 -1882
rect 5304 -2260 5313 -1884
rect 5313 -2260 5347 -1884
rect 5347 -2260 5356 -1884
rect 5496 -1884 5548 -1882
rect 5496 -2260 5505 -1884
rect 5505 -2260 5539 -1884
rect 5539 -2260 5548 -1884
rect 5688 -1884 5740 -1882
rect 5688 -2260 5697 -1884
rect 5697 -2260 5731 -1884
rect 5731 -2260 5740 -1884
rect 5880 -1884 5932 -1882
rect 5880 -2260 5889 -1884
rect 5889 -2260 5923 -1884
rect 5923 -2260 5932 -1884
rect 358 -2350 368 -2316
rect 368 -2350 402 -2316
rect 402 -2350 410 -2316
rect 358 -2368 410 -2350
rect 358 -2422 368 -2396
rect 368 -2422 402 -2396
rect 402 -2422 410 -2396
rect 358 -2448 410 -2422
rect 1170 -2376 1234 -2314
rect 1176 -2496 1250 -2426
rect 1938 -2376 2002 -2314
rect 1922 -2496 1996 -2426
rect 2762 -2350 2770 -2316
rect 2770 -2350 2804 -2316
rect 2804 -2350 2814 -2316
rect 2762 -2368 2814 -2350
rect 2762 -2422 2770 -2396
rect 2770 -2422 2804 -2396
rect 2804 -2422 2814 -2396
rect 2762 -2448 2814 -2422
rect 3238 -2350 3248 -2316
rect 3248 -2350 3282 -2316
rect 3282 -2350 3290 -2316
rect 3238 -2368 3290 -2350
rect 3238 -2422 3248 -2396
rect 3248 -2422 3282 -2396
rect 3282 -2422 3290 -2396
rect 3238 -2448 3290 -2422
rect 4050 -2376 4114 -2314
rect 4056 -2496 4130 -2426
rect 120 -2639 172 -2638
rect 120 -3335 129 -2639
rect 129 -3335 163 -2639
rect 163 -3335 172 -2639
rect 120 -3336 172 -3335
rect 312 -2639 364 -2638
rect 312 -3335 321 -2639
rect 321 -3335 355 -2639
rect 355 -3335 364 -2639
rect 312 -3336 364 -3335
rect 4818 -2376 4882 -2314
rect 4802 -2496 4876 -2426
rect 5642 -2350 5650 -2316
rect 5650 -2350 5684 -2316
rect 5684 -2350 5694 -2316
rect 5642 -2368 5694 -2350
rect 5642 -2422 5650 -2396
rect 5650 -2422 5684 -2396
rect 5684 -2422 5694 -2396
rect 5642 -2448 5694 -2422
rect 504 -2639 556 -2638
rect 504 -3335 513 -2639
rect 513 -3335 547 -2639
rect 547 -3335 556 -2639
rect 504 -3336 556 -3335
rect 696 -2639 748 -2638
rect 696 -3335 705 -2639
rect 705 -3335 739 -2639
rect 739 -3335 748 -2639
rect 696 -3336 748 -3335
rect 888 -2639 940 -2638
rect 888 -3335 897 -2639
rect 897 -3335 931 -2639
rect 931 -3335 940 -2639
rect 888 -3336 940 -3335
rect 1080 -2639 1132 -2638
rect 1080 -3335 1089 -2639
rect 1089 -3335 1123 -2639
rect 1123 -3335 1132 -2639
rect 1080 -3336 1132 -3335
rect 1272 -2639 1324 -2638
rect 1272 -3335 1281 -2639
rect 1281 -3335 1315 -2639
rect 1315 -3335 1324 -2639
rect 1272 -3336 1324 -3335
rect 1464 -2639 1516 -2638
rect 1464 -3335 1473 -2639
rect 1473 -3335 1507 -2639
rect 1507 -3335 1516 -2639
rect 1464 -3336 1516 -3335
rect 1656 -2639 1708 -2637
rect 1656 -3335 1665 -2639
rect 1665 -3335 1699 -2639
rect 1699 -3335 1708 -2639
rect 1848 -2639 1900 -2637
rect 1848 -3335 1857 -2639
rect 1857 -3335 1891 -2639
rect 1891 -3335 1900 -2639
rect 2040 -2639 2092 -2637
rect 2040 -3335 2049 -2639
rect 2049 -3335 2083 -2639
rect 2083 -3335 2092 -2639
rect 2232 -2639 2284 -2637
rect 2232 -3335 2241 -2639
rect 2241 -3335 2275 -2639
rect 2275 -3335 2284 -2639
rect 2424 -2639 2476 -2637
rect 2424 -3335 2433 -2639
rect 2433 -3335 2467 -2639
rect 2467 -3335 2476 -2639
rect 2616 -2639 2668 -2637
rect 2616 -3335 2625 -2639
rect 2625 -3335 2659 -2639
rect 2659 -3335 2668 -2639
rect 2808 -2639 2860 -2638
rect 2808 -3335 2817 -2639
rect 2817 -3335 2851 -2639
rect 2851 -3335 2860 -2639
rect 2808 -3336 2860 -3335
rect 3000 -2639 3052 -2638
rect 3000 -3335 3009 -2639
rect 3009 -3335 3043 -2639
rect 3043 -3335 3052 -2639
rect 3000 -3336 3052 -3335
rect 3192 -2639 3244 -2638
rect 3192 -3335 3201 -2639
rect 3201 -3335 3235 -2639
rect 3235 -3335 3244 -2639
rect 3192 -3336 3244 -3335
rect 3384 -2639 3436 -2638
rect 3384 -3335 3393 -2639
rect 3393 -3335 3427 -2639
rect 3427 -3335 3436 -2639
rect 3384 -3336 3436 -3335
rect 3576 -2639 3628 -2638
rect 3576 -3335 3585 -2639
rect 3585 -3335 3619 -2639
rect 3619 -3335 3628 -2639
rect 3576 -3336 3628 -3335
rect 3768 -2639 3820 -2638
rect 3768 -3335 3777 -2639
rect 3777 -3335 3811 -2639
rect 3811 -3335 3820 -2639
rect 3768 -3336 3820 -3335
rect 3960 -2639 4012 -2638
rect 3960 -3335 3969 -2639
rect 3969 -3335 4003 -2639
rect 4003 -3335 4012 -2639
rect 3960 -3336 4012 -3335
rect 4152 -2639 4204 -2638
rect 4152 -3335 4161 -2639
rect 4161 -3335 4195 -2639
rect 4195 -3335 4204 -2639
rect 4152 -3336 4204 -3335
rect 4344 -2639 4396 -2638
rect 4344 -3335 4353 -2639
rect 4353 -3335 4387 -2639
rect 4387 -3335 4396 -2639
rect 4344 -3336 4396 -3335
rect 4536 -2639 4588 -2637
rect 4536 -3335 4545 -2639
rect 4545 -3335 4579 -2639
rect 4579 -3335 4588 -2639
rect 4728 -2639 4780 -2637
rect 4728 -3335 4737 -2639
rect 4737 -3335 4771 -2639
rect 4771 -3335 4780 -2639
rect 4920 -2639 4972 -2637
rect 4920 -3335 4929 -2639
rect 4929 -3335 4963 -2639
rect 4963 -3335 4972 -2639
rect 5112 -2639 5164 -2637
rect 5112 -3335 5121 -2639
rect 5121 -3335 5155 -2639
rect 5155 -3335 5164 -2639
rect 5304 -2639 5356 -2637
rect 5304 -3335 5313 -2639
rect 5313 -3335 5347 -2639
rect 5347 -3335 5356 -2639
rect 5496 -2639 5548 -2637
rect 5496 -3335 5505 -2639
rect 5505 -3335 5539 -2639
rect 5539 -3335 5548 -2639
rect 5688 -2639 5740 -2638
rect 5688 -3335 5697 -2639
rect 5697 -3335 5731 -2639
rect 5731 -3335 5740 -2639
rect 5688 -3336 5740 -3335
rect 5880 -2639 5932 -2638
rect 5880 -3335 5889 -2639
rect 5889 -3335 5923 -2639
rect 5923 -3335 5932 -2639
rect 5880 -3336 5932 -3335
<< metal2 >>
rect 117 1916 174 1932
rect 117 1204 174 1218
rect 309 1916 366 1932
rect 309 1204 366 1218
rect 501 1916 558 1932
rect 501 1204 558 1218
rect 693 1916 750 1932
rect 693 1204 750 1218
rect 885 1916 942 1932
rect 885 1204 942 1218
rect 1077 1916 1134 1932
rect 1077 1204 1134 1218
rect 1269 1916 1326 1932
rect 1269 1204 1326 1218
rect 1461 1916 1518 1932
rect 1461 1204 1518 1218
rect 1654 1915 1711 1931
rect 1654 1203 1711 1217
rect 1846 1915 1903 1931
rect 1846 1203 1903 1217
rect 2038 1915 2095 1931
rect 2038 1203 2095 1217
rect 2230 1915 2287 1931
rect 2230 1203 2287 1217
rect 2422 1915 2479 1931
rect 2422 1203 2479 1217
rect 2614 1915 2671 1931
rect 2614 1203 2671 1217
rect 2806 1916 2863 1932
rect 2806 1204 2863 1218
rect 2997 1916 3055 1932
rect 2997 1204 3055 1218
rect 3189 1916 3246 1932
rect 3189 1204 3246 1218
rect 3381 1916 3438 1932
rect 3381 1204 3438 1218
rect 3573 1916 3630 1932
rect 3573 1204 3630 1218
rect 3765 1916 3822 1932
rect 3765 1204 3822 1218
rect 3957 1916 4014 1932
rect 3957 1204 4014 1218
rect 4149 1916 4206 1932
rect 4149 1204 4206 1218
rect 4341 1916 4398 1932
rect 4341 1204 4398 1218
rect 4534 1915 4591 1931
rect 4534 1203 4591 1217
rect 4726 1915 4783 1931
rect 4726 1203 4783 1217
rect 4918 1915 4975 1931
rect 4918 1203 4975 1217
rect 5110 1915 5167 1931
rect 5110 1203 5167 1217
rect 5302 1915 5359 1931
rect 5302 1203 5359 1217
rect 5494 1915 5551 1931
rect 5494 1203 5551 1217
rect 5686 1916 5743 1932
rect 5686 1204 5743 1218
rect 5878 1916 5935 1932
rect 5878 1204 5935 1218
rect 1166 1076 1260 1086
rect 350 1028 422 1034
rect 350 976 358 1028
rect 410 976 422 1028
rect 1166 1006 1176 1076
rect 1250 1006 1260 1076
rect 1166 996 1260 1006
rect 1912 1076 2006 1086
rect 1912 1006 1922 1076
rect 1996 1006 2006 1076
rect 4046 1076 4140 1086
rect 1912 996 2006 1006
rect 2750 1028 2822 1034
rect 350 962 422 976
rect 2750 976 2762 1028
rect 2814 976 2822 1028
rect 2750 962 2822 976
rect 3230 1028 3302 1034
rect 3230 976 3238 1028
rect 3290 976 3302 1028
rect 4046 1006 4056 1076
rect 4130 1006 4140 1076
rect 4046 996 4140 1006
rect 4792 1076 4886 1086
rect 4792 1006 4802 1076
rect 4876 1006 4886 1076
rect 4792 996 4886 1006
rect 5630 1028 5702 1034
rect 3230 962 3302 976
rect 5630 976 5642 1028
rect 5694 976 5702 1028
rect 5630 962 5702 976
rect 210 948 422 962
rect 210 896 358 948
rect 410 896 422 948
rect 210 894 422 896
rect 117 840 174 856
rect 117 448 174 462
rect 210 166 274 894
rect 309 890 422 894
rect 1170 956 1234 962
rect 309 840 366 856
rect 309 448 366 462
rect 501 840 558 856
rect 501 448 558 462
rect 693 840 750 856
rect 693 448 750 462
rect 885 840 942 856
rect 885 448 942 462
rect 1077 840 1134 856
rect 1077 448 1134 462
rect 1170 166 1234 894
rect 1938 956 2002 962
rect 1269 840 1326 856
rect 1269 448 1326 462
rect 1461 840 1518 856
rect 1461 448 1518 462
rect 1654 840 1711 856
rect 1654 448 1711 462
rect 1846 840 1903 856
rect 1846 448 1903 462
rect 1938 166 2002 894
rect 2750 948 2962 962
rect 2750 896 2762 948
rect 2814 896 2962 948
rect 2750 894 2962 896
rect 2750 890 2863 894
rect 2038 840 2095 856
rect 2038 448 2095 462
rect 2230 840 2287 856
rect 2230 448 2287 462
rect 2422 840 2479 856
rect 2422 448 2479 462
rect 2614 840 2671 856
rect 2614 448 2671 462
rect 2806 840 2863 856
rect 2806 448 2863 462
rect 2898 166 2962 894
rect 3090 948 3302 962
rect 3090 896 3238 948
rect 3290 896 3302 948
rect 3090 894 3302 896
rect 2997 840 3055 856
rect 2997 448 3055 462
rect 3090 166 3154 894
rect 3189 890 3302 894
rect 4050 956 4114 962
rect 3189 840 3246 856
rect 3189 448 3246 462
rect 3381 840 3438 856
rect 3381 448 3438 462
rect 3573 840 3630 856
rect 3573 448 3630 462
rect 3765 840 3822 856
rect 3765 448 3822 462
rect 3957 840 4014 856
rect 3957 448 4014 462
rect 4050 166 4114 894
rect 4818 956 4882 962
rect 4149 840 4206 856
rect 4149 448 4206 462
rect 4341 840 4398 856
rect 4341 448 4398 462
rect 4534 840 4591 856
rect 4534 448 4591 462
rect 4726 840 4783 856
rect 4726 448 4783 462
rect 4818 166 4882 894
rect 5630 948 5842 962
rect 5630 896 5642 948
rect 5694 896 5842 948
rect 5630 894 5842 896
rect 5630 890 5743 894
rect 4918 840 4975 856
rect 4918 448 4975 462
rect 5110 840 5167 856
rect 5110 448 5167 462
rect 5302 840 5359 856
rect 5302 448 5359 462
rect 5494 840 5551 856
rect 5494 448 5551 462
rect 5686 840 5743 856
rect 5686 448 5743 462
rect 5778 166 5842 894
rect 5878 840 5935 856
rect 5878 448 5935 462
rect 208 160 276 166
rect 208 104 214 160
rect 270 104 276 160
rect 208 78 276 104
rect 208 22 214 78
rect 270 22 276 78
rect 208 2 276 22
rect 1168 160 1236 166
rect 1168 104 1174 160
rect 1230 104 1236 160
rect 1168 78 1236 104
rect 1168 22 1174 78
rect 1230 22 1236 78
rect 1168 2 1236 22
rect 1936 160 2004 166
rect 1936 104 1942 160
rect 1998 104 2004 160
rect 1936 78 2004 104
rect 1936 22 1942 78
rect 1998 22 2004 78
rect 1936 2 2004 22
rect 2896 160 2964 166
rect 2896 104 2902 160
rect 2958 104 2964 160
rect 2896 78 2964 104
rect 2896 22 2902 78
rect 2958 22 2964 78
rect 2896 2 2964 22
rect 3088 160 3156 166
rect 3088 104 3094 160
rect 3150 104 3156 160
rect 3088 78 3156 104
rect 3088 22 3094 78
rect 3150 22 3156 78
rect 3088 2 3156 22
rect 4048 160 4116 166
rect 4048 104 4054 160
rect 4110 104 4116 160
rect 4048 78 4116 104
rect 4048 22 4054 78
rect 4110 22 4116 78
rect 4048 2 4116 22
rect 4816 160 4884 166
rect 4816 104 4822 160
rect 4878 104 4884 160
rect 4816 78 4884 104
rect 4816 22 4822 78
rect 4878 22 4884 78
rect 4816 2 4884 22
rect 5776 160 5844 166
rect 5776 104 5782 160
rect 5838 104 5844 160
rect 5776 78 5844 104
rect 5776 22 5782 78
rect 5838 22 5844 78
rect 5776 2 5844 22
rect 208 -1442 276 -1422
rect 208 -1498 214 -1442
rect 270 -1498 276 -1442
rect 208 -1524 276 -1498
rect 208 -1580 214 -1524
rect 270 -1580 276 -1524
rect 208 -1586 276 -1580
rect 1168 -1442 1236 -1422
rect 1168 -1498 1174 -1442
rect 1230 -1498 1236 -1442
rect 1168 -1524 1236 -1498
rect 1168 -1580 1174 -1524
rect 1230 -1580 1236 -1524
rect 1168 -1586 1236 -1580
rect 1936 -1442 2004 -1422
rect 1936 -1498 1942 -1442
rect 1998 -1498 2004 -1442
rect 1936 -1524 2004 -1498
rect 1936 -1580 1942 -1524
rect 1998 -1580 2004 -1524
rect 1936 -1586 2004 -1580
rect 2896 -1442 2964 -1422
rect 2896 -1498 2902 -1442
rect 2958 -1498 2964 -1442
rect 2896 -1524 2964 -1498
rect 2896 -1580 2902 -1524
rect 2958 -1580 2964 -1524
rect 2896 -1586 2964 -1580
rect 3088 -1442 3156 -1422
rect 3088 -1498 3094 -1442
rect 3150 -1498 3156 -1442
rect 3088 -1524 3156 -1498
rect 3088 -1580 3094 -1524
rect 3150 -1580 3156 -1524
rect 3088 -1586 3156 -1580
rect 4048 -1442 4116 -1422
rect 4048 -1498 4054 -1442
rect 4110 -1498 4116 -1442
rect 4048 -1524 4116 -1498
rect 4048 -1580 4054 -1524
rect 4110 -1580 4116 -1524
rect 4048 -1586 4116 -1580
rect 4816 -1442 4884 -1422
rect 4816 -1498 4822 -1442
rect 4878 -1498 4884 -1442
rect 4816 -1524 4884 -1498
rect 4816 -1580 4822 -1524
rect 4878 -1580 4884 -1524
rect 4816 -1586 4884 -1580
rect 5776 -1442 5844 -1422
rect 5776 -1498 5782 -1442
rect 5838 -1498 5844 -1442
rect 5776 -1524 5844 -1498
rect 5776 -1580 5782 -1524
rect 5838 -1580 5844 -1524
rect 5776 -1586 5844 -1580
rect 117 -1882 174 -1868
rect 117 -2276 174 -2260
rect 210 -2314 274 -1586
rect 309 -1882 366 -1868
rect 309 -2276 366 -2260
rect 501 -1882 558 -1868
rect 501 -2276 558 -2260
rect 693 -1882 750 -1868
rect 693 -2276 750 -2260
rect 885 -1882 942 -1868
rect 885 -2276 942 -2260
rect 1077 -1882 1134 -1868
rect 1077 -2276 1134 -2260
rect 309 -2314 422 -2310
rect 210 -2316 422 -2314
rect 210 -2368 358 -2316
rect 410 -2368 422 -2316
rect 210 -2382 422 -2368
rect 1170 -2314 1234 -1586
rect 1269 -1882 1326 -1868
rect 1269 -2276 1326 -2260
rect 1461 -1882 1518 -1868
rect 1461 -2276 1518 -2260
rect 1654 -1882 1711 -1868
rect 1654 -2276 1711 -2260
rect 1846 -1882 1903 -1868
rect 1846 -2276 1903 -2260
rect 1170 -2382 1234 -2376
rect 1938 -2314 2002 -1586
rect 2038 -1882 2095 -1868
rect 2038 -2276 2095 -2260
rect 2230 -1882 2287 -1868
rect 2230 -2276 2287 -2260
rect 2422 -1882 2479 -1868
rect 2422 -2276 2479 -2260
rect 2614 -1882 2671 -1868
rect 2614 -2276 2671 -2260
rect 2806 -1882 2863 -1868
rect 2806 -2276 2863 -2260
rect 1938 -2382 2002 -2376
rect 2750 -2314 2863 -2310
rect 2898 -2314 2962 -1586
rect 2997 -1882 3055 -1868
rect 2997 -2276 3055 -2260
rect 2750 -2316 2962 -2314
rect 2750 -2368 2762 -2316
rect 2814 -2368 2962 -2316
rect 2750 -2382 2962 -2368
rect 3090 -2314 3154 -1586
rect 3189 -1882 3246 -1868
rect 3189 -2276 3246 -2260
rect 3381 -1882 3438 -1868
rect 3381 -2276 3438 -2260
rect 3573 -1882 3630 -1868
rect 3573 -2276 3630 -2260
rect 3765 -1882 3822 -1868
rect 3765 -2276 3822 -2260
rect 3957 -1882 4014 -1868
rect 3957 -2276 4014 -2260
rect 3189 -2314 3302 -2310
rect 3090 -2316 3302 -2314
rect 3090 -2368 3238 -2316
rect 3290 -2368 3302 -2316
rect 3090 -2382 3302 -2368
rect 4050 -2314 4114 -1586
rect 4149 -1882 4206 -1868
rect 4149 -2276 4206 -2260
rect 4341 -1882 4398 -1868
rect 4341 -2276 4398 -2260
rect 4534 -1882 4591 -1868
rect 4534 -2276 4591 -2260
rect 4726 -1882 4783 -1868
rect 4726 -2276 4783 -2260
rect 4050 -2382 4114 -2376
rect 4818 -2314 4882 -1586
rect 4918 -1882 4975 -1868
rect 4918 -2276 4975 -2260
rect 5110 -1882 5167 -1868
rect 5110 -2276 5167 -2260
rect 5302 -1882 5359 -1868
rect 5302 -2276 5359 -2260
rect 5494 -1882 5551 -1868
rect 5494 -2276 5551 -2260
rect 5686 -1882 5743 -1868
rect 5686 -2276 5743 -2260
rect 4818 -2382 4882 -2376
rect 5630 -2314 5743 -2310
rect 5778 -2314 5842 -1586
rect 5878 -1882 5935 -1868
rect 5878 -2276 5935 -2260
rect 5630 -2316 5842 -2314
rect 5630 -2368 5642 -2316
rect 5694 -2368 5842 -2316
rect 5630 -2382 5842 -2368
rect 350 -2396 422 -2382
rect 350 -2448 358 -2396
rect 410 -2448 422 -2396
rect 2750 -2396 2822 -2382
rect 350 -2454 422 -2448
rect 1166 -2426 1260 -2416
rect 1166 -2496 1176 -2426
rect 1250 -2496 1260 -2426
rect 1166 -2506 1260 -2496
rect 1912 -2426 2006 -2416
rect 1912 -2496 1922 -2426
rect 1996 -2496 2006 -2426
rect 2750 -2448 2762 -2396
rect 2814 -2448 2822 -2396
rect 2750 -2454 2822 -2448
rect 3230 -2396 3302 -2382
rect 3230 -2448 3238 -2396
rect 3290 -2448 3302 -2396
rect 5630 -2396 5702 -2382
rect 3230 -2454 3302 -2448
rect 4046 -2426 4140 -2416
rect 1912 -2506 2006 -2496
rect 4046 -2496 4056 -2426
rect 4130 -2496 4140 -2426
rect 4046 -2506 4140 -2496
rect 4792 -2426 4886 -2416
rect 4792 -2496 4802 -2426
rect 4876 -2496 4886 -2426
rect 5630 -2448 5642 -2396
rect 5694 -2448 5702 -2396
rect 5630 -2454 5702 -2448
rect 4792 -2506 4886 -2496
rect 117 -2638 174 -2624
rect 117 -3352 174 -3336
rect 309 -2638 366 -2624
rect 309 -3352 366 -3336
rect 501 -2638 558 -2624
rect 501 -3352 558 -3336
rect 693 -2638 750 -2624
rect 693 -3352 750 -3336
rect 885 -2638 942 -2624
rect 885 -3352 942 -3336
rect 1077 -2638 1134 -2624
rect 1077 -3352 1134 -3336
rect 1269 -2638 1326 -2624
rect 1269 -3352 1326 -3336
rect 1461 -2638 1518 -2624
rect 1461 -3352 1518 -3336
rect 1654 -2637 1711 -2623
rect 1654 -3351 1711 -3335
rect 1846 -2637 1903 -2623
rect 1846 -3351 1903 -3335
rect 2038 -2637 2095 -2623
rect 2038 -3351 2095 -3335
rect 2230 -2637 2287 -2623
rect 2230 -3351 2287 -3335
rect 2422 -2637 2479 -2623
rect 2422 -3351 2479 -3335
rect 2614 -2637 2671 -2623
rect 2614 -3351 2671 -3335
rect 2806 -2638 2863 -2624
rect 2806 -3352 2863 -3336
rect 2997 -2638 3055 -2624
rect 2997 -3352 3055 -3336
rect 3189 -2638 3246 -2624
rect 3189 -3352 3246 -3336
rect 3381 -2638 3438 -2624
rect 3381 -3352 3438 -3336
rect 3573 -2638 3630 -2624
rect 3573 -3352 3630 -3336
rect 3765 -2638 3822 -2624
rect 3765 -3352 3822 -3336
rect 3957 -2638 4014 -2624
rect 3957 -3352 4014 -3336
rect 4149 -2638 4206 -2624
rect 4149 -3352 4206 -3336
rect 4341 -2638 4398 -2624
rect 4341 -3352 4398 -3336
rect 4534 -2637 4591 -2623
rect 4534 -3351 4591 -3335
rect 4726 -2637 4783 -2623
rect 4726 -3351 4783 -3335
rect 4918 -2637 4975 -2623
rect 4918 -3351 4975 -3335
rect 5110 -2637 5167 -2623
rect 5110 -3351 5167 -3335
rect 5302 -2637 5359 -2623
rect 5302 -3351 5359 -3335
rect 5494 -2637 5551 -2623
rect 5494 -3351 5551 -3335
rect 5686 -2638 5743 -2624
rect 5686 -3352 5743 -3336
rect 5878 -2638 5935 -2624
rect 5878 -3352 5935 -3336
<< via2 >>
rect 117 1218 120 1916
rect 120 1218 172 1916
rect 172 1218 174 1916
rect 309 1218 312 1916
rect 312 1218 364 1916
rect 364 1218 366 1916
rect 501 1218 504 1916
rect 504 1218 556 1916
rect 556 1218 558 1916
rect 693 1218 696 1916
rect 696 1218 748 1916
rect 748 1218 750 1916
rect 885 1218 888 1916
rect 888 1218 940 1916
rect 940 1218 942 1916
rect 1077 1218 1080 1916
rect 1080 1218 1132 1916
rect 1132 1218 1134 1916
rect 1269 1218 1272 1916
rect 1272 1218 1324 1916
rect 1324 1218 1326 1916
rect 1461 1218 1464 1916
rect 1464 1218 1516 1916
rect 1516 1218 1518 1916
rect 1654 1217 1656 1915
rect 1656 1217 1708 1915
rect 1708 1217 1711 1915
rect 1846 1217 1848 1915
rect 1848 1217 1900 1915
rect 1900 1217 1903 1915
rect 2038 1217 2040 1915
rect 2040 1217 2092 1915
rect 2092 1217 2095 1915
rect 2230 1217 2232 1915
rect 2232 1217 2284 1915
rect 2284 1217 2287 1915
rect 2422 1217 2424 1915
rect 2424 1217 2476 1915
rect 2476 1217 2479 1915
rect 2614 1217 2616 1915
rect 2616 1217 2668 1915
rect 2668 1217 2671 1915
rect 2806 1218 2808 1916
rect 2808 1218 2860 1916
rect 2860 1218 2863 1916
rect 2997 1218 3000 1916
rect 3000 1218 3052 1916
rect 3052 1218 3055 1916
rect 3189 1218 3192 1916
rect 3192 1218 3244 1916
rect 3244 1218 3246 1916
rect 3381 1218 3384 1916
rect 3384 1218 3436 1916
rect 3436 1218 3438 1916
rect 3573 1218 3576 1916
rect 3576 1218 3628 1916
rect 3628 1218 3630 1916
rect 3765 1218 3768 1916
rect 3768 1218 3820 1916
rect 3820 1218 3822 1916
rect 3957 1218 3960 1916
rect 3960 1218 4012 1916
rect 4012 1218 4014 1916
rect 4149 1218 4152 1916
rect 4152 1218 4204 1916
rect 4204 1218 4206 1916
rect 4341 1218 4344 1916
rect 4344 1218 4396 1916
rect 4396 1218 4398 1916
rect 4534 1217 4536 1915
rect 4536 1217 4588 1915
rect 4588 1217 4591 1915
rect 4726 1217 4728 1915
rect 4728 1217 4780 1915
rect 4780 1217 4783 1915
rect 4918 1217 4920 1915
rect 4920 1217 4972 1915
rect 4972 1217 4975 1915
rect 5110 1217 5112 1915
rect 5112 1217 5164 1915
rect 5164 1217 5167 1915
rect 5302 1217 5304 1915
rect 5304 1217 5356 1915
rect 5356 1217 5359 1915
rect 5494 1217 5496 1915
rect 5496 1217 5548 1915
rect 5548 1217 5551 1915
rect 5686 1218 5688 1916
rect 5688 1218 5740 1916
rect 5740 1218 5743 1916
rect 5878 1218 5880 1916
rect 5880 1218 5932 1916
rect 5932 1218 5935 1916
rect 1176 1006 1250 1076
rect 1922 1006 1996 1076
rect 4056 1006 4130 1076
rect 4802 1006 4876 1076
rect 117 462 120 840
rect 120 462 172 840
rect 172 462 174 840
rect 309 462 312 840
rect 312 462 364 840
rect 364 462 366 840
rect 501 462 504 840
rect 504 462 556 840
rect 556 462 558 840
rect 693 462 696 840
rect 696 462 748 840
rect 748 462 750 840
rect 885 462 888 840
rect 888 462 940 840
rect 940 462 942 840
rect 1077 462 1080 840
rect 1080 462 1132 840
rect 1132 462 1134 840
rect 1269 462 1272 840
rect 1272 462 1324 840
rect 1324 462 1326 840
rect 1461 462 1464 840
rect 1464 462 1516 840
rect 1516 462 1518 840
rect 1654 462 1656 840
rect 1656 462 1708 840
rect 1708 462 1711 840
rect 1846 462 1848 840
rect 1848 462 1900 840
rect 1900 462 1903 840
rect 2038 462 2040 840
rect 2040 462 2092 840
rect 2092 462 2095 840
rect 2230 462 2232 840
rect 2232 462 2284 840
rect 2284 462 2287 840
rect 2422 462 2424 840
rect 2424 462 2476 840
rect 2476 462 2479 840
rect 2614 462 2616 840
rect 2616 462 2668 840
rect 2668 462 2671 840
rect 2806 462 2808 840
rect 2808 462 2860 840
rect 2860 462 2863 840
rect 2997 462 3000 840
rect 3000 462 3052 840
rect 3052 462 3055 840
rect 3189 462 3192 840
rect 3192 462 3244 840
rect 3244 462 3246 840
rect 3381 462 3384 840
rect 3384 462 3436 840
rect 3436 462 3438 840
rect 3573 462 3576 840
rect 3576 462 3628 840
rect 3628 462 3630 840
rect 3765 462 3768 840
rect 3768 462 3820 840
rect 3820 462 3822 840
rect 3957 462 3960 840
rect 3960 462 4012 840
rect 4012 462 4014 840
rect 4149 462 4152 840
rect 4152 462 4204 840
rect 4204 462 4206 840
rect 4341 462 4344 840
rect 4344 462 4396 840
rect 4396 462 4398 840
rect 4534 462 4536 840
rect 4536 462 4588 840
rect 4588 462 4591 840
rect 4726 462 4728 840
rect 4728 462 4780 840
rect 4780 462 4783 840
rect 4918 462 4920 840
rect 4920 462 4972 840
rect 4972 462 4975 840
rect 5110 462 5112 840
rect 5112 462 5164 840
rect 5164 462 5167 840
rect 5302 462 5304 840
rect 5304 462 5356 840
rect 5356 462 5359 840
rect 5494 462 5496 840
rect 5496 462 5548 840
rect 5548 462 5551 840
rect 5686 462 5688 840
rect 5688 462 5740 840
rect 5740 462 5743 840
rect 5878 462 5880 840
rect 5880 462 5932 840
rect 5932 462 5935 840
rect 214 104 270 160
rect 214 22 270 78
rect 1174 104 1230 160
rect 1174 22 1230 78
rect 1942 104 1998 160
rect 1942 22 1998 78
rect 2902 104 2958 160
rect 2902 22 2958 78
rect 3094 104 3150 160
rect 3094 22 3150 78
rect 4054 104 4110 160
rect 4054 22 4110 78
rect 4822 104 4878 160
rect 4822 22 4878 78
rect 5782 104 5838 160
rect 5782 22 5838 78
rect 214 -1498 270 -1442
rect 214 -1580 270 -1524
rect 1174 -1498 1230 -1442
rect 1174 -1580 1230 -1524
rect 1942 -1498 1998 -1442
rect 1942 -1580 1998 -1524
rect 2902 -1498 2958 -1442
rect 2902 -1580 2958 -1524
rect 3094 -1498 3150 -1442
rect 3094 -1580 3150 -1524
rect 4054 -1498 4110 -1442
rect 4054 -1580 4110 -1524
rect 4822 -1498 4878 -1442
rect 4822 -1580 4878 -1524
rect 5782 -1498 5838 -1442
rect 5782 -1580 5838 -1524
rect 117 -2260 120 -1882
rect 120 -2260 172 -1882
rect 172 -2260 174 -1882
rect 309 -2260 312 -1882
rect 312 -2260 364 -1882
rect 364 -2260 366 -1882
rect 501 -2260 504 -1882
rect 504 -2260 556 -1882
rect 556 -2260 558 -1882
rect 693 -2260 696 -1882
rect 696 -2260 748 -1882
rect 748 -2260 750 -1882
rect 885 -2260 888 -1882
rect 888 -2260 940 -1882
rect 940 -2260 942 -1882
rect 1077 -2260 1080 -1882
rect 1080 -2260 1132 -1882
rect 1132 -2260 1134 -1882
rect 1269 -2260 1272 -1882
rect 1272 -2260 1324 -1882
rect 1324 -2260 1326 -1882
rect 1461 -2260 1464 -1882
rect 1464 -2260 1516 -1882
rect 1516 -2260 1518 -1882
rect 1654 -2260 1656 -1882
rect 1656 -2260 1708 -1882
rect 1708 -2260 1711 -1882
rect 1846 -2260 1848 -1882
rect 1848 -2260 1900 -1882
rect 1900 -2260 1903 -1882
rect 2038 -2260 2040 -1882
rect 2040 -2260 2092 -1882
rect 2092 -2260 2095 -1882
rect 2230 -2260 2232 -1882
rect 2232 -2260 2284 -1882
rect 2284 -2260 2287 -1882
rect 2422 -2260 2424 -1882
rect 2424 -2260 2476 -1882
rect 2476 -2260 2479 -1882
rect 2614 -2260 2616 -1882
rect 2616 -2260 2668 -1882
rect 2668 -2260 2671 -1882
rect 2806 -2260 2808 -1882
rect 2808 -2260 2860 -1882
rect 2860 -2260 2863 -1882
rect 2997 -2260 3000 -1882
rect 3000 -2260 3052 -1882
rect 3052 -2260 3055 -1882
rect 3189 -2260 3192 -1882
rect 3192 -2260 3244 -1882
rect 3244 -2260 3246 -1882
rect 3381 -2260 3384 -1882
rect 3384 -2260 3436 -1882
rect 3436 -2260 3438 -1882
rect 3573 -2260 3576 -1882
rect 3576 -2260 3628 -1882
rect 3628 -2260 3630 -1882
rect 3765 -2260 3768 -1882
rect 3768 -2260 3820 -1882
rect 3820 -2260 3822 -1882
rect 3957 -2260 3960 -1882
rect 3960 -2260 4012 -1882
rect 4012 -2260 4014 -1882
rect 4149 -2260 4152 -1882
rect 4152 -2260 4204 -1882
rect 4204 -2260 4206 -1882
rect 4341 -2260 4344 -1882
rect 4344 -2260 4396 -1882
rect 4396 -2260 4398 -1882
rect 4534 -2260 4536 -1882
rect 4536 -2260 4588 -1882
rect 4588 -2260 4591 -1882
rect 4726 -2260 4728 -1882
rect 4728 -2260 4780 -1882
rect 4780 -2260 4783 -1882
rect 4918 -2260 4920 -1882
rect 4920 -2260 4972 -1882
rect 4972 -2260 4975 -1882
rect 5110 -2260 5112 -1882
rect 5112 -2260 5164 -1882
rect 5164 -2260 5167 -1882
rect 5302 -2260 5304 -1882
rect 5304 -2260 5356 -1882
rect 5356 -2260 5359 -1882
rect 5494 -2260 5496 -1882
rect 5496 -2260 5548 -1882
rect 5548 -2260 5551 -1882
rect 5686 -2260 5688 -1882
rect 5688 -2260 5740 -1882
rect 5740 -2260 5743 -1882
rect 5878 -2260 5880 -1882
rect 5880 -2260 5932 -1882
rect 5932 -2260 5935 -1882
rect 1176 -2496 1250 -2426
rect 1922 -2496 1996 -2426
rect 4056 -2496 4130 -2426
rect 4802 -2496 4876 -2426
rect 117 -3336 120 -2638
rect 120 -3336 172 -2638
rect 172 -3336 174 -2638
rect 309 -3336 312 -2638
rect 312 -3336 364 -2638
rect 364 -3336 366 -2638
rect 501 -3336 504 -2638
rect 504 -3336 556 -2638
rect 556 -3336 558 -2638
rect 693 -3336 696 -2638
rect 696 -3336 748 -2638
rect 748 -3336 750 -2638
rect 885 -3336 888 -2638
rect 888 -3336 940 -2638
rect 940 -3336 942 -2638
rect 1077 -3336 1080 -2638
rect 1080 -3336 1132 -2638
rect 1132 -3336 1134 -2638
rect 1269 -3336 1272 -2638
rect 1272 -3336 1324 -2638
rect 1324 -3336 1326 -2638
rect 1461 -3336 1464 -2638
rect 1464 -3336 1516 -2638
rect 1516 -3336 1518 -2638
rect 1654 -3335 1656 -2637
rect 1656 -3335 1708 -2637
rect 1708 -3335 1711 -2637
rect 1846 -3335 1848 -2637
rect 1848 -3335 1900 -2637
rect 1900 -3335 1903 -2637
rect 2038 -3335 2040 -2637
rect 2040 -3335 2092 -2637
rect 2092 -3335 2095 -2637
rect 2230 -3335 2232 -2637
rect 2232 -3335 2284 -2637
rect 2284 -3335 2287 -2637
rect 2422 -3335 2424 -2637
rect 2424 -3335 2476 -2637
rect 2476 -3335 2479 -2637
rect 2614 -3335 2616 -2637
rect 2616 -3335 2668 -2637
rect 2668 -3335 2671 -2637
rect 2806 -3336 2808 -2638
rect 2808 -3336 2860 -2638
rect 2860 -3336 2863 -2638
rect 2997 -3336 3000 -2638
rect 3000 -3336 3052 -2638
rect 3052 -3336 3055 -2638
rect 3189 -3336 3192 -2638
rect 3192 -3336 3244 -2638
rect 3244 -3336 3246 -2638
rect 3381 -3336 3384 -2638
rect 3384 -3336 3436 -2638
rect 3436 -3336 3438 -2638
rect 3573 -3336 3576 -2638
rect 3576 -3336 3628 -2638
rect 3628 -3336 3630 -2638
rect 3765 -3336 3768 -2638
rect 3768 -3336 3820 -2638
rect 3820 -3336 3822 -2638
rect 3957 -3336 3960 -2638
rect 3960 -3336 4012 -2638
rect 4012 -3336 4014 -2638
rect 4149 -3336 4152 -2638
rect 4152 -3336 4204 -2638
rect 4204 -3336 4206 -2638
rect 4341 -3336 4344 -2638
rect 4344 -3336 4396 -2638
rect 4396 -3336 4398 -2638
rect 4534 -3335 4536 -2637
rect 4536 -3335 4588 -2637
rect 4588 -3335 4591 -2637
rect 4726 -3335 4728 -2637
rect 4728 -3335 4780 -2637
rect 4780 -3335 4783 -2637
rect 4918 -3335 4920 -2637
rect 4920 -3335 4972 -2637
rect 4972 -3335 4975 -2637
rect 5110 -3335 5112 -2637
rect 5112 -3335 5164 -2637
rect 5164 -3335 5167 -2637
rect 5302 -3335 5304 -2637
rect 5304 -3335 5356 -2637
rect 5356 -3335 5359 -2637
rect 5494 -3335 5496 -2637
rect 5496 -3335 5548 -2637
rect 5548 -3335 5551 -2637
rect 5686 -3336 5688 -2638
rect 5688 -3336 5740 -2638
rect 5740 -3336 5743 -2638
rect 5878 -3336 5880 -2638
rect 5880 -3336 5932 -2638
rect 5932 -3336 5935 -2638
<< metal3 >>
rect 112 1916 180 1932
rect 112 1218 117 1916
rect 174 1218 180 1916
rect 112 1204 180 1218
rect 304 1916 372 1932
rect 304 1218 309 1916
rect 366 1218 372 1916
rect 304 1204 372 1218
rect 496 1916 564 1932
rect 496 1218 501 1916
rect 558 1218 564 1916
rect 112 840 180 856
rect 112 462 117 840
rect 174 462 180 840
rect 112 448 180 462
rect 304 840 372 856
rect 304 462 309 840
rect 366 462 372 840
rect 304 286 372 462
rect 496 840 564 1218
rect 496 462 501 840
rect 558 462 564 840
rect 304 226 400 286
rect 496 226 564 462
rect 688 1916 756 1932
rect 688 1218 693 1916
rect 750 1218 756 1916
rect 688 840 756 1218
rect 688 462 693 840
rect 750 462 756 840
rect 688 226 756 462
rect 880 1916 948 1932
rect 880 1218 885 1916
rect 942 1218 948 1916
rect 880 840 948 1218
rect 880 462 885 840
rect 942 462 948 840
rect 880 226 948 462
rect 1072 1916 1140 1932
rect 1072 1218 1077 1916
rect 1134 1218 1140 1916
rect 1072 1086 1140 1218
rect 1264 1916 1332 1932
rect 1264 1218 1269 1916
rect 1326 1258 1332 1916
rect 1456 1916 1524 1932
rect 1326 1218 1396 1258
rect 1264 1198 1396 1218
rect 1072 1076 1260 1086
rect 1072 1006 1176 1076
rect 1250 1006 1260 1076
rect 1072 996 1260 1006
rect 1072 840 1140 996
rect 1328 852 1396 1198
rect 1072 462 1077 840
rect 1134 462 1140 840
rect 1072 286 1140 462
rect 1044 226 1140 286
rect 1264 840 1396 852
rect 1264 462 1269 840
rect 1326 790 1396 840
rect 1456 1218 1461 1916
rect 1518 1218 1524 1916
rect 1456 840 1524 1218
rect 1326 462 1332 790
rect 1264 286 1332 462
rect 1456 462 1461 840
rect 1518 462 1524 840
rect 1264 226 1360 286
rect 1456 226 1524 462
rect 204 160 280 166
rect 204 104 214 160
rect 270 104 280 160
rect 340 120 1104 226
rect 1164 160 1240 166
rect 204 78 280 104
rect 204 22 214 78
rect 270 22 280 78
rect 204 2 280 22
rect 880 -100 950 120
rect 1164 104 1174 160
rect 1230 104 1240 160
rect 1300 120 1524 226
rect 1164 78 1240 104
rect 1164 40 1174 78
rect 1160 22 1174 40
rect 1230 22 1240 78
rect 870 -110 960 -100
rect 870 -190 880 -110
rect 950 -190 960 -110
rect 870 -200 960 -190
rect 1160 -1060 1240 22
rect 1456 0 1524 120
rect 1648 1915 1716 1931
rect 1648 1217 1654 1915
rect 1711 1217 1716 1915
rect 1840 1915 1908 1931
rect 1840 1258 1846 1915
rect 1648 840 1716 1217
rect 1648 462 1654 840
rect 1711 462 1716 840
rect 1776 1217 1846 1258
rect 1903 1217 1908 1915
rect 1776 1198 1908 1217
rect 2032 1915 2100 1931
rect 2032 1217 2038 1915
rect 2095 1217 2100 1915
rect 1776 852 1844 1198
rect 2032 1086 2100 1217
rect 1912 1076 2100 1086
rect 1912 1006 1922 1076
rect 1996 1006 2100 1076
rect 1912 996 2100 1006
rect 1776 840 1908 852
rect 1776 790 1846 840
rect 1648 226 1716 462
rect 1840 462 1846 790
rect 1903 462 1908 840
rect 1840 286 1908 462
rect 1812 226 1908 286
rect 2032 840 2100 996
rect 2032 462 2038 840
rect 2095 462 2100 840
rect 2032 286 2100 462
rect 2224 1915 2292 1931
rect 2224 1217 2230 1915
rect 2287 1217 2292 1915
rect 2224 840 2292 1217
rect 2224 462 2230 840
rect 2287 462 2292 840
rect 2032 226 2128 286
rect 2224 226 2292 462
rect 2416 1915 2484 1931
rect 2416 1217 2422 1915
rect 2479 1217 2484 1915
rect 2416 840 2484 1217
rect 2416 462 2422 840
rect 2479 462 2484 840
rect 2416 226 2484 462
rect 2608 1915 2676 1931
rect 2608 1217 2614 1915
rect 2671 1217 2676 1915
rect 2608 840 2676 1217
rect 2800 1916 2868 1932
rect 2800 1218 2806 1916
rect 2863 1218 2868 1916
rect 2800 1110 2868 1218
rect 2992 1916 3060 1932
rect 2992 1218 2997 1916
rect 3055 1218 3060 1916
rect 2992 1110 3060 1218
rect 3184 1916 3252 1932
rect 3184 1218 3189 1916
rect 3246 1218 3252 1916
rect 3184 1204 3252 1218
rect 3376 1916 3444 1932
rect 3376 1218 3381 1916
rect 3438 1218 3444 1916
rect 2608 462 2614 840
rect 2671 462 2676 840
rect 2608 226 2676 462
rect 2800 840 2868 856
rect 2800 462 2806 840
rect 2863 462 2868 840
rect 2800 286 2868 462
rect 2992 840 3060 856
rect 2992 462 2997 840
rect 3055 462 3060 840
rect 2992 448 3060 462
rect 3184 840 3252 856
rect 3184 462 3189 840
rect 3246 462 3252 840
rect 2772 226 2868 286
rect 3184 286 3252 462
rect 3376 840 3444 1218
rect 3376 462 3381 840
rect 3438 462 3444 840
rect 3184 226 3280 286
rect 3376 226 3444 462
rect 3568 1916 3636 1932
rect 3568 1218 3573 1916
rect 3630 1218 3636 1916
rect 3568 840 3636 1218
rect 3568 462 3573 840
rect 3630 462 3636 840
rect 3568 226 3636 462
rect 3760 1916 3828 1932
rect 3760 1218 3765 1916
rect 3822 1218 3828 1916
rect 3760 840 3828 1218
rect 3760 462 3765 840
rect 3822 462 3828 840
rect 3760 226 3828 462
rect 3952 1916 4020 1932
rect 3952 1218 3957 1916
rect 4014 1218 4020 1916
rect 3952 1086 4020 1218
rect 4144 1916 4212 1932
rect 4144 1218 4149 1916
rect 4206 1258 4212 1916
rect 4336 1916 4404 1932
rect 4206 1218 4276 1258
rect 4144 1198 4276 1218
rect 3952 1076 4140 1086
rect 3952 1006 4056 1076
rect 4130 1006 4140 1076
rect 3952 996 4140 1006
rect 3952 840 4020 996
rect 4208 852 4276 1198
rect 3952 462 3957 840
rect 4014 462 4020 840
rect 3952 286 4020 462
rect 3924 226 4020 286
rect 4144 840 4276 852
rect 4144 462 4149 840
rect 4206 790 4276 840
rect 4336 1218 4341 1916
rect 4398 1218 4404 1916
rect 4336 840 4404 1218
rect 4206 462 4212 790
rect 4144 286 4212 462
rect 4336 462 4341 840
rect 4398 462 4404 840
rect 4144 226 4240 286
rect 4336 226 4404 462
rect 1648 120 1872 226
rect 1932 160 2008 166
rect 1460 -870 1520 -30
rect 1648 -524 1716 120
rect 1932 104 1942 160
rect 1998 104 2008 160
rect 2068 120 2832 226
rect 2892 160 2968 166
rect 1932 78 2008 104
rect 1932 22 1942 78
rect 1998 22 2008 78
rect 1932 2 2008 22
rect 1586 -966 1654 -586
rect 1456 -1034 1654 -966
rect 870 -1160 1240 -1060
rect 1350 -1070 1440 -1060
rect 1350 -1150 1360 -1070
rect 1430 -1150 1440 -1070
rect 870 -1230 960 -1160
rect 1350 -1220 1440 -1150
rect 870 -1310 880 -1230
rect 950 -1310 960 -1230
rect 870 -1320 960 -1310
rect 1160 -1320 1440 -1220
rect 204 -1442 280 -1422
rect 204 -1498 214 -1442
rect 270 -1498 280 -1442
rect 204 -1524 280 -1498
rect 204 -1580 214 -1524
rect 270 -1580 280 -1524
rect 880 -1540 950 -1320
rect 1160 -1442 1240 -1320
rect 1160 -1480 1174 -1442
rect 1164 -1498 1174 -1480
rect 1230 -1498 1240 -1442
rect 1164 -1524 1240 -1498
rect 204 -1586 280 -1580
rect 340 -1646 1104 -1540
rect 1164 -1580 1174 -1524
rect 1230 -1580 1240 -1524
rect 1456 -1540 1524 -1034
rect 1746 -1126 1814 -926
rect 1164 -1586 1240 -1580
rect 1300 -1646 1524 -1540
rect 304 -1706 400 -1646
rect 112 -1882 180 -1868
rect 112 -2260 117 -1882
rect 174 -2260 180 -1882
rect 112 -2276 180 -2260
rect 304 -1882 372 -1706
rect 304 -2260 309 -1882
rect 366 -2260 372 -1882
rect 304 -2276 372 -2260
rect 496 -1882 564 -1646
rect 496 -2260 501 -1882
rect 558 -2260 564 -1882
rect 112 -2638 180 -2624
rect 112 -3336 117 -2638
rect 174 -3336 180 -2638
rect 112 -3352 180 -3336
rect 304 -2638 372 -2624
rect 304 -3336 309 -2638
rect 366 -3336 372 -2638
rect 304 -3352 372 -3336
rect 496 -2638 564 -2260
rect 496 -3336 501 -2638
rect 558 -3336 564 -2638
rect 496 -3352 564 -3336
rect 688 -1882 756 -1646
rect 688 -2260 693 -1882
rect 750 -2260 756 -1882
rect 688 -2638 756 -2260
rect 688 -3336 693 -2638
rect 750 -3336 756 -2638
rect 688 -3352 756 -3336
rect 880 -1882 948 -1646
rect 1044 -1706 1140 -1646
rect 880 -2260 885 -1882
rect 942 -2260 948 -1882
rect 880 -2638 948 -2260
rect 880 -3336 885 -2638
rect 942 -3336 948 -2638
rect 880 -3352 948 -3336
rect 1072 -1882 1140 -1706
rect 1072 -2260 1077 -1882
rect 1134 -2260 1140 -1882
rect 1072 -2416 1140 -2260
rect 1264 -1706 1360 -1646
rect 1264 -1882 1332 -1706
rect 1264 -2260 1269 -1882
rect 1326 -2210 1332 -1882
rect 1456 -1882 1524 -1646
rect 1326 -2260 1396 -2210
rect 1264 -2272 1396 -2260
rect 1072 -2426 1260 -2416
rect 1072 -2496 1176 -2426
rect 1250 -2496 1260 -2426
rect 1072 -2506 1260 -2496
rect 1072 -2638 1140 -2506
rect 1328 -2618 1396 -2272
rect 1072 -3336 1077 -2638
rect 1134 -3336 1140 -2638
rect 1072 -3352 1140 -3336
rect 1264 -2638 1396 -2618
rect 1264 -3336 1269 -2638
rect 1326 -2678 1396 -2638
rect 1456 -2260 1461 -1882
rect 1518 -2260 1524 -1882
rect 1456 -2638 1524 -2260
rect 1326 -3336 1332 -2678
rect 1264 -3352 1332 -3336
rect 1456 -3336 1461 -2638
rect 1518 -3336 1524 -2638
rect 1456 -3352 1524 -3336
rect 1648 -1194 1814 -1126
rect 1648 -1540 1716 -1194
rect 1930 -1442 2010 -100
rect 2070 -1000 2150 50
rect 2220 2 2292 120
rect 2892 104 2902 160
rect 2958 104 2968 160
rect 2892 78 2968 104
rect 2892 22 2902 78
rect 2958 22 2968 78
rect 2892 2 2968 22
rect 3084 160 3160 166
rect 3084 104 3094 160
rect 3150 104 3160 160
rect 3220 120 3984 226
rect 4044 160 4120 166
rect 3084 78 3160 104
rect 3084 22 3094 78
rect 3150 22 3160 78
rect 3084 2 3160 22
rect 2220 -1060 2290 2
rect 2600 -270 2690 -260
rect 2600 -350 2610 -270
rect 2680 -350 2690 -270
rect 2600 -360 2690 -350
rect 2210 -1070 2300 -1060
rect 2210 -1150 2220 -1070
rect 2290 -1150 2300 -1070
rect 2210 -1160 2300 -1150
rect 1930 -1480 1942 -1442
rect 1932 -1498 1942 -1480
rect 1998 -1480 2010 -1442
rect 1998 -1498 2008 -1480
rect 1932 -1524 2008 -1498
rect 1648 -1646 1872 -1540
rect 1932 -1580 1942 -1524
rect 1998 -1580 2008 -1524
rect 2610 -1540 2680 -360
rect 3760 -420 3830 120
rect 4044 104 4054 160
rect 4110 104 4120 160
rect 4180 120 4404 226
rect 4044 80 4120 104
rect 4040 78 4120 80
rect 4040 22 4054 78
rect 4110 22 4120 78
rect 4040 -360 4120 22
rect 3750 -430 3840 -420
rect 3750 -510 3760 -430
rect 3830 -510 3840 -430
rect 3750 -520 3840 -510
rect 3750 -910 3840 -900
rect 3750 -990 3760 -910
rect 3830 -990 3840 -910
rect 3750 -1000 3840 -990
rect 2892 -1442 2968 -1422
rect 2892 -1498 2902 -1442
rect 2958 -1498 2968 -1442
rect 2892 -1524 2968 -1498
rect 1932 -1586 2008 -1580
rect 2068 -1646 2832 -1540
rect 2892 -1580 2902 -1524
rect 2958 -1580 2968 -1524
rect 2892 -1586 2968 -1580
rect 3084 -1442 3160 -1422
rect 3084 -1498 3094 -1442
rect 3150 -1498 3160 -1442
rect 3084 -1524 3160 -1498
rect 3084 -1580 3094 -1524
rect 3150 -1580 3160 -1524
rect 3760 -1540 3830 -1000
rect 4040 -1442 4130 -740
rect 4040 -1470 4054 -1442
rect 4044 -1498 4054 -1470
rect 4110 -1470 4130 -1442
rect 4216 -1436 4284 -266
rect 4336 -1144 4404 120
rect 4528 1915 4596 1931
rect 4528 1217 4534 1915
rect 4591 1217 4596 1915
rect 4720 1915 4788 1931
rect 4720 1258 4726 1915
rect 4528 840 4596 1217
rect 4528 462 4534 840
rect 4591 462 4596 840
rect 4656 1217 4726 1258
rect 4783 1217 4788 1915
rect 4656 1198 4788 1217
rect 4912 1915 4980 1931
rect 4912 1217 4918 1915
rect 4975 1217 4980 1915
rect 4656 852 4724 1198
rect 4912 1086 4980 1217
rect 4792 1076 4980 1086
rect 4792 1006 4802 1076
rect 4876 1006 4980 1076
rect 4792 996 4980 1006
rect 4656 840 4788 852
rect 4656 790 4726 840
rect 4528 226 4596 462
rect 4720 462 4726 790
rect 4783 462 4788 840
rect 4720 286 4788 462
rect 4692 226 4788 286
rect 4912 840 4980 996
rect 4912 462 4918 840
rect 4975 462 4980 840
rect 4912 286 4980 462
rect 5104 1915 5172 1931
rect 5104 1217 5110 1915
rect 5167 1217 5172 1915
rect 5104 840 5172 1217
rect 5104 462 5110 840
rect 5167 462 5172 840
rect 4912 226 5008 286
rect 5104 226 5172 462
rect 5296 1915 5364 1931
rect 5296 1217 5302 1915
rect 5359 1217 5364 1915
rect 5296 840 5364 1217
rect 5296 462 5302 840
rect 5359 462 5364 840
rect 5296 226 5364 462
rect 5488 1915 5556 1931
rect 5488 1217 5494 1915
rect 5551 1217 5556 1915
rect 5488 840 5556 1217
rect 5680 1916 5748 1932
rect 5680 1218 5686 1916
rect 5743 1218 5748 1916
rect 5680 1110 5748 1218
rect 5872 1916 5940 1932
rect 5872 1218 5878 1916
rect 5935 1218 5940 1916
rect 5872 1110 5940 1218
rect 5488 462 5494 840
rect 5551 462 5556 840
rect 5488 226 5556 462
rect 5680 840 5748 856
rect 5680 462 5686 840
rect 5743 462 5748 840
rect 5680 286 5748 462
rect 5872 840 5940 856
rect 5872 462 5878 840
rect 5935 462 5940 840
rect 5872 448 5940 462
rect 5652 226 5748 286
rect 4528 120 4752 226
rect 4812 160 4888 166
rect 4528 -184 4596 120
rect 4812 104 4822 160
rect 4878 104 4888 160
rect 4948 120 5712 226
rect 5772 160 5848 166
rect 4812 78 4888 104
rect 4812 50 4822 78
rect 4810 22 4822 50
rect 4878 50 4888 78
rect 4878 22 4900 50
rect 4336 -1436 4404 -1420
rect 4110 -1498 4120 -1470
rect 4044 -1524 4120 -1498
rect 4216 -1504 4404 -1436
rect 3084 -1586 3160 -1580
rect 3220 -1646 3984 -1540
rect 4044 -1580 4054 -1524
rect 4110 -1580 4120 -1524
rect 4336 -1540 4404 -1504
rect 4044 -1586 4120 -1580
rect 4180 -1646 4404 -1540
rect 1648 -1882 1716 -1646
rect 1812 -1706 1908 -1646
rect 1648 -2260 1654 -1882
rect 1711 -2260 1716 -1882
rect 1840 -1882 1908 -1706
rect 1840 -2210 1846 -1882
rect 1648 -2637 1716 -2260
rect 1648 -3335 1654 -2637
rect 1711 -3335 1716 -2637
rect 1776 -2260 1846 -2210
rect 1903 -2260 1908 -1882
rect 1776 -2272 1908 -2260
rect 2032 -1706 2128 -1646
rect 2032 -1882 2100 -1706
rect 2032 -2260 2038 -1882
rect 2095 -2260 2100 -1882
rect 1776 -2618 1844 -2272
rect 2032 -2416 2100 -2260
rect 1912 -2426 2100 -2416
rect 1912 -2496 1922 -2426
rect 1996 -2496 2100 -2426
rect 1912 -2506 2100 -2496
rect 1776 -2637 1908 -2618
rect 1776 -2678 1846 -2637
rect 1648 -3351 1716 -3335
rect 1840 -3335 1846 -2678
rect 1903 -3335 1908 -2637
rect 1840 -3351 1908 -3335
rect 2032 -2637 2100 -2506
rect 2032 -3335 2038 -2637
rect 2095 -3335 2100 -2637
rect 2032 -3351 2100 -3335
rect 2224 -1882 2292 -1646
rect 2224 -2260 2230 -1882
rect 2287 -2260 2292 -1882
rect 2224 -2637 2292 -2260
rect 2224 -3335 2230 -2637
rect 2287 -3335 2292 -2637
rect 2224 -3351 2292 -3335
rect 2416 -1882 2484 -1646
rect 2416 -2260 2422 -1882
rect 2479 -2260 2484 -1882
rect 2416 -2637 2484 -2260
rect 2416 -3335 2422 -2637
rect 2479 -3335 2484 -2637
rect 2416 -3351 2484 -3335
rect 2608 -1882 2676 -1646
rect 2772 -1706 2868 -1646
rect 2608 -2260 2614 -1882
rect 2671 -2260 2676 -1882
rect 2608 -2637 2676 -2260
rect 2800 -1882 2868 -1706
rect 3184 -1706 3280 -1646
rect 2800 -2260 2806 -1882
rect 2863 -2260 2868 -1882
rect 2800 -2276 2868 -2260
rect 2992 -1882 3060 -1868
rect 2992 -2260 2997 -1882
rect 3055 -2260 3060 -1882
rect 2992 -2276 3060 -2260
rect 3184 -1882 3252 -1706
rect 3184 -2260 3189 -1882
rect 3246 -2260 3252 -1882
rect 3184 -2276 3252 -2260
rect 3376 -1882 3444 -1646
rect 3376 -2260 3381 -1882
rect 3438 -2260 3444 -1882
rect 2608 -3335 2614 -2637
rect 2671 -3335 2676 -2637
rect 2608 -3351 2676 -3335
rect 2800 -2638 2868 -2530
rect 2800 -3336 2806 -2638
rect 2863 -3336 2868 -2638
rect 2800 -3352 2868 -3336
rect 2992 -2638 3060 -2530
rect 2992 -3336 2997 -2638
rect 3055 -3336 3060 -2638
rect 2992 -3352 3060 -3336
rect 3184 -2638 3252 -2624
rect 3184 -3336 3189 -2638
rect 3246 -3336 3252 -2638
rect 3184 -3352 3252 -3336
rect 3376 -2638 3444 -2260
rect 3376 -3336 3381 -2638
rect 3438 -3336 3444 -2638
rect 3376 -3352 3444 -3336
rect 3568 -1882 3636 -1646
rect 3568 -2260 3573 -1882
rect 3630 -2260 3636 -1882
rect 3568 -2638 3636 -2260
rect 3568 -3336 3573 -2638
rect 3630 -3336 3636 -2638
rect 3568 -3352 3636 -3336
rect 3760 -1882 3828 -1646
rect 3924 -1706 4020 -1646
rect 3760 -2260 3765 -1882
rect 3822 -2260 3828 -1882
rect 3760 -2638 3828 -2260
rect 3760 -3336 3765 -2638
rect 3822 -3336 3828 -2638
rect 3760 -3352 3828 -3336
rect 3952 -1882 4020 -1706
rect 3952 -2260 3957 -1882
rect 4014 -2260 4020 -1882
rect 3952 -2416 4020 -2260
rect 4144 -1706 4240 -1646
rect 4144 -1882 4212 -1706
rect 4144 -2260 4149 -1882
rect 4206 -2210 4212 -1882
rect 4336 -1882 4404 -1646
rect 4206 -2260 4276 -2210
rect 4144 -2272 4276 -2260
rect 3952 -2426 4140 -2416
rect 3952 -2496 4056 -2426
rect 4130 -2496 4140 -2426
rect 3952 -2506 4140 -2496
rect 3952 -2638 4020 -2506
rect 4208 -2618 4276 -2272
rect 3952 -3336 3957 -2638
rect 4014 -3336 4020 -2638
rect 3952 -3352 4020 -3336
rect 4144 -2638 4276 -2618
rect 4144 -3336 4149 -2638
rect 4206 -2678 4276 -2638
rect 4336 -2260 4341 -1882
rect 4398 -2260 4404 -1882
rect 4336 -2638 4404 -2260
rect 4206 -3336 4212 -2678
rect 4144 -3352 4212 -3336
rect 4336 -3336 4341 -2638
rect 4398 -3336 4404 -2638
rect 4336 -3352 4404 -3336
rect 4528 -1540 4596 -586
rect 4810 -680 4900 22
rect 4960 -1360 5030 -430
rect 5100 -740 5170 120
rect 5772 104 5782 160
rect 5838 104 5848 160
rect 5772 78 5848 104
rect 5772 22 5782 78
rect 5838 22 5848 78
rect 5772 2 5848 22
rect 5480 -590 5570 -580
rect 5480 -670 5490 -590
rect 5560 -670 5570 -590
rect 5480 -680 5570 -670
rect 5090 -750 5180 -740
rect 5090 -830 5100 -750
rect 5170 -830 5180 -750
rect 5090 -840 5180 -830
rect 4812 -1442 4888 -1422
rect 4812 -1498 4822 -1442
rect 4878 -1498 4888 -1442
rect 4812 -1524 4888 -1498
rect 4528 -1646 4752 -1540
rect 4812 -1580 4822 -1524
rect 4878 -1580 4888 -1524
rect 5490 -1540 5560 -680
rect 5772 -1442 5848 -1422
rect 5772 -1498 5782 -1442
rect 5838 -1498 5848 -1442
rect 5772 -1524 5848 -1498
rect 4812 -1586 4888 -1580
rect 4948 -1646 5712 -1540
rect 5772 -1580 5782 -1524
rect 5838 -1580 5848 -1524
rect 5772 -1586 5848 -1580
rect 4528 -1882 4596 -1646
rect 4692 -1706 4788 -1646
rect 4528 -2260 4534 -1882
rect 4591 -2260 4596 -1882
rect 4720 -1882 4788 -1706
rect 4720 -2210 4726 -1882
rect 4528 -2637 4596 -2260
rect 4528 -3335 4534 -2637
rect 4591 -3335 4596 -2637
rect 4656 -2260 4726 -2210
rect 4783 -2260 4788 -1882
rect 4656 -2272 4788 -2260
rect 4912 -1706 5008 -1646
rect 4912 -1882 4980 -1706
rect 4912 -2260 4918 -1882
rect 4975 -2260 4980 -1882
rect 4656 -2618 4724 -2272
rect 4912 -2416 4980 -2260
rect 4792 -2426 4980 -2416
rect 4792 -2496 4802 -2426
rect 4876 -2496 4980 -2426
rect 4792 -2506 4980 -2496
rect 4656 -2637 4788 -2618
rect 4656 -2678 4726 -2637
rect 4528 -3351 4596 -3335
rect 4720 -3335 4726 -2678
rect 4783 -3335 4788 -2637
rect 4720 -3351 4788 -3335
rect 4912 -2637 4980 -2506
rect 4912 -3335 4918 -2637
rect 4975 -3335 4980 -2637
rect 4912 -3351 4980 -3335
rect 5104 -1882 5172 -1646
rect 5104 -2260 5110 -1882
rect 5167 -2260 5172 -1882
rect 5104 -2637 5172 -2260
rect 5104 -3335 5110 -2637
rect 5167 -3335 5172 -2637
rect 5104 -3351 5172 -3335
rect 5296 -1882 5364 -1646
rect 5296 -2260 5302 -1882
rect 5359 -2260 5364 -1882
rect 5296 -2637 5364 -2260
rect 5296 -3335 5302 -2637
rect 5359 -3335 5364 -2637
rect 5296 -3351 5364 -3335
rect 5488 -1882 5556 -1646
rect 5652 -1706 5748 -1646
rect 5488 -2260 5494 -1882
rect 5551 -2260 5556 -1882
rect 5488 -2637 5556 -2260
rect 5680 -1882 5748 -1706
rect 5680 -2260 5686 -1882
rect 5743 -2260 5748 -1882
rect 5680 -2276 5748 -2260
rect 5872 -1882 5940 -1868
rect 5872 -2260 5878 -1882
rect 5935 -2260 5940 -1882
rect 5872 -2276 5940 -2260
rect 5488 -3335 5494 -2637
rect 5551 -3335 5556 -2637
rect 5488 -3351 5556 -3335
rect 5680 -2638 5748 -2530
rect 5680 -3336 5686 -2638
rect 5743 -3336 5748 -2638
rect 5680 -3352 5748 -3336
rect 5872 -2638 5940 -2530
rect 5872 -3336 5878 -2638
rect 5935 -3336 5940 -2638
rect 5872 -3352 5940 -3336
<< via3 >>
rect 880 -190 950 -110
rect 1360 -1150 1430 -1070
rect 880 -1310 950 -1230
rect 2610 -350 2680 -270
rect 2220 -1150 2290 -1070
rect 3760 -510 3830 -430
rect 3760 -990 3830 -910
rect 5490 -670 5560 -590
rect 5100 -830 5170 -750
<< metal4 >>
rect 100 -110 6000 -100
rect 100 -190 880 -110
rect 950 -190 6000 -110
rect 100 -200 6000 -190
rect 100 -270 6000 -260
rect 100 -350 2610 -270
rect 2680 -350 6000 -270
rect 100 -360 6000 -350
rect 100 -430 6000 -420
rect 100 -510 3760 -430
rect 3830 -510 6000 -430
rect 100 -520 6000 -510
rect 100 -590 6000 -580
rect 100 -670 5490 -590
rect 5560 -670 6000 -590
rect 100 -680 6000 -670
rect 100 -750 6000 -740
rect 100 -830 5100 -750
rect 5170 -830 6000 -750
rect 100 -840 6000 -830
rect 100 -910 6000 -900
rect 100 -990 3760 -910
rect 3830 -990 6000 -910
rect 100 -1000 6000 -990
rect 100 -1070 6000 -1060
rect 100 -1150 1360 -1070
rect 1430 -1150 2220 -1070
rect 2290 -1150 6000 -1070
rect 100 -1160 6000 -1150
rect 100 -1230 6000 -1220
rect 100 -1310 880 -1230
rect 950 -1310 6000 -1230
rect 100 -1320 6000 -1310
<< comment >>
rect 74 1994 88 2024
rect 266 1994 280 2024
rect 2892 1994 2906 2024
rect 2954 1994 2968 2024
rect 3084 1994 3098 2024
rect 3146 1994 3160 2024
rect 5772 1994 5786 2024
rect 5964 1994 5978 2024
rect -940 660 -910 670
rect -940 650 -930 660
rect -920 650 -910 660
rect -940 640 -910 650
rect -920 630 -910 640
rect -940 620 -910 630
rect -900 660 -870 670
rect -860 660 -830 670
rect -900 650 -890 660
rect -880 650 -870 660
rect -840 650 -830 660
rect -820 660 -790 670
rect -780 660 -750 670
rect -820 650 -810 660
rect -780 650 -770 660
rect -740 650 -730 670
rect -720 650 -710 670
rect -700 660 -670 670
rect -660 660 -630 670
rect -610 660 -600 670
rect -680 650 -670 660
rect -640 650 -630 660
rect -620 650 -600 660
rect -900 640 -870 650
rect -900 630 -890 640
rect -880 630 -870 640
rect -900 620 -870 630
rect -850 620 -840 650
rect -820 640 -790 650
rect -780 640 -750 650
rect -740 640 -710 650
rect -700 640 -670 650
rect -820 630 -810 640
rect -800 630 -790 640
rect -760 630 -750 640
rect -820 620 -790 630
rect -780 620 -750 630
rect -720 620 -710 640
rect -680 630 -670 640
rect -700 620 -670 630
rect -660 640 -630 650
rect -660 630 -650 640
rect -610 630 -600 650
rect -580 660 -550 670
rect -580 630 -570 660
rect -560 630 -550 660
rect -660 620 -630 630
rect -620 620 -590 630
rect -580 620 -550 630
rect 100 -160 130 -150
rect 100 -190 110 -160
rect 120 -190 130 -160
rect 100 -200 130 -190
rect 100 -330 110 -310
rect 120 -330 130 -310
rect 100 -340 130 -330
rect 140 -320 170 -310
rect 140 -330 150 -320
rect 140 -340 170 -330
rect 120 -360 130 -340
rect 160 -350 170 -340
rect 140 -360 170 -350
rect 100 -480 130 -470
rect 100 -490 110 -480
rect 120 -490 130 -480
rect 100 -500 130 -490
rect 120 -510 130 -500
rect 100 -520 130 -510
rect 140 -480 170 -470
rect 140 -510 150 -480
rect 160 -510 170 -480
rect 140 -520 170 -510
rect 110 -640 120 -630
rect 140 -640 170 -630
rect 100 -650 120 -640
rect 160 -650 170 -640
rect 110 -670 120 -650
rect 140 -660 170 -650
rect 180 -640 210 -630
rect 180 -650 190 -640
rect 180 -660 210 -650
rect 160 -670 170 -660
rect 200 -670 210 -660
rect 100 -680 130 -670
rect 140 -680 170 -670
rect 180 -680 210 -670
rect 110 -800 120 -790
rect 100 -810 120 -800
rect 110 -830 120 -810
rect 140 -800 170 -790
rect 140 -810 150 -800
rect 160 -810 170 -800
rect 140 -820 170 -810
rect 140 -830 150 -820
rect 160 -830 170 -820
rect 100 -840 130 -830
rect 140 -840 170 -830
rect 180 -800 210 -790
rect 180 -830 190 -800
rect 200 -830 210 -800
rect 180 -840 210 -830
rect 100 -960 130 -950
rect 140 -960 170 -950
rect 120 -970 130 -960
rect 160 -970 170 -960
rect 100 -980 130 -970
rect 140 -980 170 -970
rect 180 -960 210 -950
rect 180 -970 190 -960
rect 180 -980 210 -970
rect 100 -990 110 -980
rect 140 -990 150 -980
rect 200 -990 210 -980
rect 100 -1000 130 -990
rect 140 -1000 170 -990
rect 180 -1000 210 -990
rect 100 -1120 130 -1110
rect 140 -1120 170 -1110
rect 120 -1130 130 -1120
rect 160 -1130 170 -1120
rect 180 -1120 210 -1110
rect 100 -1140 130 -1130
rect 100 -1150 110 -1140
rect 100 -1160 130 -1150
rect 150 -1160 160 -1130
rect 180 -1150 190 -1120
rect 200 -1150 210 -1120
rect 180 -1160 210 -1150
rect 100 -1280 130 -1270
rect 150 -1280 160 -1270
rect 120 -1290 130 -1280
rect 140 -1290 160 -1280
rect 100 -1300 130 -1290
rect 120 -1310 130 -1300
rect 150 -1310 160 -1290
rect 180 -1280 210 -1270
rect 180 -1290 190 -1280
rect 180 -1300 210 -1290
rect 200 -1310 210 -1300
rect 100 -1320 130 -1310
rect 140 -1320 170 -1310
rect 180 -1320 210 -1310
rect 74 -3444 88 -3414
rect 266 -3444 280 -3414
rect 2892 -3444 2906 -3414
rect 2954 -3444 2968 -3414
rect 3084 -3444 3098 -3414
rect 3146 -3444 3160 -3414
rect 5772 -3444 5786 -3414
rect 5964 -3444 5978 -3414
<< end >>
