magic
tech sky130A
magscale 1 2
timestamp 1671336542
<< metal1 >>
rect -4320 -7120 -4280 -6920
rect -4200 -7120 -4160 -6920
<< metal2 >>
rect -2600 0 2000 100
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 1860 -3140 2060 -3100
rect -1060 -4320 -680 -4300
rect -1060 -4480 -1040 -4320
rect -700 -4480 -680 -4320
rect -1060 -4500 -680 -4480
rect -2840 -6200 -2340 -5800
rect -2840 -6500 -1600 -6200
rect -2840 -6700 -2340 -6500
rect -3760 -7140 -3680 -6940
rect -3320 -7000 -1600 -6700
rect 1600 -7000 2000 -5800
rect -3000 -7100 -1200 -7000
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via2 >>
rect -2500 -500 1900 0
rect -1040 -4480 -700 -4320
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< metal3 >>
rect -2600 0 2000 100
rect -7600 -7100 -4800 -200
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect -660 -4200 -620 -4180
rect 120 -4200 160 -4180
rect -1400 -4320 -680 -4300
rect -1400 -4480 -1040 -4320
rect -700 -4480 -680 -4320
rect -1400 -4500 -680 -4480
rect -3600 -5700 -2800 -5600
rect -1400 -5700 -1100 -4500
rect -3600 -5800 -1100 -5700
rect -3000 -6000 -1100 -5800
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 -1200 -7000
rect -4900 -7600 -4600 -7300
rect -4900 -7700 -4800 -7600
rect -7600 -7800 -4800 -7700
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via3 >>
rect -2500 -500 1900 0
rect -7500 -7700 -4900 -7100
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< mimcap >>
rect -7500 -340 -4900 -300
rect -7500 -6660 -7460 -340
rect -4940 -6660 -4900 -340
rect -7500 -6700 -4900 -6660
<< mimcapcontact >>
rect -7460 -6660 -4940 -340
<< metal4 >>
rect -7400 100 2000 600
rect -7400 -200 -5000 100
rect -2600 0 2000 100
rect -7600 -340 -4800 -200
rect -7600 -6660 -7460 -340
rect -4940 -6660 -4800 -340
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect -7600 -6800 -4800 -6660
rect -7600 -7100 -4800 -7000
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 2000 -7000
rect -3000 -7300 -2900 -7100
rect -4900 -7700 -2900 -7300
rect -1300 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect -7600 -7800 2000 -7700
<< via4 >>
rect -7500 -7700 -4900 -7100
<< mimcap2 >>
rect -7500 -340 -4900 -300
rect -7500 -6660 -7460 -340
rect -4940 -6660 -4900 -340
rect -7500 -6700 -4900 -6660
<< mimcap2contact >>
rect -7460 -6660 -4940 -340
<< metal5 >>
rect -7600 -340 -4800 -200
rect -7600 -6660 -7460 -340
rect -4940 -6660 -4800 -340
rect -7600 -7100 -4800 -6660
rect -7600 -7700 -7500 -7100
rect -4900 -7700 -4800 -7100
rect -7600 -7800 -4800 -7700
use cmota_1_flat_1  cmota_1_flat_1_0
timestamp 1671334909
transform 1 0 -2836 0 1 -3200
box -164 -3800 5363 2800
use gated_iref  gated_iref_0
timestamp 1671335613
transform 0 1 -4300 1 0 -7948
box 948 -100 7800 1200
<< labels >>
rlabel metal4 -3840 -7800 -3660 -7300 1 VLO
rlabel metal2 -3760 -7140 -3680 -7060 1 VREF
rlabel metal1 -4200 -7120 -4160 -7080 1 S
rlabel metal1 -4320 -7120 -4280 -7080 1 SBAR
rlabel metal4 -4220 320 -3840 600 1 VHI
rlabel metal3 -660 -4200 -620 -4180 1 VIN
rlabel metal3 120 -4200 160 -4180 1 VIP
rlabel metal2 1860 -3140 2060 -3100 1 VOP
<< end >>
