magic
tech sky130A
timestamp 1672120492
<< metal2 >>
rect 390 12760 530 12770
rect 390 12640 400 12760
rect 520 12640 530 12760
rect 390 12630 530 12640
<< via2 >>
rect 400 12640 520 12760
<< metal3 >>
rect 390 12765 865 12770
rect 390 12635 400 12765
rect 860 12635 865 12765
rect 390 12630 865 12635
rect 395 11975 865 11980
rect 395 11835 400 11975
rect 860 11835 865 11975
rect 395 11830 865 11835
<< via3 >>
rect 400 12760 860 12765
rect 400 12640 520 12760
rect 520 12640 860 12760
rect 400 12635 860 12640
rect 400 11835 860 11975
<< metal4 >>
rect -3830 12910 -3430 14750
rect -3830 12750 -3810 12910
rect -3450 12750 -3430 12910
rect -3830 600 -3430 12750
rect -3330 12540 -2930 14750
rect -3330 12380 -3310 12540
rect -2950 12380 -2930 12540
rect -3330 600 -2930 12380
rect -2830 12180 -2430 14750
rect -2830 12020 -2810 12180
rect -2450 12020 -2430 12180
rect -2830 600 -2430 12020
rect -2330 11050 -1680 14750
rect -2330 10450 -2280 11050
rect -1730 10450 -1680 11050
rect -2330 8900 -1680 10450
rect -2330 8000 -2280 8900
rect -1730 8000 -1680 8900
rect -2330 6900 -1680 8000
rect -2330 6000 -2280 6900
rect -1730 6000 -1680 6900
rect -2330 4900 -1680 6000
rect -2330 4000 -2280 4900
rect -1730 4000 -1680 4900
rect -2330 2900 -1680 4000
rect -2330 2000 -2280 2900
rect -1730 2000 -1680 2900
rect -2330 600 -1680 2000
rect -1580 12950 -930 14750
rect -730 12950 -80 14750
rect -1580 11950 -80 12950
rect 395 12765 865 12770
rect 395 12635 400 12765
rect 860 12635 865 12765
rect 395 12630 865 12635
rect -40 12540 130 12560
rect -40 12380 -20 12540
rect 110 12380 130 12540
rect -40 12230 805 12380
rect -1580 11750 -930 11950
rect -1580 11350 -1530 11750
rect -980 11350 -930 11750
rect -1580 10950 -930 11350
rect -730 11750 -80 11950
rect 395 11975 865 11980
rect 395 11835 400 11975
rect 860 11835 865 11975
rect 395 11830 865 11835
rect -730 11350 -680 11750
rect -130 11350 -80 11750
rect -730 10950 -80 11350
rect -1580 9950 -80 10950
rect -1580 8950 -930 9950
rect -730 8950 -80 9950
rect -1580 7950 -80 8950
rect -1580 6950 -930 7950
rect -730 6950 -80 7950
rect -1580 5950 -80 6950
rect -1580 4950 -930 5950
rect -730 4950 -80 5950
rect -1580 3950 -80 4950
rect -1580 2950 -930 3950
rect -730 2950 -80 3950
rect -1580 1950 -80 2950
rect -1580 600 -930 1950
rect -730 600 -80 1950
<< via4 >>
rect -3810 12750 -3450 12910
rect -3310 12380 -2950 12540
rect -2810 12020 -2450 12180
rect -2280 10450 -1730 11050
rect -2280 8000 -1730 8900
rect -2280 6000 -1730 6900
rect -2280 4000 -1730 4900
rect -2280 2000 -1730 2900
rect -20 12380 110 12540
rect -1530 11350 -980 11750
rect -680 11350 -130 11750
<< mimcap2 >>
rect -1560 10370 -950 10380
rect -1560 1880 -1550 10370
rect -960 1880 -950 10370
rect -1560 1870 -950 1880
rect -710 10370 -100 10380
rect -710 1880 -700 10370
rect -110 1880 -100 10370
rect -710 1870 -100 1880
<< mimcap2contact >>
rect -1550 1880 -960 10370
rect -700 1880 -110 10370
<< metal5 >>
rect -3830 12910 485 12930
rect -3830 12750 -3810 12910
rect -3450 12750 485 12910
rect -3830 12730 485 12750
rect 285 12600 485 12730
rect -3330 12540 125 12560
rect -3330 12380 -3310 12540
rect -2950 12380 -20 12540
rect 110 12380 125 12540
rect 285 12400 900 12600
rect -3330 12360 125 12380
rect -2830 12180 855 12200
rect -2830 12020 -2810 12180
rect -2450 12020 855 12180
rect -2830 12000 855 12020
rect -1580 11750 650 11800
rect -1580 11350 -1530 11750
rect -980 11350 -680 11750
rect -130 11350 650 11750
rect -1580 11300 650 11350
rect -2330 11050 850 11100
rect -2330 10450 -2280 11050
rect -1730 10600 850 11050
rect -1730 10450 -730 10600
rect -2330 10400 -730 10450
rect -1580 10370 -80 10400
rect -1580 8950 -1550 10370
rect -2330 8900 -1550 8950
rect -2330 8000 -2280 8900
rect -1730 8000 -1550 8900
rect -2330 7950 -1550 8000
rect -1580 6950 -1550 7950
rect -2330 6900 -1550 6950
rect -2330 6000 -2280 6900
rect -1730 6000 -1550 6900
rect -2330 5950 -1550 6000
rect -1580 4950 -1550 5950
rect -2330 4900 -1550 4950
rect -2330 4000 -2280 4900
rect -1730 4000 -1550 4900
rect -2330 3950 -1550 4000
rect -1580 2950 -1550 3950
rect -2330 2900 -1550 2950
rect -2330 2000 -2280 2900
rect -1730 2000 -1550 2900
rect -2330 1950 -1550 2000
rect -1580 1880 -1550 1950
rect -960 9950 -700 10370
rect -960 8950 -930 9950
rect -730 8950 -700 9950
rect -960 7950 -700 8950
rect -960 6950 -930 7950
rect -730 6950 -700 7950
rect -960 5950 -700 6950
rect -960 4950 -930 5950
rect -730 4950 -700 5950
rect -960 3950 -700 4950
rect -960 2950 -930 3950
rect -730 2950 -700 3950
rect -960 1950 -700 2950
rect -960 1880 -930 1950
rect -1580 1850 -930 1880
rect -730 1880 -700 1950
rect -110 1880 -80 10370
rect -730 1850 -80 1880
<< end >>
