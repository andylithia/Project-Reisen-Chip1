magic
tech sky130A
magscale 1 2
timestamp 1672205966
<< pwell >>
rect 1066 781 1734 860
rect 1066 772 1308 781
rect 1414 772 1734 781
rect 1066 744 1734 772
rect 1066 698 1730 744
rect 1066 -60 1734 698
<< nmos >>
rect 1682 150 1712 650
rect 1778 150 1808 650
rect 1874 150 1904 650
rect 1970 150 2000 650
rect 2066 150 2096 650
<< ndiff >>
rect 1620 638 1682 650
rect 1620 162 1632 638
rect 1666 162 1682 638
rect 1620 150 1682 162
rect 1712 638 1778 650
rect 1712 162 1728 638
rect 1762 162 1778 638
rect 1712 150 1778 162
rect 1808 638 1874 650
rect 1808 162 1824 638
rect 1858 162 1874 638
rect 1808 150 1874 162
rect 1904 638 1970 650
rect 1904 162 1920 638
rect 1954 162 1970 638
rect 1904 150 1970 162
rect 2000 638 2066 650
rect 2000 162 2016 638
rect 2050 162 2066 638
rect 2000 150 2066 162
rect 2096 638 2158 650
rect 2096 162 2112 638
rect 2146 162 2158 638
rect 2096 150 2158 162
<< ndiffc >>
rect 1632 162 1666 638
rect 1728 162 1762 638
rect 1824 162 1858 638
rect 1920 162 1954 638
rect 2016 162 2050 638
rect 2112 162 2146 638
<< psubdiff >>
rect 1102 790 1218 824
rect 2164 790 2260 824
rect 1102 728 1136 790
rect 2226 728 2260 790
rect 1102 10 1136 72
rect 2226 10 2260 72
rect 1102 -24 1218 10
rect 2164 -24 2260 10
<< psubdiffcont >>
rect 1218 790 2164 824
rect 1102 72 1136 728
rect 2226 72 2260 728
rect 1218 -24 2164 10
<< poly >>
rect 1682 650 1712 676
rect 1778 650 1808 676
rect 1874 650 1904 676
rect 1970 650 2000 676
rect 2066 650 2096 676
rect 1682 128 1712 150
rect 1778 128 1808 150
rect 1874 132 1904 150
rect 1682 112 1808 128
rect 1682 78 1758 112
rect 1792 78 1808 112
rect 1682 62 1808 78
rect 1857 105 1920 132
rect 1857 71 1872 105
rect 1906 71 1920 105
rect 1857 44 1920 71
rect 1970 128 2000 150
rect 2066 128 2096 150
rect 1970 112 2096 128
rect 1970 78 2046 112
rect 2080 78 2096 112
rect 1970 62 2096 78
<< polycont >>
rect 1758 78 1792 112
rect 1872 71 1906 105
rect 2046 78 2080 112
<< xpolycontact >>
rect 1278 106 1348 538
rect 1444 106 1514 538
<< xpolyres >>
rect 1278 604 1514 674
rect 1278 538 1348 604
rect 1444 538 1514 604
<< locali >>
rect 1068 960 2028 980
rect 1068 900 1088 960
rect 2008 900 2028 960
rect 1068 866 2028 900
rect 1068 858 2124 866
rect 1068 824 2294 858
rect 1068 790 1218 824
rect 2164 790 2294 824
rect 1068 728 1136 790
rect 1068 72 1102 728
rect 1632 638 1666 654
rect 1068 10 1136 72
rect 1278 90 1287 106
rect 1340 90 1348 106
rect 1278 67 1348 90
rect 1632 118 1666 162
rect 1728 638 1762 654
rect 1728 146 1762 162
rect 1824 638 1858 654
rect 1824 146 1858 162
rect 1920 638 1954 790
rect 1920 146 1954 162
rect 2016 638 2050 654
rect 2016 146 2050 162
rect 2112 638 2146 790
rect 2112 146 2146 162
rect 2226 728 2294 790
rect 1514 106 1666 118
rect 1444 67 1666 106
rect 1742 78 1758 112
rect 1792 78 1808 112
rect 1856 71 1872 105
rect 1906 71 1922 105
rect 2030 78 2046 112
rect 2080 78 2096 112
rect 2260 72 2294 728
rect 1869 10 1909 71
rect 2226 10 2294 72
rect 1068 -24 1218 10
rect 2164 -24 2294 10
rect 1068 -58 2294 -24
rect 1080 -240 1220 -58
rect 1080 -560 1280 -240
<< viali >>
rect 1088 900 2008 960
rect 1287 106 1340 522
rect 1287 90 1340 106
rect 1632 162 1666 638
rect 1728 162 1762 638
rect 1824 162 1858 638
rect 1920 162 1954 638
rect 2016 162 2050 638
rect 2112 162 2146 638
rect 1758 78 1792 112
rect 2046 78 2080 112
<< metal1 >>
rect 1068 1100 2028 1120
rect 1068 900 1088 1100
rect 2008 900 2028 1100
rect 1068 880 2028 900
rect 1626 718 1864 758
rect 1626 638 1672 718
rect 1278 522 1348 538
rect 1278 519 1287 522
rect 1340 519 1348 522
rect 1626 162 1632 638
rect 1666 162 1672 638
rect 1626 150 1672 162
rect 1719 638 1771 650
rect 1719 635 1728 638
rect 1762 635 1771 638
rect 1719 162 1728 166
rect 1762 162 1771 166
rect 1719 150 1771 162
rect 1818 638 1864 718
rect 1818 162 1824 638
rect 1858 162 1864 638
rect 1818 150 1864 162
rect 1914 638 1960 650
rect 1914 162 1920 638
rect 1954 162 1960 638
rect 1914 150 1960 162
rect 2007 638 2059 650
rect 2007 635 2016 638
rect 2050 635 2059 638
rect 2007 162 2016 166
rect 2050 162 2059 166
rect 2007 149 2059 162
rect 2106 638 2152 650
rect 2106 162 2112 638
rect 2146 162 2152 638
rect 2106 150 2152 162
rect 1278 67 1348 90
rect 1728 66 1739 118
rect 1791 112 1808 118
rect 1792 78 1808 112
rect 1791 66 1808 78
rect 2016 112 2096 118
rect 2016 78 2046 112
rect 2080 78 2096 112
rect 2016 72 2096 78
rect 2016 33 2050 72
rect 1038 -1 2050 33
rect 1039 -63 1740 -29
rect 1728 -81 1740 -63
rect 1792 -63 1809 -29
rect 1792 -81 1808 -63
<< via1 >>
rect 1088 960 2008 1100
rect 1088 900 2008 960
rect 1278 90 1287 519
rect 1287 90 1340 519
rect 1340 90 1348 519
rect 1719 166 1728 635
rect 1728 166 1762 635
rect 1762 166 1771 635
rect 2007 166 2016 635
rect 2016 166 2050 635
rect 2050 166 2059 635
rect 1739 112 1791 118
rect 1739 78 1758 112
rect 1758 78 1791 112
rect 1739 66 1791 78
rect 1740 -81 1792 -29
<< metal2 >>
rect 1068 1100 2028 1120
rect 1068 900 1088 1100
rect 2008 900 2028 1100
rect 1068 880 2028 900
rect 940 200 1060 360
rect 980 -2340 1060 200
rect 1100 -240 1220 880
rect 1719 640 2240 650
rect 1719 635 2060 640
rect 1278 519 1348 538
rect 1260 90 1278 300
rect 1771 580 2007 635
rect 1719 150 1771 166
rect 2059 500 2060 635
rect 2230 500 2240 640
rect 2059 490 2240 500
rect 2007 149 2059 166
rect 1260 67 1348 90
rect 1260 -120 1340 67
rect 1728 66 1739 118
rect 1791 66 1808 118
rect 1740 -29 1792 66
rect 1728 -81 1740 -29
rect 1792 -81 1808 -29
rect 1260 -200 2690 -120
rect 1360 -220 2690 -200
rect 1100 -560 1240 -240
rect 2590 -710 2690 -220
rect 2580 -2340 2720 -2280
rect 980 -2420 2720 -2340
<< via2 >>
rect 1088 900 2008 1100
rect 2060 500 2230 640
<< metal3 >>
rect 1068 1180 2028 1200
rect 1068 900 1088 1180
rect 2008 900 2028 1180
rect 1068 880 2028 900
rect 2200 800 7800 1200
rect 1200 770 7800 800
rect 1200 -70 1230 770
rect 1880 640 7800 770
rect 1880 500 2060 640
rect 2230 500 7800 640
rect 1880 -70 7800 500
rect 1200 -100 7800 -70
<< via3 >>
rect 1088 1100 2008 1180
rect 1088 980 2008 1100
rect 1230 -70 1880 770
<< mimcap >>
rect 2250 1150 7770 1170
rect 2250 -50 2270 1150
rect 7750 -50 7770 1150
rect 2250 -70 7770 -50
<< mimcapcontact >>
rect 2270 -50 7750 1150
<< metal4 >>
rect 1068 1180 7800 1200
rect 1068 980 1088 1180
rect 2008 1150 7800 1180
rect 2008 980 2270 1150
rect 1068 960 2270 980
rect 1200 770 1910 800
rect 1200 -70 1230 770
rect 1880 -70 1910 770
rect 1200 -100 1910 -70
rect 2200 -50 2270 960
rect 7750 -50 7800 1150
rect 2200 -100 7800 -50
<< via4 >>
rect 1230 -70 1880 770
<< mimcap2 >>
rect 2250 1150 7770 1170
rect 2250 -50 2270 1150
rect 7750 -50 7770 1150
rect 2250 -70 7770 -50
<< mimcap2contact >>
rect 2270 -50 7750 1150
<< metal5 >>
rect 2200 1150 7800 1200
rect 2200 800 2270 1150
rect 1200 770 2270 800
rect 1200 -70 1230 770
rect 1880 -50 2270 770
rect 7750 -50 7800 1150
rect 1880 -70 7800 -50
rect 1200 -100 7800 -70
<< comment >>
rect 7800 1200 7820 1220
rect 2180 940 2200 960
rect 1180 800 1200 820
rect 2276 800 2296 820
rect 1824 139 1825 145
rect 1180 -120 1200 -100
rect 7800 -120 7820 -100
use imirror2  imirror2_0
timestamp 1672168347
transform 0 1 1260 1 0 -6240
box 3897 -20 6064 3880
<< labels >>
rlabel locali 1068 862 1324 880 1 VSUB
rlabel metal1 1040 0 1064 32 1 SBAR
rlabel metal1 1040 -62 1064 -30 1 S
<< end >>
