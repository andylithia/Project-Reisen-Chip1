magic
tech sky130A
timestamp 1672298248
<< metal1 >>
rect 3000 9378 7000 9500
rect 3000 9352 3307 9378
rect 3333 9352 3467 9378
rect 3493 9352 3627 9378
rect 3653 9352 3787 9378
rect 3813 9352 3947 9378
rect 3973 9352 4107 9378
rect 4133 9352 4267 9378
rect 4293 9352 4427 9378
rect 4453 9352 4587 9378
rect 4613 9352 4747 9378
rect 4773 9352 4907 9378
rect 4933 9352 5067 9378
rect 5093 9352 5227 9378
rect 5253 9352 5387 9378
rect 5413 9352 5547 9378
rect 5573 9352 5707 9378
rect 5733 9352 5867 9378
rect 5893 9352 6027 9378
rect 6053 9352 6187 9378
rect 6213 9352 6347 9378
rect 6373 9352 6507 9378
rect 6533 9352 6667 9378
rect 6693 9352 7000 9378
rect 3000 9273 7000 9352
rect 3000 9247 3119 9273
rect 3145 9247 6852 9273
rect 6878 9247 7000 9273
rect 3000 9230 7000 9247
rect 3000 9113 3270 9230
rect 3000 9087 3119 9113
rect 3145 9087 3270 9113
rect 3000 8953 3270 9087
rect 3000 8927 3119 8953
rect 3145 8927 3270 8953
rect 3000 8793 3270 8927
rect 3000 8767 3119 8793
rect 3145 8767 3270 8793
rect 3000 8633 3270 8767
rect 3000 8607 3119 8633
rect 3145 8607 3270 8633
rect 3000 8473 3270 8607
rect 3000 8447 3119 8473
rect 3145 8447 3270 8473
rect 3000 8313 3270 8447
rect 3000 8287 3119 8313
rect 3145 8287 3270 8313
rect 3000 8153 3270 8287
rect 3000 8127 3119 8153
rect 3145 8127 3270 8153
rect 3000 7993 3270 8127
rect 3000 7967 3119 7993
rect 3145 7967 3270 7993
rect 3000 7833 3270 7967
rect 3000 7807 3119 7833
rect 3145 7807 3270 7833
rect 3000 7673 3270 7807
rect 3000 7647 3119 7673
rect 3145 7647 3270 7673
rect 3000 7513 3270 7647
rect 3000 7487 3119 7513
rect 3145 7487 3270 7513
rect 3000 7353 3270 7487
rect 3000 7327 3119 7353
rect 3145 7327 3270 7353
rect 3000 7193 3270 7327
rect 3000 7167 3119 7193
rect 3145 7167 3270 7193
rect 3000 7033 3270 7167
rect 3000 7007 3119 7033
rect 3145 7007 3270 7033
rect 3000 6873 3270 7007
rect 3000 6847 3119 6873
rect 3145 6847 3270 6873
rect 3000 6713 3270 6847
rect 3000 6687 3119 6713
rect 3145 6687 3270 6713
rect 3000 6553 3270 6687
rect 3000 6527 3119 6553
rect 3145 6527 3270 6553
rect 3000 6393 3270 6527
rect 3000 6367 3119 6393
rect 3145 6367 3270 6393
rect 3000 6233 3270 6367
rect 3000 6207 3119 6233
rect 3145 6207 3270 6233
rect 3000 6073 3270 6207
rect 3000 6047 3119 6073
rect 3145 6047 3270 6073
rect 3000 5913 3270 6047
rect 3000 5887 3119 5913
rect 3145 5887 3270 5913
rect 3000 5770 3270 5887
rect 6730 9113 7000 9230
rect 6730 9087 6852 9113
rect 6878 9087 7000 9113
rect 6730 8953 7000 9087
rect 6730 8927 6852 8953
rect 6878 8927 7000 8953
rect 6730 8793 7000 8927
rect 6730 8767 6852 8793
rect 6878 8767 7000 8793
rect 6730 8633 7000 8767
rect 6730 8607 6852 8633
rect 6878 8607 7000 8633
rect 6730 8473 7000 8607
rect 6730 8447 6852 8473
rect 6878 8447 7000 8473
rect 6730 8313 7000 8447
rect 6730 8287 6852 8313
rect 6878 8287 7000 8313
rect 6730 8153 7000 8287
rect 6730 8127 6852 8153
rect 6878 8127 7000 8153
rect 6730 7993 7000 8127
rect 6730 7967 6852 7993
rect 6878 7967 7000 7993
rect 6730 7833 7000 7967
rect 6730 7807 6852 7833
rect 6878 7807 7000 7833
rect 6730 7673 7000 7807
rect 6730 7647 6852 7673
rect 6878 7647 7000 7673
rect 6730 7513 7000 7647
rect 6730 7487 6852 7513
rect 6878 7487 7000 7513
rect 6730 7353 7000 7487
rect 6730 7327 6852 7353
rect 6878 7327 7000 7353
rect 6730 7193 7000 7327
rect 6730 7167 6852 7193
rect 6878 7167 7000 7193
rect 6730 7033 7000 7167
rect 6730 7007 6852 7033
rect 6878 7007 7000 7033
rect 6730 6873 7000 7007
rect 6730 6847 6852 6873
rect 6878 6847 7000 6873
rect 6730 6713 7000 6847
rect 6730 6687 6852 6713
rect 6878 6687 7000 6713
rect 6730 6553 7000 6687
rect 6730 6527 6852 6553
rect 6878 6527 7000 6553
rect 6730 6393 7000 6527
rect 6730 6367 6852 6393
rect 6878 6367 7000 6393
rect 6730 6233 7000 6367
rect 6730 6207 6852 6233
rect 6878 6207 7000 6233
rect 6730 6073 7000 6207
rect 6730 6047 6852 6073
rect 6878 6047 7000 6073
rect 6730 5913 7000 6047
rect 6730 5887 6852 5913
rect 6878 5887 7000 5913
rect 6730 5770 7000 5887
rect 3000 5753 7000 5770
rect 3000 5727 3119 5753
rect 3145 5727 6852 5753
rect 6878 5727 7000 5753
rect 3000 5650 7000 5727
rect 3000 5624 3307 5650
rect 3333 5624 3467 5650
rect 3493 5624 3627 5650
rect 3653 5624 3787 5650
rect 3813 5624 3947 5650
rect 3973 5624 4107 5650
rect 4133 5624 4267 5650
rect 4293 5624 4427 5650
rect 4453 5624 4587 5650
rect 4613 5624 4747 5650
rect 4773 5624 4907 5650
rect 4933 5624 5067 5650
rect 5093 5624 5227 5650
rect 5253 5624 5387 5650
rect 5413 5624 5547 5650
rect 5573 5624 5707 5650
rect 5733 5624 5867 5650
rect 5893 5624 6027 5650
rect 6053 5624 6187 5650
rect 6213 5624 6347 5650
rect 6373 5624 6507 5650
rect 6533 5624 6667 5650
rect 6693 5624 7000 5650
rect 3000 5500 7000 5624
rect 9000 9378 13000 9500
rect 9000 9352 9307 9378
rect 9333 9352 9467 9378
rect 9493 9352 9627 9378
rect 9653 9352 9787 9378
rect 9813 9352 9947 9378
rect 9973 9352 10107 9378
rect 10133 9352 10267 9378
rect 10293 9352 10427 9378
rect 10453 9352 10587 9378
rect 10613 9352 10747 9378
rect 10773 9352 10907 9378
rect 10933 9352 11067 9378
rect 11093 9352 11227 9378
rect 11253 9352 11387 9378
rect 11413 9352 11547 9378
rect 11573 9352 11707 9378
rect 11733 9352 11867 9378
rect 11893 9352 12027 9378
rect 12053 9352 12187 9378
rect 12213 9352 12347 9378
rect 12373 9352 12507 9378
rect 12533 9352 12667 9378
rect 12693 9352 13000 9378
rect 9000 9273 13000 9352
rect 9000 9247 9119 9273
rect 9145 9247 12852 9273
rect 12878 9247 13000 9273
rect 9000 9230 13000 9247
rect 9000 9113 9270 9230
rect 9000 9087 9119 9113
rect 9145 9087 9270 9113
rect 9000 8953 9270 9087
rect 9000 8927 9119 8953
rect 9145 8927 9270 8953
rect 9000 8793 9270 8927
rect 9000 8767 9119 8793
rect 9145 8767 9270 8793
rect 9000 8633 9270 8767
rect 9000 8607 9119 8633
rect 9145 8607 9270 8633
rect 9000 8473 9270 8607
rect 9000 8447 9119 8473
rect 9145 8447 9270 8473
rect 9000 8313 9270 8447
rect 9000 8287 9119 8313
rect 9145 8287 9270 8313
rect 9000 8153 9270 8287
rect 9000 8127 9119 8153
rect 9145 8127 9270 8153
rect 9000 7993 9270 8127
rect 9000 7967 9119 7993
rect 9145 7967 9270 7993
rect 9000 7833 9270 7967
rect 9000 7807 9119 7833
rect 9145 7807 9270 7833
rect 9000 7673 9270 7807
rect 9000 7647 9119 7673
rect 9145 7647 9270 7673
rect 9000 7513 9270 7647
rect 9000 7487 9119 7513
rect 9145 7487 9270 7513
rect 9000 7353 9270 7487
rect 9000 7327 9119 7353
rect 9145 7327 9270 7353
rect 9000 7193 9270 7327
rect 9000 7167 9119 7193
rect 9145 7167 9270 7193
rect 9000 7033 9270 7167
rect 9000 7007 9119 7033
rect 9145 7007 9270 7033
rect 9000 6873 9270 7007
rect 9000 6847 9119 6873
rect 9145 6847 9270 6873
rect 9000 6713 9270 6847
rect 9000 6687 9119 6713
rect 9145 6687 9270 6713
rect 9000 6553 9270 6687
rect 9000 6527 9119 6553
rect 9145 6527 9270 6553
rect 9000 6393 9270 6527
rect 9000 6367 9119 6393
rect 9145 6367 9270 6393
rect 9000 6233 9270 6367
rect 9000 6207 9119 6233
rect 9145 6207 9270 6233
rect 9000 6073 9270 6207
rect 9000 6047 9119 6073
rect 9145 6047 9270 6073
rect 9000 5913 9270 6047
rect 9000 5887 9119 5913
rect 9145 5887 9270 5913
rect 9000 5770 9270 5887
rect 12730 9113 13000 9230
rect 12730 9087 12852 9113
rect 12878 9087 13000 9113
rect 12730 8953 13000 9087
rect 12730 8927 12852 8953
rect 12878 8927 13000 8953
rect 12730 8793 13000 8927
rect 12730 8767 12852 8793
rect 12878 8767 13000 8793
rect 12730 8633 13000 8767
rect 12730 8607 12852 8633
rect 12878 8607 13000 8633
rect 12730 8473 13000 8607
rect 12730 8447 12852 8473
rect 12878 8447 13000 8473
rect 12730 8313 13000 8447
rect 12730 8287 12852 8313
rect 12878 8287 13000 8313
rect 12730 8153 13000 8287
rect 12730 8127 12852 8153
rect 12878 8127 13000 8153
rect 12730 7993 13000 8127
rect 12730 7967 12852 7993
rect 12878 7967 13000 7993
rect 12730 7833 13000 7967
rect 12730 7807 12852 7833
rect 12878 7807 13000 7833
rect 12730 7673 13000 7807
rect 12730 7647 12852 7673
rect 12878 7647 13000 7673
rect 12730 7513 13000 7647
rect 12730 7487 12852 7513
rect 12878 7487 13000 7513
rect 12730 7353 13000 7487
rect 12730 7327 12852 7353
rect 12878 7327 13000 7353
rect 12730 7193 13000 7327
rect 12730 7167 12852 7193
rect 12878 7167 13000 7193
rect 12730 7033 13000 7167
rect 12730 7007 12852 7033
rect 12878 7007 13000 7033
rect 12730 6873 13000 7007
rect 12730 6847 12852 6873
rect 12878 6847 13000 6873
rect 12730 6713 13000 6847
rect 12730 6687 12852 6713
rect 12878 6687 13000 6713
rect 12730 6553 13000 6687
rect 12730 6527 12852 6553
rect 12878 6527 13000 6553
rect 12730 6393 13000 6527
rect 12730 6367 12852 6393
rect 12878 6367 13000 6393
rect 12730 6233 13000 6367
rect 12730 6207 12852 6233
rect 12878 6207 13000 6233
rect 12730 6073 13000 6207
rect 12730 6047 12852 6073
rect 12878 6047 13000 6073
rect 12730 5913 13000 6047
rect 12730 5887 12852 5913
rect 12878 5887 13000 5913
rect 12730 5770 13000 5887
rect 9000 5753 13000 5770
rect 9000 5727 9119 5753
rect 9145 5727 12852 5753
rect 12878 5727 13000 5753
rect 9000 5650 13000 5727
rect 9000 5624 9307 5650
rect 9333 5624 9467 5650
rect 9493 5624 9627 5650
rect 9653 5624 9787 5650
rect 9813 5624 9947 5650
rect 9973 5624 10107 5650
rect 10133 5624 10267 5650
rect 10293 5624 10427 5650
rect 10453 5624 10587 5650
rect 10613 5624 10747 5650
rect 10773 5624 10907 5650
rect 10933 5624 11067 5650
rect 11093 5624 11227 5650
rect 11253 5624 11387 5650
rect 11413 5624 11547 5650
rect 11573 5624 11707 5650
rect 11733 5624 11867 5650
rect 11893 5624 12027 5650
rect 12053 5624 12187 5650
rect 12213 5624 12347 5650
rect 12373 5624 12507 5650
rect 12533 5624 12667 5650
rect 12693 5624 13000 5650
rect 9000 5500 13000 5624
rect 15000 9378 19000 9500
rect 15000 9352 15307 9378
rect 15333 9352 15467 9378
rect 15493 9352 15627 9378
rect 15653 9352 15787 9378
rect 15813 9352 15947 9378
rect 15973 9352 16107 9378
rect 16133 9352 16267 9378
rect 16293 9352 16427 9378
rect 16453 9352 16587 9378
rect 16613 9352 16747 9378
rect 16773 9352 16907 9378
rect 16933 9352 17067 9378
rect 17093 9352 17227 9378
rect 17253 9352 17387 9378
rect 17413 9352 17547 9378
rect 17573 9352 17707 9378
rect 17733 9352 17867 9378
rect 17893 9352 18027 9378
rect 18053 9352 18187 9378
rect 18213 9352 18347 9378
rect 18373 9352 18507 9378
rect 18533 9352 18667 9378
rect 18693 9352 19000 9378
rect 15000 9273 19000 9352
rect 15000 9247 15119 9273
rect 15145 9247 18852 9273
rect 18878 9247 19000 9273
rect 15000 9230 19000 9247
rect 15000 9113 15270 9230
rect 15000 9087 15119 9113
rect 15145 9087 15270 9113
rect 15000 8953 15270 9087
rect 15000 8927 15119 8953
rect 15145 8927 15270 8953
rect 15000 8793 15270 8927
rect 15000 8767 15119 8793
rect 15145 8767 15270 8793
rect 15000 8633 15270 8767
rect 15000 8607 15119 8633
rect 15145 8607 15270 8633
rect 15000 8473 15270 8607
rect 15000 8447 15119 8473
rect 15145 8447 15270 8473
rect 15000 8313 15270 8447
rect 15000 8287 15119 8313
rect 15145 8287 15270 8313
rect 15000 8153 15270 8287
rect 15000 8127 15119 8153
rect 15145 8127 15270 8153
rect 15000 7993 15270 8127
rect 15000 7967 15119 7993
rect 15145 7967 15270 7993
rect 15000 7833 15270 7967
rect 15000 7807 15119 7833
rect 15145 7807 15270 7833
rect 15000 7673 15270 7807
rect 15000 7647 15119 7673
rect 15145 7647 15270 7673
rect 15000 7513 15270 7647
rect 15000 7487 15119 7513
rect 15145 7487 15270 7513
rect 15000 7353 15270 7487
rect 15000 7327 15119 7353
rect 15145 7327 15270 7353
rect 15000 7193 15270 7327
rect 15000 7167 15119 7193
rect 15145 7167 15270 7193
rect 15000 7033 15270 7167
rect 15000 7007 15119 7033
rect 15145 7007 15270 7033
rect 15000 6873 15270 7007
rect 15000 6847 15119 6873
rect 15145 6847 15270 6873
rect 15000 6713 15270 6847
rect 15000 6687 15119 6713
rect 15145 6687 15270 6713
rect 15000 6553 15270 6687
rect 15000 6527 15119 6553
rect 15145 6527 15270 6553
rect 15000 6393 15270 6527
rect 15000 6367 15119 6393
rect 15145 6367 15270 6393
rect 15000 6233 15270 6367
rect 15000 6207 15119 6233
rect 15145 6207 15270 6233
rect 15000 6073 15270 6207
rect 15000 6047 15119 6073
rect 15145 6047 15270 6073
rect 15000 5913 15270 6047
rect 15000 5887 15119 5913
rect 15145 5887 15270 5913
rect 15000 5770 15270 5887
rect 18730 9113 19000 9230
rect 18730 9087 18852 9113
rect 18878 9087 19000 9113
rect 18730 8953 19000 9087
rect 18730 8927 18852 8953
rect 18878 8927 19000 8953
rect 18730 8793 19000 8927
rect 18730 8767 18852 8793
rect 18878 8767 19000 8793
rect 18730 8633 19000 8767
rect 18730 8607 18852 8633
rect 18878 8607 19000 8633
rect 18730 8473 19000 8607
rect 18730 8447 18852 8473
rect 18878 8447 19000 8473
rect 18730 8313 19000 8447
rect 18730 8287 18852 8313
rect 18878 8287 19000 8313
rect 18730 8153 19000 8287
rect 18730 8127 18852 8153
rect 18878 8127 19000 8153
rect 18730 7993 19000 8127
rect 18730 7967 18852 7993
rect 18878 7967 19000 7993
rect 18730 7833 19000 7967
rect 18730 7807 18852 7833
rect 18878 7807 19000 7833
rect 18730 7673 19000 7807
rect 18730 7647 18852 7673
rect 18878 7647 19000 7673
rect 18730 7513 19000 7647
rect 18730 7487 18852 7513
rect 18878 7487 19000 7513
rect 18730 7353 19000 7487
rect 18730 7327 18852 7353
rect 18878 7327 19000 7353
rect 18730 7193 19000 7327
rect 18730 7167 18852 7193
rect 18878 7167 19000 7193
rect 18730 7033 19000 7167
rect 18730 7007 18852 7033
rect 18878 7007 19000 7033
rect 18730 6873 19000 7007
rect 18730 6847 18852 6873
rect 18878 6847 19000 6873
rect 18730 6713 19000 6847
rect 18730 6687 18852 6713
rect 18878 6687 19000 6713
rect 18730 6553 19000 6687
rect 18730 6527 18852 6553
rect 18878 6527 19000 6553
rect 18730 6393 19000 6527
rect 18730 6367 18852 6393
rect 18878 6367 19000 6393
rect 18730 6233 19000 6367
rect 18730 6207 18852 6233
rect 18878 6207 19000 6233
rect 18730 6073 19000 6207
rect 18730 6047 18852 6073
rect 18878 6047 19000 6073
rect 18730 5913 19000 6047
rect 18730 5887 18852 5913
rect 18878 5887 19000 5913
rect 18730 5770 19000 5887
rect 15000 5753 19000 5770
rect 15000 5727 15119 5753
rect 15145 5727 18852 5753
rect 18878 5727 19000 5753
rect 15000 5650 19000 5727
rect 15000 5624 15307 5650
rect 15333 5624 15467 5650
rect 15493 5624 15627 5650
rect 15653 5624 15787 5650
rect 15813 5624 15947 5650
rect 15973 5624 16107 5650
rect 16133 5624 16267 5650
rect 16293 5624 16427 5650
rect 16453 5624 16587 5650
rect 16613 5624 16747 5650
rect 16773 5624 16907 5650
rect 16933 5624 17067 5650
rect 17093 5624 17227 5650
rect 17253 5624 17387 5650
rect 17413 5624 17547 5650
rect 17573 5624 17707 5650
rect 17733 5624 17867 5650
rect 17893 5624 18027 5650
rect 18053 5624 18187 5650
rect 18213 5624 18347 5650
rect 18373 5624 18507 5650
rect 18533 5624 18667 5650
rect 18693 5624 19000 5650
rect 15000 5500 19000 5624
rect 21000 9378 25000 9500
rect 21000 9352 21307 9378
rect 21333 9352 21467 9378
rect 21493 9352 21627 9378
rect 21653 9352 21787 9378
rect 21813 9352 21947 9378
rect 21973 9352 22107 9378
rect 22133 9352 22267 9378
rect 22293 9352 22427 9378
rect 22453 9352 22587 9378
rect 22613 9352 22747 9378
rect 22773 9352 22907 9378
rect 22933 9352 23067 9378
rect 23093 9352 23227 9378
rect 23253 9352 23387 9378
rect 23413 9352 23547 9378
rect 23573 9352 23707 9378
rect 23733 9352 23867 9378
rect 23893 9352 24027 9378
rect 24053 9352 24187 9378
rect 24213 9352 24347 9378
rect 24373 9352 24507 9378
rect 24533 9352 24667 9378
rect 24693 9352 25000 9378
rect 21000 9273 25000 9352
rect 21000 9247 21119 9273
rect 21145 9247 24852 9273
rect 24878 9247 25000 9273
rect 21000 9230 25000 9247
rect 21000 9113 21270 9230
rect 21000 9087 21119 9113
rect 21145 9087 21270 9113
rect 21000 8953 21270 9087
rect 21000 8927 21119 8953
rect 21145 8927 21270 8953
rect 21000 8793 21270 8927
rect 21000 8767 21119 8793
rect 21145 8767 21270 8793
rect 21000 8633 21270 8767
rect 21000 8607 21119 8633
rect 21145 8607 21270 8633
rect 21000 8473 21270 8607
rect 21000 8447 21119 8473
rect 21145 8447 21270 8473
rect 21000 8313 21270 8447
rect 21000 8287 21119 8313
rect 21145 8287 21270 8313
rect 21000 8153 21270 8287
rect 21000 8127 21119 8153
rect 21145 8127 21270 8153
rect 21000 7993 21270 8127
rect 21000 7967 21119 7993
rect 21145 7967 21270 7993
rect 21000 7833 21270 7967
rect 21000 7807 21119 7833
rect 21145 7807 21270 7833
rect 21000 7673 21270 7807
rect 21000 7647 21119 7673
rect 21145 7647 21270 7673
rect 21000 7513 21270 7647
rect 21000 7487 21119 7513
rect 21145 7487 21270 7513
rect 21000 7353 21270 7487
rect 21000 7327 21119 7353
rect 21145 7327 21270 7353
rect 21000 7193 21270 7327
rect 21000 7167 21119 7193
rect 21145 7167 21270 7193
rect 21000 7033 21270 7167
rect 21000 7007 21119 7033
rect 21145 7007 21270 7033
rect 21000 6873 21270 7007
rect 21000 6847 21119 6873
rect 21145 6847 21270 6873
rect 21000 6713 21270 6847
rect 21000 6687 21119 6713
rect 21145 6687 21270 6713
rect 21000 6553 21270 6687
rect 21000 6527 21119 6553
rect 21145 6527 21270 6553
rect 21000 6393 21270 6527
rect 21000 6367 21119 6393
rect 21145 6367 21270 6393
rect 21000 6233 21270 6367
rect 21000 6207 21119 6233
rect 21145 6207 21270 6233
rect 21000 6073 21270 6207
rect 21000 6047 21119 6073
rect 21145 6047 21270 6073
rect 21000 5913 21270 6047
rect 21000 5887 21119 5913
rect 21145 5887 21270 5913
rect 21000 5770 21270 5887
rect 24730 9113 25000 9230
rect 24730 9087 24852 9113
rect 24878 9087 25000 9113
rect 24730 8953 25000 9087
rect 24730 8927 24852 8953
rect 24878 8927 25000 8953
rect 24730 8793 25000 8927
rect 24730 8767 24852 8793
rect 24878 8767 25000 8793
rect 24730 8633 25000 8767
rect 24730 8607 24852 8633
rect 24878 8607 25000 8633
rect 24730 8473 25000 8607
rect 24730 8447 24852 8473
rect 24878 8447 25000 8473
rect 24730 8313 25000 8447
rect 24730 8287 24852 8313
rect 24878 8287 25000 8313
rect 24730 8153 25000 8287
rect 24730 8127 24852 8153
rect 24878 8127 25000 8153
rect 24730 7993 25000 8127
rect 24730 7967 24852 7993
rect 24878 7967 25000 7993
rect 24730 7833 25000 7967
rect 24730 7807 24852 7833
rect 24878 7807 25000 7833
rect 24730 7673 25000 7807
rect 24730 7647 24852 7673
rect 24878 7647 25000 7673
rect 24730 7513 25000 7647
rect 24730 7487 24852 7513
rect 24878 7487 25000 7513
rect 24730 7353 25000 7487
rect 24730 7327 24852 7353
rect 24878 7327 25000 7353
rect 24730 7193 25000 7327
rect 24730 7167 24852 7193
rect 24878 7167 25000 7193
rect 24730 7033 25000 7167
rect 24730 7007 24852 7033
rect 24878 7007 25000 7033
rect 24730 6873 25000 7007
rect 24730 6847 24852 6873
rect 24878 6847 25000 6873
rect 24730 6713 25000 6847
rect 24730 6687 24852 6713
rect 24878 6687 25000 6713
rect 24730 6553 25000 6687
rect 24730 6527 24852 6553
rect 24878 6527 25000 6553
rect 24730 6393 25000 6527
rect 24730 6367 24852 6393
rect 24878 6367 25000 6393
rect 24730 6233 25000 6367
rect 24730 6207 24852 6233
rect 24878 6207 25000 6233
rect 24730 6073 25000 6207
rect 24730 6047 24852 6073
rect 24878 6047 25000 6073
rect 24730 5913 25000 6047
rect 24730 5887 24852 5913
rect 24878 5887 25000 5913
rect 24730 5770 25000 5887
rect 21000 5753 25000 5770
rect 21000 5727 21119 5753
rect 21145 5727 24852 5753
rect 24878 5727 25000 5753
rect 21000 5650 25000 5727
rect 21000 5624 21307 5650
rect 21333 5624 21467 5650
rect 21493 5624 21627 5650
rect 21653 5624 21787 5650
rect 21813 5624 21947 5650
rect 21973 5624 22107 5650
rect 22133 5624 22267 5650
rect 22293 5624 22427 5650
rect 22453 5624 22587 5650
rect 22613 5624 22747 5650
rect 22773 5624 22907 5650
rect 22933 5624 23067 5650
rect 23093 5624 23227 5650
rect 23253 5624 23387 5650
rect 23413 5624 23547 5650
rect 23573 5624 23707 5650
rect 23733 5624 23867 5650
rect 23893 5624 24027 5650
rect 24053 5624 24187 5650
rect 24213 5624 24347 5650
rect 24373 5624 24507 5650
rect 24533 5624 24667 5650
rect 24693 5624 25000 5650
rect 21000 5500 25000 5624
rect 3000 3378 7000 3500
rect 3000 3352 3307 3378
rect 3333 3352 3467 3378
rect 3493 3352 3627 3378
rect 3653 3352 3787 3378
rect 3813 3352 3947 3378
rect 3973 3352 4107 3378
rect 4133 3352 4267 3378
rect 4293 3352 4427 3378
rect 4453 3352 4587 3378
rect 4613 3352 4747 3378
rect 4773 3352 4907 3378
rect 4933 3352 5067 3378
rect 5093 3352 5227 3378
rect 5253 3352 5387 3378
rect 5413 3352 5547 3378
rect 5573 3352 5707 3378
rect 5733 3352 5867 3378
rect 5893 3352 6027 3378
rect 6053 3352 6187 3378
rect 6213 3352 6347 3378
rect 6373 3352 6507 3378
rect 6533 3352 6667 3378
rect 6693 3352 7000 3378
rect 3000 3273 7000 3352
rect 3000 3247 3119 3273
rect 3145 3247 6852 3273
rect 6878 3247 7000 3273
rect 3000 3230 7000 3247
rect 3000 3113 3270 3230
rect 3000 3087 3119 3113
rect 3145 3087 3270 3113
rect 3000 2953 3270 3087
rect 3000 2927 3119 2953
rect 3145 2927 3270 2953
rect 3000 2793 3270 2927
rect 3000 2767 3119 2793
rect 3145 2767 3270 2793
rect 3000 2633 3270 2767
rect 3000 2607 3119 2633
rect 3145 2607 3270 2633
rect 3000 2473 3270 2607
rect 3000 2447 3119 2473
rect 3145 2447 3270 2473
rect 3000 2313 3270 2447
rect 3000 2287 3119 2313
rect 3145 2287 3270 2313
rect 3000 2153 3270 2287
rect 3000 2127 3119 2153
rect 3145 2127 3270 2153
rect 3000 1993 3270 2127
rect 3000 1967 3119 1993
rect 3145 1967 3270 1993
rect 3000 1833 3270 1967
rect 3000 1807 3119 1833
rect 3145 1807 3270 1833
rect 3000 1673 3270 1807
rect 3000 1647 3119 1673
rect 3145 1647 3270 1673
rect 3000 1513 3270 1647
rect 3000 1487 3119 1513
rect 3145 1487 3270 1513
rect 3000 1353 3270 1487
rect 3000 1327 3119 1353
rect 3145 1327 3270 1353
rect 3000 1193 3270 1327
rect 3000 1167 3119 1193
rect 3145 1167 3270 1193
rect 3000 1033 3270 1167
rect 3000 1007 3119 1033
rect 3145 1007 3270 1033
rect 3000 873 3270 1007
rect 3000 847 3119 873
rect 3145 847 3270 873
rect 3000 713 3270 847
rect 3000 687 3119 713
rect 3145 687 3270 713
rect 3000 553 3270 687
rect 3000 527 3119 553
rect 3145 527 3270 553
rect 3000 393 3270 527
rect 3000 367 3119 393
rect 3145 367 3270 393
rect 3000 233 3270 367
rect 3000 207 3119 233
rect 3145 207 3270 233
rect 3000 73 3270 207
rect 3000 47 3119 73
rect 3145 47 3270 73
rect 3000 -87 3270 47
rect 3000 -113 3119 -87
rect 3145 -113 3270 -87
rect 3000 -230 3270 -113
rect 6730 3113 7000 3230
rect 6730 3087 6852 3113
rect 6878 3087 7000 3113
rect 6730 2953 7000 3087
rect 6730 2927 6852 2953
rect 6878 2927 7000 2953
rect 6730 2793 7000 2927
rect 6730 2767 6852 2793
rect 6878 2767 7000 2793
rect 6730 2633 7000 2767
rect 6730 2607 6852 2633
rect 6878 2607 7000 2633
rect 6730 2473 7000 2607
rect 6730 2447 6852 2473
rect 6878 2447 7000 2473
rect 6730 2313 7000 2447
rect 6730 2287 6852 2313
rect 6878 2287 7000 2313
rect 6730 2153 7000 2287
rect 6730 2127 6852 2153
rect 6878 2127 7000 2153
rect 6730 1993 7000 2127
rect 6730 1967 6852 1993
rect 6878 1967 7000 1993
rect 6730 1833 7000 1967
rect 6730 1807 6852 1833
rect 6878 1807 7000 1833
rect 6730 1673 7000 1807
rect 6730 1647 6852 1673
rect 6878 1647 7000 1673
rect 6730 1513 7000 1647
rect 6730 1487 6852 1513
rect 6878 1487 7000 1513
rect 6730 1353 7000 1487
rect 6730 1327 6852 1353
rect 6878 1327 7000 1353
rect 6730 1193 7000 1327
rect 6730 1167 6852 1193
rect 6878 1167 7000 1193
rect 6730 1033 7000 1167
rect 6730 1007 6852 1033
rect 6878 1007 7000 1033
rect 6730 873 7000 1007
rect 6730 847 6852 873
rect 6878 847 7000 873
rect 6730 713 7000 847
rect 6730 687 6852 713
rect 6878 687 7000 713
rect 6730 553 7000 687
rect 6730 527 6852 553
rect 6878 527 7000 553
rect 6730 393 7000 527
rect 6730 367 6852 393
rect 6878 367 7000 393
rect 6730 233 7000 367
rect 6730 207 6852 233
rect 6878 207 7000 233
rect 6730 73 7000 207
rect 6730 47 6852 73
rect 6878 47 7000 73
rect 6730 -87 7000 47
rect 6730 -113 6852 -87
rect 6878 -113 7000 -87
rect 6730 -230 7000 -113
rect 3000 -247 7000 -230
rect 3000 -273 3119 -247
rect 3145 -273 6852 -247
rect 6878 -273 7000 -247
rect 3000 -350 7000 -273
rect 3000 -376 3307 -350
rect 3333 -376 3467 -350
rect 3493 -376 3627 -350
rect 3653 -376 3787 -350
rect 3813 -376 3947 -350
rect 3973 -376 4107 -350
rect 4133 -376 4267 -350
rect 4293 -376 4427 -350
rect 4453 -376 4587 -350
rect 4613 -376 4747 -350
rect 4773 -376 4907 -350
rect 4933 -376 5067 -350
rect 5093 -376 5227 -350
rect 5253 -376 5387 -350
rect 5413 -376 5547 -350
rect 5573 -376 5707 -350
rect 5733 -376 5867 -350
rect 5893 -376 6027 -350
rect 6053 -376 6187 -350
rect 6213 -376 6347 -350
rect 6373 -376 6507 -350
rect 6533 -376 6667 -350
rect 6693 -376 7000 -350
rect 3000 -500 7000 -376
rect 9000 3378 13000 3500
rect 9000 3352 9307 3378
rect 9333 3352 9467 3378
rect 9493 3352 9627 3378
rect 9653 3352 9787 3378
rect 9813 3352 9947 3378
rect 9973 3352 10107 3378
rect 10133 3352 10267 3378
rect 10293 3352 10427 3378
rect 10453 3352 10587 3378
rect 10613 3352 10747 3378
rect 10773 3352 10907 3378
rect 10933 3352 11067 3378
rect 11093 3352 11227 3378
rect 11253 3352 11387 3378
rect 11413 3352 11547 3378
rect 11573 3352 11707 3378
rect 11733 3352 11867 3378
rect 11893 3352 12027 3378
rect 12053 3352 12187 3378
rect 12213 3352 12347 3378
rect 12373 3352 12507 3378
rect 12533 3352 12667 3378
rect 12693 3352 13000 3378
rect 9000 3273 13000 3352
rect 9000 3247 9119 3273
rect 9145 3247 12852 3273
rect 12878 3247 13000 3273
rect 9000 3230 13000 3247
rect 9000 3113 9270 3230
rect 9000 3087 9119 3113
rect 9145 3087 9270 3113
rect 9000 2953 9270 3087
rect 9000 2927 9119 2953
rect 9145 2927 9270 2953
rect 9000 2793 9270 2927
rect 9000 2767 9119 2793
rect 9145 2767 9270 2793
rect 9000 2633 9270 2767
rect 9000 2607 9119 2633
rect 9145 2607 9270 2633
rect 9000 2473 9270 2607
rect 9000 2447 9119 2473
rect 9145 2447 9270 2473
rect 9000 2313 9270 2447
rect 9000 2287 9119 2313
rect 9145 2287 9270 2313
rect 9000 2153 9270 2287
rect 9000 2127 9119 2153
rect 9145 2127 9270 2153
rect 9000 1993 9270 2127
rect 9000 1967 9119 1993
rect 9145 1967 9270 1993
rect 9000 1833 9270 1967
rect 9000 1807 9119 1833
rect 9145 1807 9270 1833
rect 9000 1673 9270 1807
rect 9000 1647 9119 1673
rect 9145 1647 9270 1673
rect 9000 1513 9270 1647
rect 9000 1487 9119 1513
rect 9145 1487 9270 1513
rect 9000 1353 9270 1487
rect 9000 1327 9119 1353
rect 9145 1327 9270 1353
rect 9000 1193 9270 1327
rect 9000 1167 9119 1193
rect 9145 1167 9270 1193
rect 9000 1033 9270 1167
rect 9000 1007 9119 1033
rect 9145 1007 9270 1033
rect 9000 873 9270 1007
rect 9000 847 9119 873
rect 9145 847 9270 873
rect 9000 713 9270 847
rect 9000 687 9119 713
rect 9145 687 9270 713
rect 9000 553 9270 687
rect 9000 527 9119 553
rect 9145 527 9270 553
rect 9000 393 9270 527
rect 9000 367 9119 393
rect 9145 367 9270 393
rect 9000 233 9270 367
rect 9000 207 9119 233
rect 9145 207 9270 233
rect 9000 73 9270 207
rect 9000 47 9119 73
rect 9145 47 9270 73
rect 9000 -87 9270 47
rect 9000 -113 9119 -87
rect 9145 -113 9270 -87
rect 9000 -230 9270 -113
rect 12730 3113 13000 3230
rect 12730 3087 12852 3113
rect 12878 3087 13000 3113
rect 12730 2953 13000 3087
rect 12730 2927 12852 2953
rect 12878 2927 13000 2953
rect 12730 2793 13000 2927
rect 12730 2767 12852 2793
rect 12878 2767 13000 2793
rect 12730 2633 13000 2767
rect 12730 2607 12852 2633
rect 12878 2607 13000 2633
rect 12730 2473 13000 2607
rect 12730 2447 12852 2473
rect 12878 2447 13000 2473
rect 12730 2313 13000 2447
rect 12730 2287 12852 2313
rect 12878 2287 13000 2313
rect 12730 2153 13000 2287
rect 12730 2127 12852 2153
rect 12878 2127 13000 2153
rect 12730 1993 13000 2127
rect 12730 1967 12852 1993
rect 12878 1967 13000 1993
rect 12730 1833 13000 1967
rect 12730 1807 12852 1833
rect 12878 1807 13000 1833
rect 12730 1673 13000 1807
rect 12730 1647 12852 1673
rect 12878 1647 13000 1673
rect 12730 1513 13000 1647
rect 12730 1487 12852 1513
rect 12878 1487 13000 1513
rect 12730 1353 13000 1487
rect 12730 1327 12852 1353
rect 12878 1327 13000 1353
rect 12730 1193 13000 1327
rect 12730 1167 12852 1193
rect 12878 1167 13000 1193
rect 12730 1033 13000 1167
rect 12730 1007 12852 1033
rect 12878 1007 13000 1033
rect 12730 873 13000 1007
rect 12730 847 12852 873
rect 12878 847 13000 873
rect 12730 713 13000 847
rect 12730 687 12852 713
rect 12878 687 13000 713
rect 12730 553 13000 687
rect 12730 527 12852 553
rect 12878 527 13000 553
rect 12730 393 13000 527
rect 12730 367 12852 393
rect 12878 367 13000 393
rect 12730 233 13000 367
rect 12730 207 12852 233
rect 12878 207 13000 233
rect 12730 73 13000 207
rect 12730 47 12852 73
rect 12878 47 13000 73
rect 12730 -87 13000 47
rect 12730 -113 12852 -87
rect 12878 -113 13000 -87
rect 12730 -230 13000 -113
rect 9000 -247 13000 -230
rect 9000 -273 9119 -247
rect 9145 -273 12852 -247
rect 12878 -273 13000 -247
rect 9000 -350 13000 -273
rect 9000 -376 9307 -350
rect 9333 -376 9467 -350
rect 9493 -376 9627 -350
rect 9653 -376 9787 -350
rect 9813 -376 9947 -350
rect 9973 -376 10107 -350
rect 10133 -376 10267 -350
rect 10293 -376 10427 -350
rect 10453 -376 10587 -350
rect 10613 -376 10747 -350
rect 10773 -376 10907 -350
rect 10933 -376 11067 -350
rect 11093 -376 11227 -350
rect 11253 -376 11387 -350
rect 11413 -376 11547 -350
rect 11573 -376 11707 -350
rect 11733 -376 11867 -350
rect 11893 -376 12027 -350
rect 12053 -376 12187 -350
rect 12213 -376 12347 -350
rect 12373 -376 12507 -350
rect 12533 -376 12667 -350
rect 12693 -376 13000 -350
rect 9000 -500 13000 -376
rect 15000 3378 19000 3500
rect 15000 3352 15307 3378
rect 15333 3352 15467 3378
rect 15493 3352 15627 3378
rect 15653 3352 15787 3378
rect 15813 3352 15947 3378
rect 15973 3352 16107 3378
rect 16133 3352 16267 3378
rect 16293 3352 16427 3378
rect 16453 3352 16587 3378
rect 16613 3352 16747 3378
rect 16773 3352 16907 3378
rect 16933 3352 17067 3378
rect 17093 3352 17227 3378
rect 17253 3352 17387 3378
rect 17413 3352 17547 3378
rect 17573 3352 17707 3378
rect 17733 3352 17867 3378
rect 17893 3352 18027 3378
rect 18053 3352 18187 3378
rect 18213 3352 18347 3378
rect 18373 3352 18507 3378
rect 18533 3352 18667 3378
rect 18693 3352 19000 3378
rect 15000 3273 19000 3352
rect 15000 3247 15119 3273
rect 15145 3247 18852 3273
rect 18878 3247 19000 3273
rect 15000 3230 19000 3247
rect 15000 3113 15270 3230
rect 15000 3087 15119 3113
rect 15145 3087 15270 3113
rect 15000 2953 15270 3087
rect 15000 2927 15119 2953
rect 15145 2927 15270 2953
rect 15000 2793 15270 2927
rect 15000 2767 15119 2793
rect 15145 2767 15270 2793
rect 15000 2633 15270 2767
rect 15000 2607 15119 2633
rect 15145 2607 15270 2633
rect 15000 2473 15270 2607
rect 15000 2447 15119 2473
rect 15145 2447 15270 2473
rect 15000 2313 15270 2447
rect 15000 2287 15119 2313
rect 15145 2287 15270 2313
rect 15000 2153 15270 2287
rect 15000 2127 15119 2153
rect 15145 2127 15270 2153
rect 15000 1993 15270 2127
rect 15000 1967 15119 1993
rect 15145 1967 15270 1993
rect 15000 1833 15270 1967
rect 15000 1807 15119 1833
rect 15145 1807 15270 1833
rect 15000 1673 15270 1807
rect 15000 1647 15119 1673
rect 15145 1647 15270 1673
rect 15000 1513 15270 1647
rect 15000 1487 15119 1513
rect 15145 1487 15270 1513
rect 15000 1353 15270 1487
rect 15000 1327 15119 1353
rect 15145 1327 15270 1353
rect 15000 1193 15270 1327
rect 15000 1167 15119 1193
rect 15145 1167 15270 1193
rect 15000 1033 15270 1167
rect 15000 1007 15119 1033
rect 15145 1007 15270 1033
rect 15000 873 15270 1007
rect 15000 847 15119 873
rect 15145 847 15270 873
rect 15000 713 15270 847
rect 15000 687 15119 713
rect 15145 687 15270 713
rect 15000 553 15270 687
rect 15000 527 15119 553
rect 15145 527 15270 553
rect 15000 393 15270 527
rect 15000 367 15119 393
rect 15145 367 15270 393
rect 15000 233 15270 367
rect 15000 207 15119 233
rect 15145 207 15270 233
rect 15000 73 15270 207
rect 15000 47 15119 73
rect 15145 47 15270 73
rect 15000 -87 15270 47
rect 15000 -113 15119 -87
rect 15145 -113 15270 -87
rect 15000 -230 15270 -113
rect 18730 3113 19000 3230
rect 18730 3087 18852 3113
rect 18878 3087 19000 3113
rect 18730 2953 19000 3087
rect 18730 2927 18852 2953
rect 18878 2927 19000 2953
rect 18730 2793 19000 2927
rect 18730 2767 18852 2793
rect 18878 2767 19000 2793
rect 18730 2633 19000 2767
rect 18730 2607 18852 2633
rect 18878 2607 19000 2633
rect 18730 2473 19000 2607
rect 18730 2447 18852 2473
rect 18878 2447 19000 2473
rect 18730 2313 19000 2447
rect 18730 2287 18852 2313
rect 18878 2287 19000 2313
rect 18730 2153 19000 2287
rect 18730 2127 18852 2153
rect 18878 2127 19000 2153
rect 18730 1993 19000 2127
rect 18730 1967 18852 1993
rect 18878 1967 19000 1993
rect 18730 1833 19000 1967
rect 18730 1807 18852 1833
rect 18878 1807 19000 1833
rect 18730 1673 19000 1807
rect 18730 1647 18852 1673
rect 18878 1647 19000 1673
rect 18730 1513 19000 1647
rect 18730 1487 18852 1513
rect 18878 1487 19000 1513
rect 18730 1353 19000 1487
rect 18730 1327 18852 1353
rect 18878 1327 19000 1353
rect 18730 1193 19000 1327
rect 18730 1167 18852 1193
rect 18878 1167 19000 1193
rect 18730 1033 19000 1167
rect 18730 1007 18852 1033
rect 18878 1007 19000 1033
rect 18730 873 19000 1007
rect 18730 847 18852 873
rect 18878 847 19000 873
rect 18730 713 19000 847
rect 18730 687 18852 713
rect 18878 687 19000 713
rect 18730 553 19000 687
rect 18730 527 18852 553
rect 18878 527 19000 553
rect 18730 393 19000 527
rect 18730 367 18852 393
rect 18878 367 19000 393
rect 18730 233 19000 367
rect 18730 207 18852 233
rect 18878 207 19000 233
rect 18730 73 19000 207
rect 18730 47 18852 73
rect 18878 47 19000 73
rect 18730 -87 19000 47
rect 18730 -113 18852 -87
rect 18878 -113 19000 -87
rect 18730 -230 19000 -113
rect 15000 -247 19000 -230
rect 15000 -273 15119 -247
rect 15145 -273 18852 -247
rect 18878 -273 19000 -247
rect 15000 -350 19000 -273
rect 15000 -376 15307 -350
rect 15333 -376 15467 -350
rect 15493 -376 15627 -350
rect 15653 -376 15787 -350
rect 15813 -376 15947 -350
rect 15973 -376 16107 -350
rect 16133 -376 16267 -350
rect 16293 -376 16427 -350
rect 16453 -376 16587 -350
rect 16613 -376 16747 -350
rect 16773 -376 16907 -350
rect 16933 -376 17067 -350
rect 17093 -376 17227 -350
rect 17253 -376 17387 -350
rect 17413 -376 17547 -350
rect 17573 -376 17707 -350
rect 17733 -376 17867 -350
rect 17893 -376 18027 -350
rect 18053 -376 18187 -350
rect 18213 -376 18347 -350
rect 18373 -376 18507 -350
rect 18533 -376 18667 -350
rect 18693 -376 19000 -350
rect 15000 -500 19000 -376
rect 21000 3378 25000 3500
rect 21000 3352 21307 3378
rect 21333 3352 21467 3378
rect 21493 3352 21627 3378
rect 21653 3352 21787 3378
rect 21813 3352 21947 3378
rect 21973 3352 22107 3378
rect 22133 3352 22267 3378
rect 22293 3352 22427 3378
rect 22453 3352 22587 3378
rect 22613 3352 22747 3378
rect 22773 3352 22907 3378
rect 22933 3352 23067 3378
rect 23093 3352 23227 3378
rect 23253 3352 23387 3378
rect 23413 3352 23547 3378
rect 23573 3352 23707 3378
rect 23733 3352 23867 3378
rect 23893 3352 24027 3378
rect 24053 3352 24187 3378
rect 24213 3352 24347 3378
rect 24373 3352 24507 3378
rect 24533 3352 24667 3378
rect 24693 3352 25000 3378
rect 21000 3273 25000 3352
rect 21000 3247 21119 3273
rect 21145 3247 24852 3273
rect 24878 3247 25000 3273
rect 21000 3230 25000 3247
rect 21000 3113 21270 3230
rect 21000 3087 21119 3113
rect 21145 3087 21270 3113
rect 21000 2953 21270 3087
rect 21000 2927 21119 2953
rect 21145 2927 21270 2953
rect 21000 2793 21270 2927
rect 21000 2767 21119 2793
rect 21145 2767 21270 2793
rect 21000 2633 21270 2767
rect 21000 2607 21119 2633
rect 21145 2607 21270 2633
rect 21000 2473 21270 2607
rect 21000 2447 21119 2473
rect 21145 2447 21270 2473
rect 21000 2313 21270 2447
rect 21000 2287 21119 2313
rect 21145 2287 21270 2313
rect 21000 2153 21270 2287
rect 21000 2127 21119 2153
rect 21145 2127 21270 2153
rect 21000 1993 21270 2127
rect 21000 1967 21119 1993
rect 21145 1967 21270 1993
rect 21000 1833 21270 1967
rect 21000 1807 21119 1833
rect 21145 1807 21270 1833
rect 21000 1673 21270 1807
rect 21000 1647 21119 1673
rect 21145 1647 21270 1673
rect 21000 1513 21270 1647
rect 21000 1487 21119 1513
rect 21145 1487 21270 1513
rect 21000 1353 21270 1487
rect 21000 1327 21119 1353
rect 21145 1327 21270 1353
rect 21000 1193 21270 1327
rect 21000 1167 21119 1193
rect 21145 1167 21270 1193
rect 21000 1033 21270 1167
rect 21000 1007 21119 1033
rect 21145 1007 21270 1033
rect 21000 873 21270 1007
rect 21000 847 21119 873
rect 21145 847 21270 873
rect 21000 713 21270 847
rect 21000 687 21119 713
rect 21145 687 21270 713
rect 21000 553 21270 687
rect 21000 527 21119 553
rect 21145 527 21270 553
rect 21000 393 21270 527
rect 21000 367 21119 393
rect 21145 367 21270 393
rect 21000 233 21270 367
rect 21000 207 21119 233
rect 21145 207 21270 233
rect 21000 73 21270 207
rect 21000 47 21119 73
rect 21145 47 21270 73
rect 21000 -87 21270 47
rect 21000 -113 21119 -87
rect 21145 -113 21270 -87
rect 21000 -230 21270 -113
rect 24730 3113 25000 3230
rect 24730 3087 24852 3113
rect 24878 3087 25000 3113
rect 24730 2953 25000 3087
rect 24730 2927 24852 2953
rect 24878 2927 25000 2953
rect 24730 2793 25000 2927
rect 24730 2767 24852 2793
rect 24878 2767 25000 2793
rect 24730 2633 25000 2767
rect 24730 2607 24852 2633
rect 24878 2607 25000 2633
rect 24730 2473 25000 2607
rect 24730 2447 24852 2473
rect 24878 2447 25000 2473
rect 24730 2313 25000 2447
rect 24730 2287 24852 2313
rect 24878 2287 25000 2313
rect 24730 2153 25000 2287
rect 24730 2127 24852 2153
rect 24878 2127 25000 2153
rect 24730 1993 25000 2127
rect 24730 1967 24852 1993
rect 24878 1967 25000 1993
rect 24730 1833 25000 1967
rect 24730 1807 24852 1833
rect 24878 1807 25000 1833
rect 24730 1673 25000 1807
rect 24730 1647 24852 1673
rect 24878 1647 25000 1673
rect 24730 1513 25000 1647
rect 24730 1487 24852 1513
rect 24878 1487 25000 1513
rect 24730 1353 25000 1487
rect 24730 1327 24852 1353
rect 24878 1327 25000 1353
rect 24730 1193 25000 1327
rect 24730 1167 24852 1193
rect 24878 1167 25000 1193
rect 24730 1033 25000 1167
rect 24730 1007 24852 1033
rect 24878 1007 25000 1033
rect 24730 873 25000 1007
rect 24730 847 24852 873
rect 24878 847 25000 873
rect 24730 713 25000 847
rect 24730 687 24852 713
rect 24878 687 25000 713
rect 24730 553 25000 687
rect 24730 527 24852 553
rect 24878 527 25000 553
rect 24730 393 25000 527
rect 24730 367 24852 393
rect 24878 367 25000 393
rect 24730 233 25000 367
rect 24730 207 24852 233
rect 24878 207 25000 233
rect 24730 73 25000 207
rect 24730 47 24852 73
rect 24878 47 25000 73
rect 24730 -87 25000 47
rect 24730 -113 24852 -87
rect 24878 -113 25000 -87
rect 24730 -230 25000 -113
rect 21000 -247 25000 -230
rect 21000 -273 21119 -247
rect 21145 -273 24852 -247
rect 24878 -273 25000 -247
rect 21000 -350 25000 -273
rect 21000 -376 21307 -350
rect 21333 -376 21467 -350
rect 21493 -376 21627 -350
rect 21653 -376 21787 -350
rect 21813 -376 21947 -350
rect 21973 -376 22107 -350
rect 22133 -376 22267 -350
rect 22293 -376 22427 -350
rect 22453 -376 22587 -350
rect 22613 -376 22747 -350
rect 22773 -376 22907 -350
rect 22933 -376 23067 -350
rect 23093 -376 23227 -350
rect 23253 -376 23387 -350
rect 23413 -376 23547 -350
rect 23573 -376 23707 -350
rect 23733 -376 23867 -350
rect 23893 -376 24027 -350
rect 24053 -376 24187 -350
rect 24213 -376 24347 -350
rect 24373 -376 24507 -350
rect 24533 -376 24667 -350
rect 24693 -376 25000 -350
rect 21000 -500 25000 -376
rect 19240 -575 19300 -570
rect 19240 -745 19245 -575
rect 19290 -745 19300 -575
rect 19595 -575 19650 -570
rect 19430 -630 19490 -625
rect 19430 -690 19435 -630
rect 19485 -690 19490 -630
rect 19430 -695 19490 -690
rect 19240 -750 19300 -745
rect 19595 -745 19600 -575
rect 19645 -745 19650 -575
rect 19595 -750 19650 -745
rect 20030 -1140 20070 -1135
rect 20030 -1170 20035 -1140
rect 20065 -1170 20070 -1140
rect 20030 -1175 20070 -1170
rect 20030 -1225 20050 -1175
rect 20065 -1210 20105 -1205
rect 20065 -1240 20070 -1210
rect 20100 -1240 20105 -1210
rect 20065 -1245 20105 -1240
rect 16200 -2050 16250 -1950
rect 16350 -2050 16400 -1950
rect 16150 -2180 16155 -2140
rect 16225 -2180 16230 -2140
rect 16290 -2180 16295 -2140
rect 16365 -2180 16370 -2140
rect 16200 -2400 16250 -2300
rect 16350 -2400 16400 -2300
rect 11600 -3700 11650 -3600
rect 11750 -3700 11800 -3600
rect 11630 -3860 11635 -3820
rect 11705 -3860 11710 -3820
rect 11770 -3860 11775 -3820
rect 11845 -3860 11850 -3820
rect 11600 -4050 11650 -3950
rect 11750 -4050 11800 -3950
rect 8195 -4760 8235 -4755
rect 8195 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8195 -4795 8235 -4790
rect 8250 -4825 8270 -4775
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 8350 -5255 8405 -5250
rect 8350 -5425 8355 -5255
rect 8400 -5425 8405 -5255
rect 8700 -5255 8760 -5250
rect 8510 -5310 8570 -5305
rect 8510 -5370 8515 -5310
rect 8565 -5370 8570 -5310
rect 8510 -5375 8570 -5370
rect 8350 -5430 8405 -5425
rect 8700 -5425 8710 -5255
rect 8755 -5425 8760 -5255
rect 8700 -5430 8760 -5425
rect 3000 -5624 7000 -5500
rect 3000 -5650 3307 -5624
rect 3333 -5650 3467 -5624
rect 3493 -5650 3627 -5624
rect 3653 -5650 3787 -5624
rect 3813 -5650 3947 -5624
rect 3973 -5650 4107 -5624
rect 4133 -5650 4267 -5624
rect 4293 -5650 4427 -5624
rect 4453 -5650 4587 -5624
rect 4613 -5650 4747 -5624
rect 4773 -5650 4907 -5624
rect 4933 -5650 5067 -5624
rect 5093 -5650 5227 -5624
rect 5253 -5650 5387 -5624
rect 5413 -5650 5547 -5624
rect 5573 -5650 5707 -5624
rect 5733 -5650 5867 -5624
rect 5893 -5650 6027 -5624
rect 6053 -5650 6187 -5624
rect 6213 -5650 6347 -5624
rect 6373 -5650 6507 -5624
rect 6533 -5650 6667 -5624
rect 6693 -5650 7000 -5624
rect 3000 -5727 7000 -5650
rect 3000 -5753 3122 -5727
rect 3148 -5753 6855 -5727
rect 6881 -5753 7000 -5727
rect 3000 -5770 7000 -5753
rect 3000 -5887 3270 -5770
rect 3000 -5913 3122 -5887
rect 3148 -5913 3270 -5887
rect 3000 -6047 3270 -5913
rect 3000 -6073 3122 -6047
rect 3148 -6073 3270 -6047
rect 3000 -6207 3270 -6073
rect 3000 -6233 3122 -6207
rect 3148 -6233 3270 -6207
rect 3000 -6367 3270 -6233
rect 3000 -6393 3122 -6367
rect 3148 -6393 3270 -6367
rect 3000 -6527 3270 -6393
rect 3000 -6553 3122 -6527
rect 3148 -6553 3270 -6527
rect 3000 -6687 3270 -6553
rect 3000 -6713 3122 -6687
rect 3148 -6713 3270 -6687
rect 3000 -6847 3270 -6713
rect 3000 -6873 3122 -6847
rect 3148 -6873 3270 -6847
rect 3000 -7007 3270 -6873
rect 3000 -7033 3122 -7007
rect 3148 -7033 3270 -7007
rect 3000 -7167 3270 -7033
rect 3000 -7193 3122 -7167
rect 3148 -7193 3270 -7167
rect 3000 -7327 3270 -7193
rect 3000 -7353 3122 -7327
rect 3148 -7353 3270 -7327
rect 3000 -7487 3270 -7353
rect 3000 -7513 3122 -7487
rect 3148 -7513 3270 -7487
rect 3000 -7647 3270 -7513
rect 3000 -7673 3122 -7647
rect 3148 -7673 3270 -7647
rect 3000 -7807 3270 -7673
rect 3000 -7833 3122 -7807
rect 3148 -7833 3270 -7807
rect 3000 -7967 3270 -7833
rect 3000 -7993 3122 -7967
rect 3148 -7993 3270 -7967
rect 3000 -8127 3270 -7993
rect 3000 -8153 3122 -8127
rect 3148 -8153 3270 -8127
rect 3000 -8287 3270 -8153
rect 3000 -8313 3122 -8287
rect 3148 -8313 3270 -8287
rect 3000 -8447 3270 -8313
rect 3000 -8473 3122 -8447
rect 3148 -8473 3270 -8447
rect 3000 -8607 3270 -8473
rect 3000 -8633 3122 -8607
rect 3148 -8633 3270 -8607
rect 3000 -8767 3270 -8633
rect 3000 -8793 3122 -8767
rect 3148 -8793 3270 -8767
rect 3000 -8927 3270 -8793
rect 3000 -8953 3122 -8927
rect 3148 -8953 3270 -8927
rect 3000 -9087 3270 -8953
rect 3000 -9113 3122 -9087
rect 3148 -9113 3270 -9087
rect 3000 -9230 3270 -9113
rect 6730 -5887 7000 -5770
rect 6730 -5913 6855 -5887
rect 6881 -5913 7000 -5887
rect 6730 -6047 7000 -5913
rect 6730 -6073 6855 -6047
rect 6881 -6073 7000 -6047
rect 6730 -6207 7000 -6073
rect 6730 -6233 6855 -6207
rect 6881 -6233 7000 -6207
rect 6730 -6367 7000 -6233
rect 6730 -6393 6855 -6367
rect 6881 -6393 7000 -6367
rect 6730 -6527 7000 -6393
rect 6730 -6553 6855 -6527
rect 6881 -6553 7000 -6527
rect 6730 -6687 7000 -6553
rect 6730 -6713 6855 -6687
rect 6881 -6713 7000 -6687
rect 6730 -6847 7000 -6713
rect 6730 -6873 6855 -6847
rect 6881 -6873 7000 -6847
rect 6730 -7007 7000 -6873
rect 6730 -7033 6855 -7007
rect 6881 -7033 7000 -7007
rect 6730 -7167 7000 -7033
rect 6730 -7193 6855 -7167
rect 6881 -7193 7000 -7167
rect 6730 -7327 7000 -7193
rect 6730 -7353 6855 -7327
rect 6881 -7353 7000 -7327
rect 6730 -7487 7000 -7353
rect 6730 -7513 6855 -7487
rect 6881 -7513 7000 -7487
rect 6730 -7647 7000 -7513
rect 6730 -7673 6855 -7647
rect 6881 -7673 7000 -7647
rect 6730 -7807 7000 -7673
rect 6730 -7833 6855 -7807
rect 6881 -7833 7000 -7807
rect 6730 -7967 7000 -7833
rect 6730 -7993 6855 -7967
rect 6881 -7993 7000 -7967
rect 6730 -8127 7000 -7993
rect 6730 -8153 6855 -8127
rect 6881 -8153 7000 -8127
rect 6730 -8287 7000 -8153
rect 6730 -8313 6855 -8287
rect 6881 -8313 7000 -8287
rect 6730 -8447 7000 -8313
rect 6730 -8473 6855 -8447
rect 6881 -8473 7000 -8447
rect 6730 -8607 7000 -8473
rect 6730 -8633 6855 -8607
rect 6881 -8633 7000 -8607
rect 6730 -8767 7000 -8633
rect 6730 -8793 6855 -8767
rect 6881 -8793 7000 -8767
rect 6730 -8927 7000 -8793
rect 6730 -8953 6855 -8927
rect 6881 -8953 7000 -8927
rect 6730 -9087 7000 -8953
rect 6730 -9113 6855 -9087
rect 6881 -9113 7000 -9087
rect 6730 -9230 7000 -9113
rect 3000 -9247 7000 -9230
rect 3000 -9273 3122 -9247
rect 3148 -9273 6855 -9247
rect 6881 -9273 7000 -9247
rect 3000 -9352 7000 -9273
rect 3000 -9378 3307 -9352
rect 3333 -9378 3467 -9352
rect 3493 -9378 3627 -9352
rect 3653 -9378 3787 -9352
rect 3813 -9378 3947 -9352
rect 3973 -9378 4107 -9352
rect 4133 -9378 4267 -9352
rect 4293 -9378 4427 -9352
rect 4453 -9378 4587 -9352
rect 4613 -9378 4747 -9352
rect 4773 -9378 4907 -9352
rect 4933 -9378 5067 -9352
rect 5093 -9378 5227 -9352
rect 5253 -9378 5387 -9352
rect 5413 -9378 5547 -9352
rect 5573 -9378 5707 -9352
rect 5733 -9378 5867 -9352
rect 5893 -9378 6027 -9352
rect 6053 -9378 6187 -9352
rect 6213 -9378 6347 -9352
rect 6373 -9378 6507 -9352
rect 6533 -9378 6667 -9352
rect 6693 -9378 7000 -9352
rect 3000 -9500 7000 -9378
rect 9000 -5624 13000 -5500
rect 9000 -5650 9307 -5624
rect 9333 -5650 9467 -5624
rect 9493 -5650 9627 -5624
rect 9653 -5650 9787 -5624
rect 9813 -5650 9947 -5624
rect 9973 -5650 10107 -5624
rect 10133 -5650 10267 -5624
rect 10293 -5650 10427 -5624
rect 10453 -5650 10587 -5624
rect 10613 -5650 10747 -5624
rect 10773 -5650 10907 -5624
rect 10933 -5650 11067 -5624
rect 11093 -5650 11227 -5624
rect 11253 -5650 11387 -5624
rect 11413 -5650 11547 -5624
rect 11573 -5650 11707 -5624
rect 11733 -5650 11867 -5624
rect 11893 -5650 12027 -5624
rect 12053 -5650 12187 -5624
rect 12213 -5650 12347 -5624
rect 12373 -5650 12507 -5624
rect 12533 -5650 12667 -5624
rect 12693 -5650 13000 -5624
rect 9000 -5727 13000 -5650
rect 9000 -5753 9122 -5727
rect 9148 -5753 12855 -5727
rect 12881 -5753 13000 -5727
rect 9000 -5770 13000 -5753
rect 9000 -5887 9270 -5770
rect 9000 -5913 9122 -5887
rect 9148 -5913 9270 -5887
rect 9000 -6047 9270 -5913
rect 9000 -6073 9122 -6047
rect 9148 -6073 9270 -6047
rect 9000 -6207 9270 -6073
rect 9000 -6233 9122 -6207
rect 9148 -6233 9270 -6207
rect 9000 -6367 9270 -6233
rect 9000 -6393 9122 -6367
rect 9148 -6393 9270 -6367
rect 9000 -6527 9270 -6393
rect 9000 -6553 9122 -6527
rect 9148 -6553 9270 -6527
rect 9000 -6687 9270 -6553
rect 9000 -6713 9122 -6687
rect 9148 -6713 9270 -6687
rect 9000 -6847 9270 -6713
rect 9000 -6873 9122 -6847
rect 9148 -6873 9270 -6847
rect 9000 -7007 9270 -6873
rect 9000 -7033 9122 -7007
rect 9148 -7033 9270 -7007
rect 9000 -7167 9270 -7033
rect 9000 -7193 9122 -7167
rect 9148 -7193 9270 -7167
rect 9000 -7327 9270 -7193
rect 9000 -7353 9122 -7327
rect 9148 -7353 9270 -7327
rect 9000 -7487 9270 -7353
rect 9000 -7513 9122 -7487
rect 9148 -7513 9270 -7487
rect 9000 -7647 9270 -7513
rect 9000 -7673 9122 -7647
rect 9148 -7673 9270 -7647
rect 9000 -7807 9270 -7673
rect 9000 -7833 9122 -7807
rect 9148 -7833 9270 -7807
rect 9000 -7967 9270 -7833
rect 9000 -7993 9122 -7967
rect 9148 -7993 9270 -7967
rect 9000 -8127 9270 -7993
rect 9000 -8153 9122 -8127
rect 9148 -8153 9270 -8127
rect 9000 -8287 9270 -8153
rect 9000 -8313 9122 -8287
rect 9148 -8313 9270 -8287
rect 9000 -8447 9270 -8313
rect 9000 -8473 9122 -8447
rect 9148 -8473 9270 -8447
rect 9000 -8607 9270 -8473
rect 9000 -8633 9122 -8607
rect 9148 -8633 9270 -8607
rect 9000 -8767 9270 -8633
rect 9000 -8793 9122 -8767
rect 9148 -8793 9270 -8767
rect 9000 -8927 9270 -8793
rect 9000 -8953 9122 -8927
rect 9148 -8953 9270 -8927
rect 9000 -9087 9270 -8953
rect 9000 -9113 9122 -9087
rect 9148 -9113 9270 -9087
rect 9000 -9230 9270 -9113
rect 12730 -5887 13000 -5770
rect 12730 -5913 12855 -5887
rect 12881 -5913 13000 -5887
rect 12730 -6047 13000 -5913
rect 12730 -6073 12855 -6047
rect 12881 -6073 13000 -6047
rect 12730 -6207 13000 -6073
rect 12730 -6233 12855 -6207
rect 12881 -6233 13000 -6207
rect 12730 -6367 13000 -6233
rect 12730 -6393 12855 -6367
rect 12881 -6393 13000 -6367
rect 12730 -6527 13000 -6393
rect 12730 -6553 12855 -6527
rect 12881 -6553 13000 -6527
rect 12730 -6687 13000 -6553
rect 12730 -6713 12855 -6687
rect 12881 -6713 13000 -6687
rect 12730 -6847 13000 -6713
rect 12730 -6873 12855 -6847
rect 12881 -6873 13000 -6847
rect 12730 -7007 13000 -6873
rect 12730 -7033 12855 -7007
rect 12881 -7033 13000 -7007
rect 12730 -7167 13000 -7033
rect 12730 -7193 12855 -7167
rect 12881 -7193 13000 -7167
rect 12730 -7327 13000 -7193
rect 12730 -7353 12855 -7327
rect 12881 -7353 13000 -7327
rect 12730 -7487 13000 -7353
rect 12730 -7513 12855 -7487
rect 12881 -7513 13000 -7487
rect 12730 -7647 13000 -7513
rect 12730 -7673 12855 -7647
rect 12881 -7673 13000 -7647
rect 12730 -7807 13000 -7673
rect 12730 -7833 12855 -7807
rect 12881 -7833 13000 -7807
rect 12730 -7967 13000 -7833
rect 12730 -7993 12855 -7967
rect 12881 -7993 13000 -7967
rect 12730 -8127 13000 -7993
rect 12730 -8153 12855 -8127
rect 12881 -8153 13000 -8127
rect 12730 -8287 13000 -8153
rect 12730 -8313 12855 -8287
rect 12881 -8313 13000 -8287
rect 12730 -8447 13000 -8313
rect 12730 -8473 12855 -8447
rect 12881 -8473 13000 -8447
rect 12730 -8607 13000 -8473
rect 12730 -8633 12855 -8607
rect 12881 -8633 13000 -8607
rect 12730 -8767 13000 -8633
rect 12730 -8793 12855 -8767
rect 12881 -8793 13000 -8767
rect 12730 -8927 13000 -8793
rect 12730 -8953 12855 -8927
rect 12881 -8953 13000 -8927
rect 12730 -9087 13000 -8953
rect 12730 -9113 12855 -9087
rect 12881 -9113 13000 -9087
rect 12730 -9230 13000 -9113
rect 9000 -9247 13000 -9230
rect 9000 -9273 9122 -9247
rect 9148 -9273 12855 -9247
rect 12881 -9273 13000 -9247
rect 9000 -9352 13000 -9273
rect 9000 -9378 9307 -9352
rect 9333 -9378 9467 -9352
rect 9493 -9378 9627 -9352
rect 9653 -9378 9787 -9352
rect 9813 -9378 9947 -9352
rect 9973 -9378 10107 -9352
rect 10133 -9378 10267 -9352
rect 10293 -9378 10427 -9352
rect 10453 -9378 10587 -9352
rect 10613 -9378 10747 -9352
rect 10773 -9378 10907 -9352
rect 10933 -9378 11067 -9352
rect 11093 -9378 11227 -9352
rect 11253 -9378 11387 -9352
rect 11413 -9378 11547 -9352
rect 11573 -9378 11707 -9352
rect 11733 -9378 11867 -9352
rect 11893 -9378 12027 -9352
rect 12053 -9378 12187 -9352
rect 12213 -9378 12347 -9352
rect 12373 -9378 12507 -9352
rect 12533 -9378 12667 -9352
rect 12693 -9378 13000 -9352
rect 9000 -9500 13000 -9378
rect 15000 -5624 19000 -5500
rect 15000 -5650 15307 -5624
rect 15333 -5650 15467 -5624
rect 15493 -5650 15627 -5624
rect 15653 -5650 15787 -5624
rect 15813 -5650 15947 -5624
rect 15973 -5650 16107 -5624
rect 16133 -5650 16267 -5624
rect 16293 -5650 16427 -5624
rect 16453 -5650 16587 -5624
rect 16613 -5650 16747 -5624
rect 16773 -5650 16907 -5624
rect 16933 -5650 17067 -5624
rect 17093 -5650 17227 -5624
rect 17253 -5650 17387 -5624
rect 17413 -5650 17547 -5624
rect 17573 -5650 17707 -5624
rect 17733 -5650 17867 -5624
rect 17893 -5650 18027 -5624
rect 18053 -5650 18187 -5624
rect 18213 -5650 18347 -5624
rect 18373 -5650 18507 -5624
rect 18533 -5650 18667 -5624
rect 18693 -5650 19000 -5624
rect 15000 -5727 19000 -5650
rect 15000 -5753 15122 -5727
rect 15148 -5753 18855 -5727
rect 18881 -5753 19000 -5727
rect 15000 -5770 19000 -5753
rect 15000 -5887 15270 -5770
rect 15000 -5913 15122 -5887
rect 15148 -5913 15270 -5887
rect 15000 -6047 15270 -5913
rect 15000 -6073 15122 -6047
rect 15148 -6073 15270 -6047
rect 15000 -6207 15270 -6073
rect 15000 -6233 15122 -6207
rect 15148 -6233 15270 -6207
rect 15000 -6367 15270 -6233
rect 15000 -6393 15122 -6367
rect 15148 -6393 15270 -6367
rect 15000 -6527 15270 -6393
rect 15000 -6553 15122 -6527
rect 15148 -6553 15270 -6527
rect 15000 -6687 15270 -6553
rect 15000 -6713 15122 -6687
rect 15148 -6713 15270 -6687
rect 15000 -6847 15270 -6713
rect 15000 -6873 15122 -6847
rect 15148 -6873 15270 -6847
rect 15000 -7007 15270 -6873
rect 15000 -7033 15122 -7007
rect 15148 -7033 15270 -7007
rect 15000 -7167 15270 -7033
rect 15000 -7193 15122 -7167
rect 15148 -7193 15270 -7167
rect 15000 -7327 15270 -7193
rect 15000 -7353 15122 -7327
rect 15148 -7353 15270 -7327
rect 15000 -7487 15270 -7353
rect 15000 -7513 15122 -7487
rect 15148 -7513 15270 -7487
rect 15000 -7647 15270 -7513
rect 15000 -7673 15122 -7647
rect 15148 -7673 15270 -7647
rect 15000 -7807 15270 -7673
rect 15000 -7833 15122 -7807
rect 15148 -7833 15270 -7807
rect 15000 -7967 15270 -7833
rect 15000 -7993 15122 -7967
rect 15148 -7993 15270 -7967
rect 15000 -8127 15270 -7993
rect 15000 -8153 15122 -8127
rect 15148 -8153 15270 -8127
rect 15000 -8287 15270 -8153
rect 15000 -8313 15122 -8287
rect 15148 -8313 15270 -8287
rect 15000 -8447 15270 -8313
rect 15000 -8473 15122 -8447
rect 15148 -8473 15270 -8447
rect 15000 -8607 15270 -8473
rect 15000 -8633 15122 -8607
rect 15148 -8633 15270 -8607
rect 15000 -8767 15270 -8633
rect 15000 -8793 15122 -8767
rect 15148 -8793 15270 -8767
rect 15000 -8927 15270 -8793
rect 15000 -8953 15122 -8927
rect 15148 -8953 15270 -8927
rect 15000 -9087 15270 -8953
rect 15000 -9113 15122 -9087
rect 15148 -9113 15270 -9087
rect 15000 -9230 15270 -9113
rect 18730 -5887 19000 -5770
rect 18730 -5913 18855 -5887
rect 18881 -5913 19000 -5887
rect 18730 -6047 19000 -5913
rect 18730 -6073 18855 -6047
rect 18881 -6073 19000 -6047
rect 18730 -6207 19000 -6073
rect 18730 -6233 18855 -6207
rect 18881 -6233 19000 -6207
rect 18730 -6367 19000 -6233
rect 18730 -6393 18855 -6367
rect 18881 -6393 19000 -6367
rect 18730 -6527 19000 -6393
rect 18730 -6553 18855 -6527
rect 18881 -6553 19000 -6527
rect 18730 -6687 19000 -6553
rect 18730 -6713 18855 -6687
rect 18881 -6713 19000 -6687
rect 18730 -6847 19000 -6713
rect 18730 -6873 18855 -6847
rect 18881 -6873 19000 -6847
rect 18730 -7007 19000 -6873
rect 18730 -7033 18855 -7007
rect 18881 -7033 19000 -7007
rect 18730 -7167 19000 -7033
rect 18730 -7193 18855 -7167
rect 18881 -7193 19000 -7167
rect 18730 -7327 19000 -7193
rect 18730 -7353 18855 -7327
rect 18881 -7353 19000 -7327
rect 18730 -7487 19000 -7353
rect 18730 -7513 18855 -7487
rect 18881 -7513 19000 -7487
rect 18730 -7647 19000 -7513
rect 18730 -7673 18855 -7647
rect 18881 -7673 19000 -7647
rect 18730 -7807 19000 -7673
rect 18730 -7833 18855 -7807
rect 18881 -7833 19000 -7807
rect 18730 -7967 19000 -7833
rect 18730 -7993 18855 -7967
rect 18881 -7993 19000 -7967
rect 18730 -8127 19000 -7993
rect 18730 -8153 18855 -8127
rect 18881 -8153 19000 -8127
rect 18730 -8287 19000 -8153
rect 18730 -8313 18855 -8287
rect 18881 -8313 19000 -8287
rect 18730 -8447 19000 -8313
rect 18730 -8473 18855 -8447
rect 18881 -8473 19000 -8447
rect 18730 -8607 19000 -8473
rect 18730 -8633 18855 -8607
rect 18881 -8633 19000 -8607
rect 18730 -8767 19000 -8633
rect 18730 -8793 18855 -8767
rect 18881 -8793 19000 -8767
rect 18730 -8927 19000 -8793
rect 18730 -8953 18855 -8927
rect 18881 -8953 19000 -8927
rect 18730 -9087 19000 -8953
rect 18730 -9113 18855 -9087
rect 18881 -9113 19000 -9087
rect 18730 -9230 19000 -9113
rect 15000 -9247 19000 -9230
rect 15000 -9273 15122 -9247
rect 15148 -9273 18855 -9247
rect 18881 -9273 19000 -9247
rect 15000 -9352 19000 -9273
rect 15000 -9378 15307 -9352
rect 15333 -9378 15467 -9352
rect 15493 -9378 15627 -9352
rect 15653 -9378 15787 -9352
rect 15813 -9378 15947 -9352
rect 15973 -9378 16107 -9352
rect 16133 -9378 16267 -9352
rect 16293 -9378 16427 -9352
rect 16453 -9378 16587 -9352
rect 16613 -9378 16747 -9352
rect 16773 -9378 16907 -9352
rect 16933 -9378 17067 -9352
rect 17093 -9378 17227 -9352
rect 17253 -9378 17387 -9352
rect 17413 -9378 17547 -9352
rect 17573 -9378 17707 -9352
rect 17733 -9378 17867 -9352
rect 17893 -9378 18027 -9352
rect 18053 -9378 18187 -9352
rect 18213 -9378 18347 -9352
rect 18373 -9378 18507 -9352
rect 18533 -9378 18667 -9352
rect 18693 -9378 19000 -9352
rect 15000 -9500 19000 -9378
rect 21000 -5624 25000 -5500
rect 21000 -5650 21307 -5624
rect 21333 -5650 21467 -5624
rect 21493 -5650 21627 -5624
rect 21653 -5650 21787 -5624
rect 21813 -5650 21947 -5624
rect 21973 -5650 22107 -5624
rect 22133 -5650 22267 -5624
rect 22293 -5650 22427 -5624
rect 22453 -5650 22587 -5624
rect 22613 -5650 22747 -5624
rect 22773 -5650 22907 -5624
rect 22933 -5650 23067 -5624
rect 23093 -5650 23227 -5624
rect 23253 -5650 23387 -5624
rect 23413 -5650 23547 -5624
rect 23573 -5650 23707 -5624
rect 23733 -5650 23867 -5624
rect 23893 -5650 24027 -5624
rect 24053 -5650 24187 -5624
rect 24213 -5650 24347 -5624
rect 24373 -5650 24507 -5624
rect 24533 -5650 24667 -5624
rect 24693 -5650 25000 -5624
rect 21000 -5727 25000 -5650
rect 21000 -5753 21122 -5727
rect 21148 -5753 24855 -5727
rect 24881 -5753 25000 -5727
rect 21000 -5770 25000 -5753
rect 21000 -5887 21270 -5770
rect 21000 -5913 21122 -5887
rect 21148 -5913 21270 -5887
rect 21000 -6047 21270 -5913
rect 21000 -6073 21122 -6047
rect 21148 -6073 21270 -6047
rect 21000 -6207 21270 -6073
rect 21000 -6233 21122 -6207
rect 21148 -6233 21270 -6207
rect 21000 -6367 21270 -6233
rect 21000 -6393 21122 -6367
rect 21148 -6393 21270 -6367
rect 21000 -6527 21270 -6393
rect 21000 -6553 21122 -6527
rect 21148 -6553 21270 -6527
rect 21000 -6687 21270 -6553
rect 21000 -6713 21122 -6687
rect 21148 -6713 21270 -6687
rect 21000 -6847 21270 -6713
rect 21000 -6873 21122 -6847
rect 21148 -6873 21270 -6847
rect 21000 -7007 21270 -6873
rect 21000 -7033 21122 -7007
rect 21148 -7033 21270 -7007
rect 21000 -7167 21270 -7033
rect 21000 -7193 21122 -7167
rect 21148 -7193 21270 -7167
rect 21000 -7327 21270 -7193
rect 21000 -7353 21122 -7327
rect 21148 -7353 21270 -7327
rect 21000 -7487 21270 -7353
rect 21000 -7513 21122 -7487
rect 21148 -7513 21270 -7487
rect 21000 -7647 21270 -7513
rect 21000 -7673 21122 -7647
rect 21148 -7673 21270 -7647
rect 21000 -7807 21270 -7673
rect 21000 -7833 21122 -7807
rect 21148 -7833 21270 -7807
rect 21000 -7967 21270 -7833
rect 21000 -7993 21122 -7967
rect 21148 -7993 21270 -7967
rect 21000 -8127 21270 -7993
rect 21000 -8153 21122 -8127
rect 21148 -8153 21270 -8127
rect 21000 -8287 21270 -8153
rect 21000 -8313 21122 -8287
rect 21148 -8313 21270 -8287
rect 21000 -8447 21270 -8313
rect 21000 -8473 21122 -8447
rect 21148 -8473 21270 -8447
rect 21000 -8607 21270 -8473
rect 21000 -8633 21122 -8607
rect 21148 -8633 21270 -8607
rect 21000 -8767 21270 -8633
rect 21000 -8793 21122 -8767
rect 21148 -8793 21270 -8767
rect 21000 -8927 21270 -8793
rect 21000 -8953 21122 -8927
rect 21148 -8953 21270 -8927
rect 21000 -9087 21270 -8953
rect 21000 -9113 21122 -9087
rect 21148 -9113 21270 -9087
rect 21000 -9230 21270 -9113
rect 24730 -5887 25000 -5770
rect 24730 -5913 24855 -5887
rect 24881 -5913 25000 -5887
rect 24730 -6047 25000 -5913
rect 24730 -6073 24855 -6047
rect 24881 -6073 25000 -6047
rect 24730 -6207 25000 -6073
rect 24730 -6233 24855 -6207
rect 24881 -6233 25000 -6207
rect 24730 -6367 25000 -6233
rect 24730 -6393 24855 -6367
rect 24881 -6393 25000 -6367
rect 24730 -6527 25000 -6393
rect 24730 -6553 24855 -6527
rect 24881 -6553 25000 -6527
rect 24730 -6687 25000 -6553
rect 24730 -6713 24855 -6687
rect 24881 -6713 25000 -6687
rect 24730 -6847 25000 -6713
rect 24730 -6873 24855 -6847
rect 24881 -6873 25000 -6847
rect 24730 -7007 25000 -6873
rect 24730 -7033 24855 -7007
rect 24881 -7033 25000 -7007
rect 24730 -7167 25000 -7033
rect 24730 -7193 24855 -7167
rect 24881 -7193 25000 -7167
rect 24730 -7327 25000 -7193
rect 24730 -7353 24855 -7327
rect 24881 -7353 25000 -7327
rect 24730 -7487 25000 -7353
rect 24730 -7513 24855 -7487
rect 24881 -7513 25000 -7487
rect 24730 -7647 25000 -7513
rect 24730 -7673 24855 -7647
rect 24881 -7673 25000 -7647
rect 24730 -7807 25000 -7673
rect 24730 -7833 24855 -7807
rect 24881 -7833 25000 -7807
rect 24730 -7967 25000 -7833
rect 24730 -7993 24855 -7967
rect 24881 -7993 25000 -7967
rect 24730 -8127 25000 -7993
rect 24730 -8153 24855 -8127
rect 24881 -8153 25000 -8127
rect 24730 -8287 25000 -8153
rect 24730 -8313 24855 -8287
rect 24881 -8313 25000 -8287
rect 24730 -8447 25000 -8313
rect 24730 -8473 24855 -8447
rect 24881 -8473 25000 -8447
rect 24730 -8607 25000 -8473
rect 24730 -8633 24855 -8607
rect 24881 -8633 25000 -8607
rect 24730 -8767 25000 -8633
rect 24730 -8793 24855 -8767
rect 24881 -8793 25000 -8767
rect 24730 -8927 25000 -8793
rect 24730 -8953 24855 -8927
rect 24881 -8953 25000 -8927
rect 24730 -9087 25000 -8953
rect 24730 -9113 24855 -9087
rect 24881 -9113 25000 -9087
rect 24730 -9230 25000 -9113
rect 21000 -9247 25000 -9230
rect 21000 -9273 21122 -9247
rect 21148 -9273 24855 -9247
rect 24881 -9273 25000 -9247
rect 21000 -9352 25000 -9273
rect 21000 -9378 21307 -9352
rect 21333 -9378 21467 -9352
rect 21493 -9378 21627 -9352
rect 21653 -9378 21787 -9352
rect 21813 -9378 21947 -9352
rect 21973 -9378 22107 -9352
rect 22133 -9378 22267 -9352
rect 22293 -9378 22427 -9352
rect 22453 -9378 22587 -9352
rect 22613 -9378 22747 -9352
rect 22773 -9378 22907 -9352
rect 22933 -9378 23067 -9352
rect 23093 -9378 23227 -9352
rect 23253 -9378 23387 -9352
rect 23413 -9378 23547 -9352
rect 23573 -9378 23707 -9352
rect 23733 -9378 23867 -9352
rect 23893 -9378 24027 -9352
rect 24053 -9378 24187 -9352
rect 24213 -9378 24347 -9352
rect 24373 -9378 24507 -9352
rect 24533 -9378 24667 -9352
rect 24693 -9378 25000 -9352
rect 21000 -9500 25000 -9378
rect 3000 -11624 7000 -11500
rect 3000 -11650 3307 -11624
rect 3333 -11650 3467 -11624
rect 3493 -11650 3627 -11624
rect 3653 -11650 3787 -11624
rect 3813 -11650 3947 -11624
rect 3973 -11650 4107 -11624
rect 4133 -11650 4267 -11624
rect 4293 -11650 4427 -11624
rect 4453 -11650 4587 -11624
rect 4613 -11650 4747 -11624
rect 4773 -11650 4907 -11624
rect 4933 -11650 5067 -11624
rect 5093 -11650 5227 -11624
rect 5253 -11650 5387 -11624
rect 5413 -11650 5547 -11624
rect 5573 -11650 5707 -11624
rect 5733 -11650 5867 -11624
rect 5893 -11650 6027 -11624
rect 6053 -11650 6187 -11624
rect 6213 -11650 6347 -11624
rect 6373 -11650 6507 -11624
rect 6533 -11650 6667 -11624
rect 6693 -11650 7000 -11624
rect 3000 -11727 7000 -11650
rect 3000 -11753 3122 -11727
rect 3148 -11753 6855 -11727
rect 6881 -11753 7000 -11727
rect 3000 -11770 7000 -11753
rect 3000 -11887 3270 -11770
rect 3000 -11913 3122 -11887
rect 3148 -11913 3270 -11887
rect 3000 -12047 3270 -11913
rect 3000 -12073 3122 -12047
rect 3148 -12073 3270 -12047
rect 3000 -12207 3270 -12073
rect 3000 -12233 3122 -12207
rect 3148 -12233 3270 -12207
rect 3000 -12367 3270 -12233
rect 3000 -12393 3122 -12367
rect 3148 -12393 3270 -12367
rect 3000 -12527 3270 -12393
rect 3000 -12553 3122 -12527
rect 3148 -12553 3270 -12527
rect 3000 -12687 3270 -12553
rect 3000 -12713 3122 -12687
rect 3148 -12713 3270 -12687
rect 3000 -12847 3270 -12713
rect 3000 -12873 3122 -12847
rect 3148 -12873 3270 -12847
rect 3000 -13007 3270 -12873
rect 3000 -13033 3122 -13007
rect 3148 -13033 3270 -13007
rect 3000 -13167 3270 -13033
rect 3000 -13193 3122 -13167
rect 3148 -13193 3270 -13167
rect 3000 -13327 3270 -13193
rect 3000 -13353 3122 -13327
rect 3148 -13353 3270 -13327
rect 3000 -13487 3270 -13353
rect 3000 -13513 3122 -13487
rect 3148 -13513 3270 -13487
rect 3000 -13647 3270 -13513
rect 3000 -13673 3122 -13647
rect 3148 -13673 3270 -13647
rect 3000 -13807 3270 -13673
rect 3000 -13833 3122 -13807
rect 3148 -13833 3270 -13807
rect 3000 -13967 3270 -13833
rect 3000 -13993 3122 -13967
rect 3148 -13993 3270 -13967
rect 3000 -14127 3270 -13993
rect 3000 -14153 3122 -14127
rect 3148 -14153 3270 -14127
rect 3000 -14287 3270 -14153
rect 3000 -14313 3122 -14287
rect 3148 -14313 3270 -14287
rect 3000 -14447 3270 -14313
rect 3000 -14473 3122 -14447
rect 3148 -14473 3270 -14447
rect 3000 -14607 3270 -14473
rect 3000 -14633 3122 -14607
rect 3148 -14633 3270 -14607
rect 3000 -14767 3270 -14633
rect 3000 -14793 3122 -14767
rect 3148 -14793 3270 -14767
rect 3000 -14927 3270 -14793
rect 3000 -14953 3122 -14927
rect 3148 -14953 3270 -14927
rect 3000 -15087 3270 -14953
rect 3000 -15113 3122 -15087
rect 3148 -15113 3270 -15087
rect 3000 -15230 3270 -15113
rect 6730 -11887 7000 -11770
rect 6730 -11913 6855 -11887
rect 6881 -11913 7000 -11887
rect 6730 -12047 7000 -11913
rect 6730 -12073 6855 -12047
rect 6881 -12073 7000 -12047
rect 6730 -12207 7000 -12073
rect 6730 -12233 6855 -12207
rect 6881 -12233 7000 -12207
rect 6730 -12367 7000 -12233
rect 6730 -12393 6855 -12367
rect 6881 -12393 7000 -12367
rect 6730 -12527 7000 -12393
rect 6730 -12553 6855 -12527
rect 6881 -12553 7000 -12527
rect 6730 -12687 7000 -12553
rect 6730 -12713 6855 -12687
rect 6881 -12713 7000 -12687
rect 6730 -12847 7000 -12713
rect 6730 -12873 6855 -12847
rect 6881 -12873 7000 -12847
rect 6730 -13007 7000 -12873
rect 6730 -13033 6855 -13007
rect 6881 -13033 7000 -13007
rect 6730 -13167 7000 -13033
rect 6730 -13193 6855 -13167
rect 6881 -13193 7000 -13167
rect 6730 -13327 7000 -13193
rect 6730 -13353 6855 -13327
rect 6881 -13353 7000 -13327
rect 6730 -13487 7000 -13353
rect 6730 -13513 6855 -13487
rect 6881 -13513 7000 -13487
rect 6730 -13647 7000 -13513
rect 6730 -13673 6855 -13647
rect 6881 -13673 7000 -13647
rect 6730 -13807 7000 -13673
rect 6730 -13833 6855 -13807
rect 6881 -13833 7000 -13807
rect 6730 -13967 7000 -13833
rect 6730 -13993 6855 -13967
rect 6881 -13993 7000 -13967
rect 6730 -14127 7000 -13993
rect 6730 -14153 6855 -14127
rect 6881 -14153 7000 -14127
rect 6730 -14287 7000 -14153
rect 6730 -14313 6855 -14287
rect 6881 -14313 7000 -14287
rect 6730 -14447 7000 -14313
rect 6730 -14473 6855 -14447
rect 6881 -14473 7000 -14447
rect 6730 -14607 7000 -14473
rect 6730 -14633 6855 -14607
rect 6881 -14633 7000 -14607
rect 6730 -14767 7000 -14633
rect 6730 -14793 6855 -14767
rect 6881 -14793 7000 -14767
rect 6730 -14927 7000 -14793
rect 6730 -14953 6855 -14927
rect 6881 -14953 7000 -14927
rect 6730 -15087 7000 -14953
rect 6730 -15113 6855 -15087
rect 6881 -15113 7000 -15087
rect 6730 -15230 7000 -15113
rect 3000 -15247 7000 -15230
rect 3000 -15273 3122 -15247
rect 3148 -15273 6855 -15247
rect 6881 -15273 7000 -15247
rect 3000 -15352 7000 -15273
rect 3000 -15378 3307 -15352
rect 3333 -15378 3467 -15352
rect 3493 -15378 3627 -15352
rect 3653 -15378 3787 -15352
rect 3813 -15378 3947 -15352
rect 3973 -15378 4107 -15352
rect 4133 -15378 4267 -15352
rect 4293 -15378 4427 -15352
rect 4453 -15378 4587 -15352
rect 4613 -15378 4747 -15352
rect 4773 -15378 4907 -15352
rect 4933 -15378 5067 -15352
rect 5093 -15378 5227 -15352
rect 5253 -15378 5387 -15352
rect 5413 -15378 5547 -15352
rect 5573 -15378 5707 -15352
rect 5733 -15378 5867 -15352
rect 5893 -15378 6027 -15352
rect 6053 -15378 6187 -15352
rect 6213 -15378 6347 -15352
rect 6373 -15378 6507 -15352
rect 6533 -15378 6667 -15352
rect 6693 -15378 7000 -15352
rect 3000 -15500 7000 -15378
rect 9000 -11624 13000 -11500
rect 9000 -11650 9307 -11624
rect 9333 -11650 9467 -11624
rect 9493 -11650 9627 -11624
rect 9653 -11650 9787 -11624
rect 9813 -11650 9947 -11624
rect 9973 -11650 10107 -11624
rect 10133 -11650 10267 -11624
rect 10293 -11650 10427 -11624
rect 10453 -11650 10587 -11624
rect 10613 -11650 10747 -11624
rect 10773 -11650 10907 -11624
rect 10933 -11650 11067 -11624
rect 11093 -11650 11227 -11624
rect 11253 -11650 11387 -11624
rect 11413 -11650 11547 -11624
rect 11573 -11650 11707 -11624
rect 11733 -11650 11867 -11624
rect 11893 -11650 12027 -11624
rect 12053 -11650 12187 -11624
rect 12213 -11650 12347 -11624
rect 12373 -11650 12507 -11624
rect 12533 -11650 12667 -11624
rect 12693 -11650 13000 -11624
rect 9000 -11727 13000 -11650
rect 9000 -11753 9122 -11727
rect 9148 -11753 12855 -11727
rect 12881 -11753 13000 -11727
rect 9000 -11770 13000 -11753
rect 9000 -11887 9270 -11770
rect 9000 -11913 9122 -11887
rect 9148 -11913 9270 -11887
rect 9000 -12047 9270 -11913
rect 9000 -12073 9122 -12047
rect 9148 -12073 9270 -12047
rect 9000 -12207 9270 -12073
rect 9000 -12233 9122 -12207
rect 9148 -12233 9270 -12207
rect 9000 -12367 9270 -12233
rect 9000 -12393 9122 -12367
rect 9148 -12393 9270 -12367
rect 9000 -12527 9270 -12393
rect 9000 -12553 9122 -12527
rect 9148 -12553 9270 -12527
rect 9000 -12687 9270 -12553
rect 9000 -12713 9122 -12687
rect 9148 -12713 9270 -12687
rect 9000 -12847 9270 -12713
rect 9000 -12873 9122 -12847
rect 9148 -12873 9270 -12847
rect 9000 -13007 9270 -12873
rect 9000 -13033 9122 -13007
rect 9148 -13033 9270 -13007
rect 9000 -13167 9270 -13033
rect 9000 -13193 9122 -13167
rect 9148 -13193 9270 -13167
rect 9000 -13327 9270 -13193
rect 9000 -13353 9122 -13327
rect 9148 -13353 9270 -13327
rect 9000 -13487 9270 -13353
rect 9000 -13513 9122 -13487
rect 9148 -13513 9270 -13487
rect 9000 -13647 9270 -13513
rect 9000 -13673 9122 -13647
rect 9148 -13673 9270 -13647
rect 9000 -13807 9270 -13673
rect 9000 -13833 9122 -13807
rect 9148 -13833 9270 -13807
rect 9000 -13967 9270 -13833
rect 9000 -13993 9122 -13967
rect 9148 -13993 9270 -13967
rect 9000 -14127 9270 -13993
rect 9000 -14153 9122 -14127
rect 9148 -14153 9270 -14127
rect 9000 -14287 9270 -14153
rect 9000 -14313 9122 -14287
rect 9148 -14313 9270 -14287
rect 9000 -14447 9270 -14313
rect 9000 -14473 9122 -14447
rect 9148 -14473 9270 -14447
rect 9000 -14607 9270 -14473
rect 9000 -14633 9122 -14607
rect 9148 -14633 9270 -14607
rect 9000 -14767 9270 -14633
rect 9000 -14793 9122 -14767
rect 9148 -14793 9270 -14767
rect 9000 -14927 9270 -14793
rect 9000 -14953 9122 -14927
rect 9148 -14953 9270 -14927
rect 9000 -15087 9270 -14953
rect 9000 -15113 9122 -15087
rect 9148 -15113 9270 -15087
rect 9000 -15230 9270 -15113
rect 12730 -11887 13000 -11770
rect 12730 -11913 12855 -11887
rect 12881 -11913 13000 -11887
rect 12730 -12047 13000 -11913
rect 12730 -12073 12855 -12047
rect 12881 -12073 13000 -12047
rect 12730 -12207 13000 -12073
rect 12730 -12233 12855 -12207
rect 12881 -12233 13000 -12207
rect 12730 -12367 13000 -12233
rect 12730 -12393 12855 -12367
rect 12881 -12393 13000 -12367
rect 12730 -12527 13000 -12393
rect 12730 -12553 12855 -12527
rect 12881 -12553 13000 -12527
rect 12730 -12687 13000 -12553
rect 12730 -12713 12855 -12687
rect 12881 -12713 13000 -12687
rect 12730 -12847 13000 -12713
rect 12730 -12873 12855 -12847
rect 12881 -12873 13000 -12847
rect 12730 -13007 13000 -12873
rect 12730 -13033 12855 -13007
rect 12881 -13033 13000 -13007
rect 12730 -13167 13000 -13033
rect 12730 -13193 12855 -13167
rect 12881 -13193 13000 -13167
rect 12730 -13327 13000 -13193
rect 12730 -13353 12855 -13327
rect 12881 -13353 13000 -13327
rect 12730 -13487 13000 -13353
rect 12730 -13513 12855 -13487
rect 12881 -13513 13000 -13487
rect 12730 -13647 13000 -13513
rect 12730 -13673 12855 -13647
rect 12881 -13673 13000 -13647
rect 12730 -13807 13000 -13673
rect 12730 -13833 12855 -13807
rect 12881 -13833 13000 -13807
rect 12730 -13967 13000 -13833
rect 12730 -13993 12855 -13967
rect 12881 -13993 13000 -13967
rect 12730 -14127 13000 -13993
rect 12730 -14153 12855 -14127
rect 12881 -14153 13000 -14127
rect 12730 -14287 13000 -14153
rect 12730 -14313 12855 -14287
rect 12881 -14313 13000 -14287
rect 12730 -14447 13000 -14313
rect 12730 -14473 12855 -14447
rect 12881 -14473 13000 -14447
rect 12730 -14607 13000 -14473
rect 12730 -14633 12855 -14607
rect 12881 -14633 13000 -14607
rect 12730 -14767 13000 -14633
rect 12730 -14793 12855 -14767
rect 12881 -14793 13000 -14767
rect 12730 -14927 13000 -14793
rect 12730 -14953 12855 -14927
rect 12881 -14953 13000 -14927
rect 12730 -15087 13000 -14953
rect 12730 -15113 12855 -15087
rect 12881 -15113 13000 -15087
rect 12730 -15230 13000 -15113
rect 9000 -15247 13000 -15230
rect 9000 -15273 9122 -15247
rect 9148 -15273 12855 -15247
rect 12881 -15273 13000 -15247
rect 9000 -15352 13000 -15273
rect 9000 -15378 9307 -15352
rect 9333 -15378 9467 -15352
rect 9493 -15378 9627 -15352
rect 9653 -15378 9787 -15352
rect 9813 -15378 9947 -15352
rect 9973 -15378 10107 -15352
rect 10133 -15378 10267 -15352
rect 10293 -15378 10427 -15352
rect 10453 -15378 10587 -15352
rect 10613 -15378 10747 -15352
rect 10773 -15378 10907 -15352
rect 10933 -15378 11067 -15352
rect 11093 -15378 11227 -15352
rect 11253 -15378 11387 -15352
rect 11413 -15378 11547 -15352
rect 11573 -15378 11707 -15352
rect 11733 -15378 11867 -15352
rect 11893 -15378 12027 -15352
rect 12053 -15378 12187 -15352
rect 12213 -15378 12347 -15352
rect 12373 -15378 12507 -15352
rect 12533 -15378 12667 -15352
rect 12693 -15378 13000 -15352
rect 9000 -15500 13000 -15378
rect 15000 -11624 19000 -11500
rect 15000 -11650 15307 -11624
rect 15333 -11650 15467 -11624
rect 15493 -11650 15627 -11624
rect 15653 -11650 15787 -11624
rect 15813 -11650 15947 -11624
rect 15973 -11650 16107 -11624
rect 16133 -11650 16267 -11624
rect 16293 -11650 16427 -11624
rect 16453 -11650 16587 -11624
rect 16613 -11650 16747 -11624
rect 16773 -11650 16907 -11624
rect 16933 -11650 17067 -11624
rect 17093 -11650 17227 -11624
rect 17253 -11650 17387 -11624
rect 17413 -11650 17547 -11624
rect 17573 -11650 17707 -11624
rect 17733 -11650 17867 -11624
rect 17893 -11650 18027 -11624
rect 18053 -11650 18187 -11624
rect 18213 -11650 18347 -11624
rect 18373 -11650 18507 -11624
rect 18533 -11650 18667 -11624
rect 18693 -11650 19000 -11624
rect 15000 -11727 19000 -11650
rect 15000 -11753 15122 -11727
rect 15148 -11753 18855 -11727
rect 18881 -11753 19000 -11727
rect 15000 -11770 19000 -11753
rect 15000 -11887 15270 -11770
rect 15000 -11913 15122 -11887
rect 15148 -11913 15270 -11887
rect 15000 -12047 15270 -11913
rect 15000 -12073 15122 -12047
rect 15148 -12073 15270 -12047
rect 15000 -12207 15270 -12073
rect 15000 -12233 15122 -12207
rect 15148 -12233 15270 -12207
rect 15000 -12367 15270 -12233
rect 15000 -12393 15122 -12367
rect 15148 -12393 15270 -12367
rect 15000 -12527 15270 -12393
rect 15000 -12553 15122 -12527
rect 15148 -12553 15270 -12527
rect 15000 -12687 15270 -12553
rect 15000 -12713 15122 -12687
rect 15148 -12713 15270 -12687
rect 15000 -12847 15270 -12713
rect 15000 -12873 15122 -12847
rect 15148 -12873 15270 -12847
rect 15000 -13007 15270 -12873
rect 15000 -13033 15122 -13007
rect 15148 -13033 15270 -13007
rect 15000 -13167 15270 -13033
rect 15000 -13193 15122 -13167
rect 15148 -13193 15270 -13167
rect 15000 -13327 15270 -13193
rect 15000 -13353 15122 -13327
rect 15148 -13353 15270 -13327
rect 15000 -13487 15270 -13353
rect 15000 -13513 15122 -13487
rect 15148 -13513 15270 -13487
rect 15000 -13647 15270 -13513
rect 15000 -13673 15122 -13647
rect 15148 -13673 15270 -13647
rect 15000 -13807 15270 -13673
rect 15000 -13833 15122 -13807
rect 15148 -13833 15270 -13807
rect 15000 -13967 15270 -13833
rect 15000 -13993 15122 -13967
rect 15148 -13993 15270 -13967
rect 15000 -14127 15270 -13993
rect 15000 -14153 15122 -14127
rect 15148 -14153 15270 -14127
rect 15000 -14287 15270 -14153
rect 15000 -14313 15122 -14287
rect 15148 -14313 15270 -14287
rect 15000 -14447 15270 -14313
rect 15000 -14473 15122 -14447
rect 15148 -14473 15270 -14447
rect 15000 -14607 15270 -14473
rect 15000 -14633 15122 -14607
rect 15148 -14633 15270 -14607
rect 15000 -14767 15270 -14633
rect 15000 -14793 15122 -14767
rect 15148 -14793 15270 -14767
rect 15000 -14927 15270 -14793
rect 15000 -14953 15122 -14927
rect 15148 -14953 15270 -14927
rect 15000 -15087 15270 -14953
rect 15000 -15113 15122 -15087
rect 15148 -15113 15270 -15087
rect 15000 -15230 15270 -15113
rect 18730 -11887 19000 -11770
rect 18730 -11913 18855 -11887
rect 18881 -11913 19000 -11887
rect 18730 -12047 19000 -11913
rect 18730 -12073 18855 -12047
rect 18881 -12073 19000 -12047
rect 18730 -12207 19000 -12073
rect 18730 -12233 18855 -12207
rect 18881 -12233 19000 -12207
rect 18730 -12367 19000 -12233
rect 18730 -12393 18855 -12367
rect 18881 -12393 19000 -12367
rect 18730 -12527 19000 -12393
rect 18730 -12553 18855 -12527
rect 18881 -12553 19000 -12527
rect 18730 -12687 19000 -12553
rect 18730 -12713 18855 -12687
rect 18881 -12713 19000 -12687
rect 18730 -12847 19000 -12713
rect 18730 -12873 18855 -12847
rect 18881 -12873 19000 -12847
rect 18730 -13007 19000 -12873
rect 18730 -13033 18855 -13007
rect 18881 -13033 19000 -13007
rect 18730 -13167 19000 -13033
rect 18730 -13193 18855 -13167
rect 18881 -13193 19000 -13167
rect 18730 -13327 19000 -13193
rect 18730 -13353 18855 -13327
rect 18881 -13353 19000 -13327
rect 18730 -13487 19000 -13353
rect 18730 -13513 18855 -13487
rect 18881 -13513 19000 -13487
rect 18730 -13647 19000 -13513
rect 18730 -13673 18855 -13647
rect 18881 -13673 19000 -13647
rect 18730 -13807 19000 -13673
rect 18730 -13833 18855 -13807
rect 18881 -13833 19000 -13807
rect 18730 -13967 19000 -13833
rect 18730 -13993 18855 -13967
rect 18881 -13993 19000 -13967
rect 18730 -14127 19000 -13993
rect 18730 -14153 18855 -14127
rect 18881 -14153 19000 -14127
rect 18730 -14287 19000 -14153
rect 18730 -14313 18855 -14287
rect 18881 -14313 19000 -14287
rect 18730 -14447 19000 -14313
rect 18730 -14473 18855 -14447
rect 18881 -14473 19000 -14447
rect 18730 -14607 19000 -14473
rect 18730 -14633 18855 -14607
rect 18881 -14633 19000 -14607
rect 18730 -14767 19000 -14633
rect 18730 -14793 18855 -14767
rect 18881 -14793 19000 -14767
rect 18730 -14927 19000 -14793
rect 18730 -14953 18855 -14927
rect 18881 -14953 19000 -14927
rect 18730 -15087 19000 -14953
rect 18730 -15113 18855 -15087
rect 18881 -15113 19000 -15087
rect 18730 -15230 19000 -15113
rect 15000 -15247 19000 -15230
rect 15000 -15273 15122 -15247
rect 15148 -15273 18855 -15247
rect 18881 -15273 19000 -15247
rect 15000 -15352 19000 -15273
rect 15000 -15378 15307 -15352
rect 15333 -15378 15467 -15352
rect 15493 -15378 15627 -15352
rect 15653 -15378 15787 -15352
rect 15813 -15378 15947 -15352
rect 15973 -15378 16107 -15352
rect 16133 -15378 16267 -15352
rect 16293 -15378 16427 -15352
rect 16453 -15378 16587 -15352
rect 16613 -15378 16747 -15352
rect 16773 -15378 16907 -15352
rect 16933 -15378 17067 -15352
rect 17093 -15378 17227 -15352
rect 17253 -15378 17387 -15352
rect 17413 -15378 17547 -15352
rect 17573 -15378 17707 -15352
rect 17733 -15378 17867 -15352
rect 17893 -15378 18027 -15352
rect 18053 -15378 18187 -15352
rect 18213 -15378 18347 -15352
rect 18373 -15378 18507 -15352
rect 18533 -15378 18667 -15352
rect 18693 -15378 19000 -15352
rect 15000 -15500 19000 -15378
rect 21000 -11624 25000 -11500
rect 21000 -11650 21307 -11624
rect 21333 -11650 21467 -11624
rect 21493 -11650 21627 -11624
rect 21653 -11650 21787 -11624
rect 21813 -11650 21947 -11624
rect 21973 -11650 22107 -11624
rect 22133 -11650 22267 -11624
rect 22293 -11650 22427 -11624
rect 22453 -11650 22587 -11624
rect 22613 -11650 22747 -11624
rect 22773 -11650 22907 -11624
rect 22933 -11650 23067 -11624
rect 23093 -11650 23227 -11624
rect 23253 -11650 23387 -11624
rect 23413 -11650 23547 -11624
rect 23573 -11650 23707 -11624
rect 23733 -11650 23867 -11624
rect 23893 -11650 24027 -11624
rect 24053 -11650 24187 -11624
rect 24213 -11650 24347 -11624
rect 24373 -11650 24507 -11624
rect 24533 -11650 24667 -11624
rect 24693 -11650 25000 -11624
rect 21000 -11727 25000 -11650
rect 21000 -11753 21122 -11727
rect 21148 -11753 24855 -11727
rect 24881 -11753 25000 -11727
rect 21000 -11770 25000 -11753
rect 21000 -11887 21270 -11770
rect 21000 -11913 21122 -11887
rect 21148 -11913 21270 -11887
rect 21000 -12047 21270 -11913
rect 21000 -12073 21122 -12047
rect 21148 -12073 21270 -12047
rect 21000 -12207 21270 -12073
rect 21000 -12233 21122 -12207
rect 21148 -12233 21270 -12207
rect 21000 -12367 21270 -12233
rect 21000 -12393 21122 -12367
rect 21148 -12393 21270 -12367
rect 21000 -12527 21270 -12393
rect 21000 -12553 21122 -12527
rect 21148 -12553 21270 -12527
rect 21000 -12687 21270 -12553
rect 21000 -12713 21122 -12687
rect 21148 -12713 21270 -12687
rect 21000 -12847 21270 -12713
rect 21000 -12873 21122 -12847
rect 21148 -12873 21270 -12847
rect 21000 -13007 21270 -12873
rect 21000 -13033 21122 -13007
rect 21148 -13033 21270 -13007
rect 21000 -13167 21270 -13033
rect 21000 -13193 21122 -13167
rect 21148 -13193 21270 -13167
rect 21000 -13327 21270 -13193
rect 21000 -13353 21122 -13327
rect 21148 -13353 21270 -13327
rect 21000 -13487 21270 -13353
rect 21000 -13513 21122 -13487
rect 21148 -13513 21270 -13487
rect 21000 -13647 21270 -13513
rect 21000 -13673 21122 -13647
rect 21148 -13673 21270 -13647
rect 21000 -13807 21270 -13673
rect 21000 -13833 21122 -13807
rect 21148 -13833 21270 -13807
rect 21000 -13967 21270 -13833
rect 21000 -13993 21122 -13967
rect 21148 -13993 21270 -13967
rect 21000 -14127 21270 -13993
rect 21000 -14153 21122 -14127
rect 21148 -14153 21270 -14127
rect 21000 -14287 21270 -14153
rect 21000 -14313 21122 -14287
rect 21148 -14313 21270 -14287
rect 21000 -14447 21270 -14313
rect 21000 -14473 21122 -14447
rect 21148 -14473 21270 -14447
rect 21000 -14607 21270 -14473
rect 21000 -14633 21122 -14607
rect 21148 -14633 21270 -14607
rect 21000 -14767 21270 -14633
rect 21000 -14793 21122 -14767
rect 21148 -14793 21270 -14767
rect 21000 -14927 21270 -14793
rect 21000 -14953 21122 -14927
rect 21148 -14953 21270 -14927
rect 21000 -15087 21270 -14953
rect 21000 -15113 21122 -15087
rect 21148 -15113 21270 -15087
rect 21000 -15230 21270 -15113
rect 24730 -11887 25000 -11770
rect 24730 -11913 24855 -11887
rect 24881 -11913 25000 -11887
rect 24730 -12047 25000 -11913
rect 24730 -12073 24855 -12047
rect 24881 -12073 25000 -12047
rect 24730 -12207 25000 -12073
rect 24730 -12233 24855 -12207
rect 24881 -12233 25000 -12207
rect 24730 -12367 25000 -12233
rect 24730 -12393 24855 -12367
rect 24881 -12393 25000 -12367
rect 24730 -12527 25000 -12393
rect 24730 -12553 24855 -12527
rect 24881 -12553 25000 -12527
rect 24730 -12687 25000 -12553
rect 24730 -12713 24855 -12687
rect 24881 -12713 25000 -12687
rect 24730 -12847 25000 -12713
rect 24730 -12873 24855 -12847
rect 24881 -12873 25000 -12847
rect 24730 -13007 25000 -12873
rect 24730 -13033 24855 -13007
rect 24881 -13033 25000 -13007
rect 24730 -13167 25000 -13033
rect 24730 -13193 24855 -13167
rect 24881 -13193 25000 -13167
rect 24730 -13327 25000 -13193
rect 24730 -13353 24855 -13327
rect 24881 -13353 25000 -13327
rect 24730 -13487 25000 -13353
rect 24730 -13513 24855 -13487
rect 24881 -13513 25000 -13487
rect 24730 -13647 25000 -13513
rect 24730 -13673 24855 -13647
rect 24881 -13673 25000 -13647
rect 24730 -13807 25000 -13673
rect 24730 -13833 24855 -13807
rect 24881 -13833 25000 -13807
rect 24730 -13967 25000 -13833
rect 24730 -13993 24855 -13967
rect 24881 -13993 25000 -13967
rect 24730 -14127 25000 -13993
rect 24730 -14153 24855 -14127
rect 24881 -14153 25000 -14127
rect 24730 -14287 25000 -14153
rect 24730 -14313 24855 -14287
rect 24881 -14313 25000 -14287
rect 24730 -14447 25000 -14313
rect 24730 -14473 24855 -14447
rect 24881 -14473 25000 -14447
rect 24730 -14607 25000 -14473
rect 24730 -14633 24855 -14607
rect 24881 -14633 25000 -14607
rect 24730 -14767 25000 -14633
rect 24730 -14793 24855 -14767
rect 24881 -14793 25000 -14767
rect 24730 -14927 25000 -14793
rect 24730 -14953 24855 -14927
rect 24881 -14953 25000 -14927
rect 24730 -15087 25000 -14953
rect 24730 -15113 24855 -15087
rect 24881 -15113 25000 -15087
rect 24730 -15230 25000 -15113
rect 21000 -15247 25000 -15230
rect 21000 -15273 21122 -15247
rect 21148 -15273 24855 -15247
rect 24881 -15273 25000 -15247
rect 21000 -15352 25000 -15273
rect 21000 -15378 21307 -15352
rect 21333 -15378 21467 -15352
rect 21493 -15378 21627 -15352
rect 21653 -15378 21787 -15352
rect 21813 -15378 21947 -15352
rect 21973 -15378 22107 -15352
rect 22133 -15378 22267 -15352
rect 22293 -15378 22427 -15352
rect 22453 -15378 22587 -15352
rect 22613 -15378 22747 -15352
rect 22773 -15378 22907 -15352
rect 22933 -15378 23067 -15352
rect 23093 -15378 23227 -15352
rect 23253 -15378 23387 -15352
rect 23413 -15378 23547 -15352
rect 23573 -15378 23707 -15352
rect 23733 -15378 23867 -15352
rect 23893 -15378 24027 -15352
rect 24053 -15378 24187 -15352
rect 24213 -15378 24347 -15352
rect 24373 -15378 24507 -15352
rect 24533 -15378 24667 -15352
rect 24693 -15378 25000 -15352
rect 21000 -15500 25000 -15378
<< via1 >>
rect 3307 9352 3333 9378
rect 3467 9352 3493 9378
rect 3627 9352 3653 9378
rect 3787 9352 3813 9378
rect 3947 9352 3973 9378
rect 4107 9352 4133 9378
rect 4267 9352 4293 9378
rect 4427 9352 4453 9378
rect 4587 9352 4613 9378
rect 4747 9352 4773 9378
rect 4907 9352 4933 9378
rect 5067 9352 5093 9378
rect 5227 9352 5253 9378
rect 5387 9352 5413 9378
rect 5547 9352 5573 9378
rect 5707 9352 5733 9378
rect 5867 9352 5893 9378
rect 6027 9352 6053 9378
rect 6187 9352 6213 9378
rect 6347 9352 6373 9378
rect 6507 9352 6533 9378
rect 6667 9352 6693 9378
rect 3119 9247 3145 9273
rect 6852 9247 6878 9273
rect 3119 9087 3145 9113
rect 3119 8927 3145 8953
rect 3119 8767 3145 8793
rect 3119 8607 3145 8633
rect 3119 8447 3145 8473
rect 3119 8287 3145 8313
rect 3119 8127 3145 8153
rect 3119 7967 3145 7993
rect 3119 7807 3145 7833
rect 3119 7647 3145 7673
rect 3119 7487 3145 7513
rect 3119 7327 3145 7353
rect 3119 7167 3145 7193
rect 3119 7007 3145 7033
rect 3119 6847 3145 6873
rect 3119 6687 3145 6713
rect 3119 6527 3145 6553
rect 3119 6367 3145 6393
rect 3119 6207 3145 6233
rect 3119 6047 3145 6073
rect 3119 5887 3145 5913
rect 6852 9087 6878 9113
rect 6852 8927 6878 8953
rect 6852 8767 6878 8793
rect 6852 8607 6878 8633
rect 6852 8447 6878 8473
rect 6852 8287 6878 8313
rect 6852 8127 6878 8153
rect 6852 7967 6878 7993
rect 6852 7807 6878 7833
rect 6852 7647 6878 7673
rect 6852 7487 6878 7513
rect 6852 7327 6878 7353
rect 6852 7167 6878 7193
rect 6852 7007 6878 7033
rect 6852 6847 6878 6873
rect 6852 6687 6878 6713
rect 6852 6527 6878 6553
rect 6852 6367 6878 6393
rect 6852 6207 6878 6233
rect 6852 6047 6878 6073
rect 6852 5887 6878 5913
rect 3119 5727 3145 5753
rect 6852 5727 6878 5753
rect 3307 5624 3333 5650
rect 3467 5624 3493 5650
rect 3627 5624 3653 5650
rect 3787 5624 3813 5650
rect 3947 5624 3973 5650
rect 4107 5624 4133 5650
rect 4267 5624 4293 5650
rect 4427 5624 4453 5650
rect 4587 5624 4613 5650
rect 4747 5624 4773 5650
rect 4907 5624 4933 5650
rect 5067 5624 5093 5650
rect 5227 5624 5253 5650
rect 5387 5624 5413 5650
rect 5547 5624 5573 5650
rect 5707 5624 5733 5650
rect 5867 5624 5893 5650
rect 6027 5624 6053 5650
rect 6187 5624 6213 5650
rect 6347 5624 6373 5650
rect 6507 5624 6533 5650
rect 6667 5624 6693 5650
rect 9307 9352 9333 9378
rect 9467 9352 9493 9378
rect 9627 9352 9653 9378
rect 9787 9352 9813 9378
rect 9947 9352 9973 9378
rect 10107 9352 10133 9378
rect 10267 9352 10293 9378
rect 10427 9352 10453 9378
rect 10587 9352 10613 9378
rect 10747 9352 10773 9378
rect 10907 9352 10933 9378
rect 11067 9352 11093 9378
rect 11227 9352 11253 9378
rect 11387 9352 11413 9378
rect 11547 9352 11573 9378
rect 11707 9352 11733 9378
rect 11867 9352 11893 9378
rect 12027 9352 12053 9378
rect 12187 9352 12213 9378
rect 12347 9352 12373 9378
rect 12507 9352 12533 9378
rect 12667 9352 12693 9378
rect 9119 9247 9145 9273
rect 12852 9247 12878 9273
rect 9119 9087 9145 9113
rect 9119 8927 9145 8953
rect 9119 8767 9145 8793
rect 9119 8607 9145 8633
rect 9119 8447 9145 8473
rect 9119 8287 9145 8313
rect 9119 8127 9145 8153
rect 9119 7967 9145 7993
rect 9119 7807 9145 7833
rect 9119 7647 9145 7673
rect 9119 7487 9145 7513
rect 9119 7327 9145 7353
rect 9119 7167 9145 7193
rect 9119 7007 9145 7033
rect 9119 6847 9145 6873
rect 9119 6687 9145 6713
rect 9119 6527 9145 6553
rect 9119 6367 9145 6393
rect 9119 6207 9145 6233
rect 9119 6047 9145 6073
rect 9119 5887 9145 5913
rect 12852 9087 12878 9113
rect 12852 8927 12878 8953
rect 12852 8767 12878 8793
rect 12852 8607 12878 8633
rect 12852 8447 12878 8473
rect 12852 8287 12878 8313
rect 12852 8127 12878 8153
rect 12852 7967 12878 7993
rect 12852 7807 12878 7833
rect 12852 7647 12878 7673
rect 12852 7487 12878 7513
rect 12852 7327 12878 7353
rect 12852 7167 12878 7193
rect 12852 7007 12878 7033
rect 12852 6847 12878 6873
rect 12852 6687 12878 6713
rect 12852 6527 12878 6553
rect 12852 6367 12878 6393
rect 12852 6207 12878 6233
rect 12852 6047 12878 6073
rect 12852 5887 12878 5913
rect 9119 5727 9145 5753
rect 12852 5727 12878 5753
rect 9307 5624 9333 5650
rect 9467 5624 9493 5650
rect 9627 5624 9653 5650
rect 9787 5624 9813 5650
rect 9947 5624 9973 5650
rect 10107 5624 10133 5650
rect 10267 5624 10293 5650
rect 10427 5624 10453 5650
rect 10587 5624 10613 5650
rect 10747 5624 10773 5650
rect 10907 5624 10933 5650
rect 11067 5624 11093 5650
rect 11227 5624 11253 5650
rect 11387 5624 11413 5650
rect 11547 5624 11573 5650
rect 11707 5624 11733 5650
rect 11867 5624 11893 5650
rect 12027 5624 12053 5650
rect 12187 5624 12213 5650
rect 12347 5624 12373 5650
rect 12507 5624 12533 5650
rect 12667 5624 12693 5650
rect 15307 9352 15333 9378
rect 15467 9352 15493 9378
rect 15627 9352 15653 9378
rect 15787 9352 15813 9378
rect 15947 9352 15973 9378
rect 16107 9352 16133 9378
rect 16267 9352 16293 9378
rect 16427 9352 16453 9378
rect 16587 9352 16613 9378
rect 16747 9352 16773 9378
rect 16907 9352 16933 9378
rect 17067 9352 17093 9378
rect 17227 9352 17253 9378
rect 17387 9352 17413 9378
rect 17547 9352 17573 9378
rect 17707 9352 17733 9378
rect 17867 9352 17893 9378
rect 18027 9352 18053 9378
rect 18187 9352 18213 9378
rect 18347 9352 18373 9378
rect 18507 9352 18533 9378
rect 18667 9352 18693 9378
rect 15119 9247 15145 9273
rect 18852 9247 18878 9273
rect 15119 9087 15145 9113
rect 15119 8927 15145 8953
rect 15119 8767 15145 8793
rect 15119 8607 15145 8633
rect 15119 8447 15145 8473
rect 15119 8287 15145 8313
rect 15119 8127 15145 8153
rect 15119 7967 15145 7993
rect 15119 7807 15145 7833
rect 15119 7647 15145 7673
rect 15119 7487 15145 7513
rect 15119 7327 15145 7353
rect 15119 7167 15145 7193
rect 15119 7007 15145 7033
rect 15119 6847 15145 6873
rect 15119 6687 15145 6713
rect 15119 6527 15145 6553
rect 15119 6367 15145 6393
rect 15119 6207 15145 6233
rect 15119 6047 15145 6073
rect 15119 5887 15145 5913
rect 18852 9087 18878 9113
rect 18852 8927 18878 8953
rect 18852 8767 18878 8793
rect 18852 8607 18878 8633
rect 18852 8447 18878 8473
rect 18852 8287 18878 8313
rect 18852 8127 18878 8153
rect 18852 7967 18878 7993
rect 18852 7807 18878 7833
rect 18852 7647 18878 7673
rect 18852 7487 18878 7513
rect 18852 7327 18878 7353
rect 18852 7167 18878 7193
rect 18852 7007 18878 7033
rect 18852 6847 18878 6873
rect 18852 6687 18878 6713
rect 18852 6527 18878 6553
rect 18852 6367 18878 6393
rect 18852 6207 18878 6233
rect 18852 6047 18878 6073
rect 18852 5887 18878 5913
rect 15119 5727 15145 5753
rect 18852 5727 18878 5753
rect 15307 5624 15333 5650
rect 15467 5624 15493 5650
rect 15627 5624 15653 5650
rect 15787 5624 15813 5650
rect 15947 5624 15973 5650
rect 16107 5624 16133 5650
rect 16267 5624 16293 5650
rect 16427 5624 16453 5650
rect 16587 5624 16613 5650
rect 16747 5624 16773 5650
rect 16907 5624 16933 5650
rect 17067 5624 17093 5650
rect 17227 5624 17253 5650
rect 17387 5624 17413 5650
rect 17547 5624 17573 5650
rect 17707 5624 17733 5650
rect 17867 5624 17893 5650
rect 18027 5624 18053 5650
rect 18187 5624 18213 5650
rect 18347 5624 18373 5650
rect 18507 5624 18533 5650
rect 18667 5624 18693 5650
rect 21307 9352 21333 9378
rect 21467 9352 21493 9378
rect 21627 9352 21653 9378
rect 21787 9352 21813 9378
rect 21947 9352 21973 9378
rect 22107 9352 22133 9378
rect 22267 9352 22293 9378
rect 22427 9352 22453 9378
rect 22587 9352 22613 9378
rect 22747 9352 22773 9378
rect 22907 9352 22933 9378
rect 23067 9352 23093 9378
rect 23227 9352 23253 9378
rect 23387 9352 23413 9378
rect 23547 9352 23573 9378
rect 23707 9352 23733 9378
rect 23867 9352 23893 9378
rect 24027 9352 24053 9378
rect 24187 9352 24213 9378
rect 24347 9352 24373 9378
rect 24507 9352 24533 9378
rect 24667 9352 24693 9378
rect 21119 9247 21145 9273
rect 24852 9247 24878 9273
rect 21119 9087 21145 9113
rect 21119 8927 21145 8953
rect 21119 8767 21145 8793
rect 21119 8607 21145 8633
rect 21119 8447 21145 8473
rect 21119 8287 21145 8313
rect 21119 8127 21145 8153
rect 21119 7967 21145 7993
rect 21119 7807 21145 7833
rect 21119 7647 21145 7673
rect 21119 7487 21145 7513
rect 21119 7327 21145 7353
rect 21119 7167 21145 7193
rect 21119 7007 21145 7033
rect 21119 6847 21145 6873
rect 21119 6687 21145 6713
rect 21119 6527 21145 6553
rect 21119 6367 21145 6393
rect 21119 6207 21145 6233
rect 21119 6047 21145 6073
rect 21119 5887 21145 5913
rect 24852 9087 24878 9113
rect 24852 8927 24878 8953
rect 24852 8767 24878 8793
rect 24852 8607 24878 8633
rect 24852 8447 24878 8473
rect 24852 8287 24878 8313
rect 24852 8127 24878 8153
rect 24852 7967 24878 7993
rect 24852 7807 24878 7833
rect 24852 7647 24878 7673
rect 24852 7487 24878 7513
rect 24852 7327 24878 7353
rect 24852 7167 24878 7193
rect 24852 7007 24878 7033
rect 24852 6847 24878 6873
rect 24852 6687 24878 6713
rect 24852 6527 24878 6553
rect 24852 6367 24878 6393
rect 24852 6207 24878 6233
rect 24852 6047 24878 6073
rect 24852 5887 24878 5913
rect 21119 5727 21145 5753
rect 24852 5727 24878 5753
rect 21307 5624 21333 5650
rect 21467 5624 21493 5650
rect 21627 5624 21653 5650
rect 21787 5624 21813 5650
rect 21947 5624 21973 5650
rect 22107 5624 22133 5650
rect 22267 5624 22293 5650
rect 22427 5624 22453 5650
rect 22587 5624 22613 5650
rect 22747 5624 22773 5650
rect 22907 5624 22933 5650
rect 23067 5624 23093 5650
rect 23227 5624 23253 5650
rect 23387 5624 23413 5650
rect 23547 5624 23573 5650
rect 23707 5624 23733 5650
rect 23867 5624 23893 5650
rect 24027 5624 24053 5650
rect 24187 5624 24213 5650
rect 24347 5624 24373 5650
rect 24507 5624 24533 5650
rect 24667 5624 24693 5650
rect 3307 3352 3333 3378
rect 3467 3352 3493 3378
rect 3627 3352 3653 3378
rect 3787 3352 3813 3378
rect 3947 3352 3973 3378
rect 4107 3352 4133 3378
rect 4267 3352 4293 3378
rect 4427 3352 4453 3378
rect 4587 3352 4613 3378
rect 4747 3352 4773 3378
rect 4907 3352 4933 3378
rect 5067 3352 5093 3378
rect 5227 3352 5253 3378
rect 5387 3352 5413 3378
rect 5547 3352 5573 3378
rect 5707 3352 5733 3378
rect 5867 3352 5893 3378
rect 6027 3352 6053 3378
rect 6187 3352 6213 3378
rect 6347 3352 6373 3378
rect 6507 3352 6533 3378
rect 6667 3352 6693 3378
rect 3119 3247 3145 3273
rect 6852 3247 6878 3273
rect 3119 3087 3145 3113
rect 3119 2927 3145 2953
rect 3119 2767 3145 2793
rect 3119 2607 3145 2633
rect 3119 2447 3145 2473
rect 3119 2287 3145 2313
rect 3119 2127 3145 2153
rect 3119 1967 3145 1993
rect 3119 1807 3145 1833
rect 3119 1647 3145 1673
rect 3119 1487 3145 1513
rect 3119 1327 3145 1353
rect 3119 1167 3145 1193
rect 3119 1007 3145 1033
rect 3119 847 3145 873
rect 3119 687 3145 713
rect 3119 527 3145 553
rect 3119 367 3145 393
rect 3119 207 3145 233
rect 3119 47 3145 73
rect 3119 -113 3145 -87
rect 6852 3087 6878 3113
rect 6852 2927 6878 2953
rect 6852 2767 6878 2793
rect 6852 2607 6878 2633
rect 6852 2447 6878 2473
rect 6852 2287 6878 2313
rect 6852 2127 6878 2153
rect 6852 1967 6878 1993
rect 6852 1807 6878 1833
rect 6852 1647 6878 1673
rect 6852 1487 6878 1513
rect 6852 1327 6878 1353
rect 6852 1167 6878 1193
rect 6852 1007 6878 1033
rect 6852 847 6878 873
rect 6852 687 6878 713
rect 6852 527 6878 553
rect 6852 367 6878 393
rect 6852 207 6878 233
rect 6852 47 6878 73
rect 6852 -113 6878 -87
rect 3119 -273 3145 -247
rect 6852 -273 6878 -247
rect 3307 -376 3333 -350
rect 3467 -376 3493 -350
rect 3627 -376 3653 -350
rect 3787 -376 3813 -350
rect 3947 -376 3973 -350
rect 4107 -376 4133 -350
rect 4267 -376 4293 -350
rect 4427 -376 4453 -350
rect 4587 -376 4613 -350
rect 4747 -376 4773 -350
rect 4907 -376 4933 -350
rect 5067 -376 5093 -350
rect 5227 -376 5253 -350
rect 5387 -376 5413 -350
rect 5547 -376 5573 -350
rect 5707 -376 5733 -350
rect 5867 -376 5893 -350
rect 6027 -376 6053 -350
rect 6187 -376 6213 -350
rect 6347 -376 6373 -350
rect 6507 -376 6533 -350
rect 6667 -376 6693 -350
rect 9307 3352 9333 3378
rect 9467 3352 9493 3378
rect 9627 3352 9653 3378
rect 9787 3352 9813 3378
rect 9947 3352 9973 3378
rect 10107 3352 10133 3378
rect 10267 3352 10293 3378
rect 10427 3352 10453 3378
rect 10587 3352 10613 3378
rect 10747 3352 10773 3378
rect 10907 3352 10933 3378
rect 11067 3352 11093 3378
rect 11227 3352 11253 3378
rect 11387 3352 11413 3378
rect 11547 3352 11573 3378
rect 11707 3352 11733 3378
rect 11867 3352 11893 3378
rect 12027 3352 12053 3378
rect 12187 3352 12213 3378
rect 12347 3352 12373 3378
rect 12507 3352 12533 3378
rect 12667 3352 12693 3378
rect 9119 3247 9145 3273
rect 12852 3247 12878 3273
rect 9119 3087 9145 3113
rect 9119 2927 9145 2953
rect 9119 2767 9145 2793
rect 9119 2607 9145 2633
rect 9119 2447 9145 2473
rect 9119 2287 9145 2313
rect 9119 2127 9145 2153
rect 9119 1967 9145 1993
rect 9119 1807 9145 1833
rect 9119 1647 9145 1673
rect 9119 1487 9145 1513
rect 9119 1327 9145 1353
rect 9119 1167 9145 1193
rect 9119 1007 9145 1033
rect 9119 847 9145 873
rect 9119 687 9145 713
rect 9119 527 9145 553
rect 9119 367 9145 393
rect 9119 207 9145 233
rect 9119 47 9145 73
rect 9119 -113 9145 -87
rect 12852 3087 12878 3113
rect 12852 2927 12878 2953
rect 12852 2767 12878 2793
rect 12852 2607 12878 2633
rect 12852 2447 12878 2473
rect 12852 2287 12878 2313
rect 12852 2127 12878 2153
rect 12852 1967 12878 1993
rect 12852 1807 12878 1833
rect 12852 1647 12878 1673
rect 12852 1487 12878 1513
rect 12852 1327 12878 1353
rect 12852 1167 12878 1193
rect 12852 1007 12878 1033
rect 12852 847 12878 873
rect 12852 687 12878 713
rect 12852 527 12878 553
rect 12852 367 12878 393
rect 12852 207 12878 233
rect 12852 47 12878 73
rect 12852 -113 12878 -87
rect 9119 -273 9145 -247
rect 12852 -273 12878 -247
rect 9307 -376 9333 -350
rect 9467 -376 9493 -350
rect 9627 -376 9653 -350
rect 9787 -376 9813 -350
rect 9947 -376 9973 -350
rect 10107 -376 10133 -350
rect 10267 -376 10293 -350
rect 10427 -376 10453 -350
rect 10587 -376 10613 -350
rect 10747 -376 10773 -350
rect 10907 -376 10933 -350
rect 11067 -376 11093 -350
rect 11227 -376 11253 -350
rect 11387 -376 11413 -350
rect 11547 -376 11573 -350
rect 11707 -376 11733 -350
rect 11867 -376 11893 -350
rect 12027 -376 12053 -350
rect 12187 -376 12213 -350
rect 12347 -376 12373 -350
rect 12507 -376 12533 -350
rect 12667 -376 12693 -350
rect 15307 3352 15333 3378
rect 15467 3352 15493 3378
rect 15627 3352 15653 3378
rect 15787 3352 15813 3378
rect 15947 3352 15973 3378
rect 16107 3352 16133 3378
rect 16267 3352 16293 3378
rect 16427 3352 16453 3378
rect 16587 3352 16613 3378
rect 16747 3352 16773 3378
rect 16907 3352 16933 3378
rect 17067 3352 17093 3378
rect 17227 3352 17253 3378
rect 17387 3352 17413 3378
rect 17547 3352 17573 3378
rect 17707 3352 17733 3378
rect 17867 3352 17893 3378
rect 18027 3352 18053 3378
rect 18187 3352 18213 3378
rect 18347 3352 18373 3378
rect 18507 3352 18533 3378
rect 18667 3352 18693 3378
rect 15119 3247 15145 3273
rect 18852 3247 18878 3273
rect 15119 3087 15145 3113
rect 15119 2927 15145 2953
rect 15119 2767 15145 2793
rect 15119 2607 15145 2633
rect 15119 2447 15145 2473
rect 15119 2287 15145 2313
rect 15119 2127 15145 2153
rect 15119 1967 15145 1993
rect 15119 1807 15145 1833
rect 15119 1647 15145 1673
rect 15119 1487 15145 1513
rect 15119 1327 15145 1353
rect 15119 1167 15145 1193
rect 15119 1007 15145 1033
rect 15119 847 15145 873
rect 15119 687 15145 713
rect 15119 527 15145 553
rect 15119 367 15145 393
rect 15119 207 15145 233
rect 15119 47 15145 73
rect 15119 -113 15145 -87
rect 18852 3087 18878 3113
rect 18852 2927 18878 2953
rect 18852 2767 18878 2793
rect 18852 2607 18878 2633
rect 18852 2447 18878 2473
rect 18852 2287 18878 2313
rect 18852 2127 18878 2153
rect 18852 1967 18878 1993
rect 18852 1807 18878 1833
rect 18852 1647 18878 1673
rect 18852 1487 18878 1513
rect 18852 1327 18878 1353
rect 18852 1167 18878 1193
rect 18852 1007 18878 1033
rect 18852 847 18878 873
rect 18852 687 18878 713
rect 18852 527 18878 553
rect 18852 367 18878 393
rect 18852 207 18878 233
rect 18852 47 18878 73
rect 18852 -113 18878 -87
rect 15119 -273 15145 -247
rect 18852 -273 18878 -247
rect 15307 -376 15333 -350
rect 15467 -376 15493 -350
rect 15627 -376 15653 -350
rect 15787 -376 15813 -350
rect 15947 -376 15973 -350
rect 16107 -376 16133 -350
rect 16267 -376 16293 -350
rect 16427 -376 16453 -350
rect 16587 -376 16613 -350
rect 16747 -376 16773 -350
rect 16907 -376 16933 -350
rect 17067 -376 17093 -350
rect 17227 -376 17253 -350
rect 17387 -376 17413 -350
rect 17547 -376 17573 -350
rect 17707 -376 17733 -350
rect 17867 -376 17893 -350
rect 18027 -376 18053 -350
rect 18187 -376 18213 -350
rect 18347 -376 18373 -350
rect 18507 -376 18533 -350
rect 18667 -376 18693 -350
rect 21307 3352 21333 3378
rect 21467 3352 21493 3378
rect 21627 3352 21653 3378
rect 21787 3352 21813 3378
rect 21947 3352 21973 3378
rect 22107 3352 22133 3378
rect 22267 3352 22293 3378
rect 22427 3352 22453 3378
rect 22587 3352 22613 3378
rect 22747 3352 22773 3378
rect 22907 3352 22933 3378
rect 23067 3352 23093 3378
rect 23227 3352 23253 3378
rect 23387 3352 23413 3378
rect 23547 3352 23573 3378
rect 23707 3352 23733 3378
rect 23867 3352 23893 3378
rect 24027 3352 24053 3378
rect 24187 3352 24213 3378
rect 24347 3352 24373 3378
rect 24507 3352 24533 3378
rect 24667 3352 24693 3378
rect 21119 3247 21145 3273
rect 24852 3247 24878 3273
rect 21119 3087 21145 3113
rect 21119 2927 21145 2953
rect 21119 2767 21145 2793
rect 21119 2607 21145 2633
rect 21119 2447 21145 2473
rect 21119 2287 21145 2313
rect 21119 2127 21145 2153
rect 21119 1967 21145 1993
rect 21119 1807 21145 1833
rect 21119 1647 21145 1673
rect 21119 1487 21145 1513
rect 21119 1327 21145 1353
rect 21119 1167 21145 1193
rect 21119 1007 21145 1033
rect 21119 847 21145 873
rect 21119 687 21145 713
rect 21119 527 21145 553
rect 21119 367 21145 393
rect 21119 207 21145 233
rect 21119 47 21145 73
rect 21119 -113 21145 -87
rect 24852 3087 24878 3113
rect 24852 2927 24878 2953
rect 24852 2767 24878 2793
rect 24852 2607 24878 2633
rect 24852 2447 24878 2473
rect 24852 2287 24878 2313
rect 24852 2127 24878 2153
rect 24852 1967 24878 1993
rect 24852 1807 24878 1833
rect 24852 1647 24878 1673
rect 24852 1487 24878 1513
rect 24852 1327 24878 1353
rect 24852 1167 24878 1193
rect 24852 1007 24878 1033
rect 24852 847 24878 873
rect 24852 687 24878 713
rect 24852 527 24878 553
rect 24852 367 24878 393
rect 24852 207 24878 233
rect 24852 47 24878 73
rect 24852 -113 24878 -87
rect 21119 -273 21145 -247
rect 24852 -273 24878 -247
rect 21307 -376 21333 -350
rect 21467 -376 21493 -350
rect 21627 -376 21653 -350
rect 21787 -376 21813 -350
rect 21947 -376 21973 -350
rect 22107 -376 22133 -350
rect 22267 -376 22293 -350
rect 22427 -376 22453 -350
rect 22587 -376 22613 -350
rect 22747 -376 22773 -350
rect 22907 -376 22933 -350
rect 23067 -376 23093 -350
rect 23227 -376 23253 -350
rect 23387 -376 23413 -350
rect 23547 -376 23573 -350
rect 23707 -376 23733 -350
rect 23867 -376 23893 -350
rect 24027 -376 24053 -350
rect 24187 -376 24213 -350
rect 24347 -376 24373 -350
rect 24507 -376 24533 -350
rect 24667 -376 24693 -350
rect 19245 -745 19290 -575
rect 19435 -690 19485 -630
rect 19600 -745 19645 -575
rect 20035 -1170 20065 -1140
rect 20070 -1240 20100 -1210
rect 16250 -2050 16350 -1950
rect 16155 -2180 16225 -2140
rect 16295 -2180 16365 -2140
rect 16250 -2400 16350 -2300
rect 11650 -3700 11750 -3600
rect 11635 -3860 11705 -3820
rect 11775 -3860 11845 -3820
rect 11650 -4050 11750 -3950
rect 8200 -4790 8230 -4760
rect 8235 -4860 8265 -4830
rect 8355 -5425 8400 -5255
rect 8515 -5370 8565 -5310
rect 8710 -5425 8755 -5255
rect 3307 -5650 3333 -5624
rect 3467 -5650 3493 -5624
rect 3627 -5650 3653 -5624
rect 3787 -5650 3813 -5624
rect 3947 -5650 3973 -5624
rect 4107 -5650 4133 -5624
rect 4267 -5650 4293 -5624
rect 4427 -5650 4453 -5624
rect 4587 -5650 4613 -5624
rect 4747 -5650 4773 -5624
rect 4907 -5650 4933 -5624
rect 5067 -5650 5093 -5624
rect 5227 -5650 5253 -5624
rect 5387 -5650 5413 -5624
rect 5547 -5650 5573 -5624
rect 5707 -5650 5733 -5624
rect 5867 -5650 5893 -5624
rect 6027 -5650 6053 -5624
rect 6187 -5650 6213 -5624
rect 6347 -5650 6373 -5624
rect 6507 -5650 6533 -5624
rect 6667 -5650 6693 -5624
rect 3122 -5753 3148 -5727
rect 6855 -5753 6881 -5727
rect 3122 -5913 3148 -5887
rect 3122 -6073 3148 -6047
rect 3122 -6233 3148 -6207
rect 3122 -6393 3148 -6367
rect 3122 -6553 3148 -6527
rect 3122 -6713 3148 -6687
rect 3122 -6873 3148 -6847
rect 3122 -7033 3148 -7007
rect 3122 -7193 3148 -7167
rect 3122 -7353 3148 -7327
rect 3122 -7513 3148 -7487
rect 3122 -7673 3148 -7647
rect 3122 -7833 3148 -7807
rect 3122 -7993 3148 -7967
rect 3122 -8153 3148 -8127
rect 3122 -8313 3148 -8287
rect 3122 -8473 3148 -8447
rect 3122 -8633 3148 -8607
rect 3122 -8793 3148 -8767
rect 3122 -8953 3148 -8927
rect 3122 -9113 3148 -9087
rect 6855 -5913 6881 -5887
rect 6855 -6073 6881 -6047
rect 6855 -6233 6881 -6207
rect 6855 -6393 6881 -6367
rect 6855 -6553 6881 -6527
rect 6855 -6713 6881 -6687
rect 6855 -6873 6881 -6847
rect 6855 -7033 6881 -7007
rect 6855 -7193 6881 -7167
rect 6855 -7353 6881 -7327
rect 6855 -7513 6881 -7487
rect 6855 -7673 6881 -7647
rect 6855 -7833 6881 -7807
rect 6855 -7993 6881 -7967
rect 6855 -8153 6881 -8127
rect 6855 -8313 6881 -8287
rect 6855 -8473 6881 -8447
rect 6855 -8633 6881 -8607
rect 6855 -8793 6881 -8767
rect 6855 -8953 6881 -8927
rect 6855 -9113 6881 -9087
rect 3122 -9273 3148 -9247
rect 6855 -9273 6881 -9247
rect 3307 -9378 3333 -9352
rect 3467 -9378 3493 -9352
rect 3627 -9378 3653 -9352
rect 3787 -9378 3813 -9352
rect 3947 -9378 3973 -9352
rect 4107 -9378 4133 -9352
rect 4267 -9378 4293 -9352
rect 4427 -9378 4453 -9352
rect 4587 -9378 4613 -9352
rect 4747 -9378 4773 -9352
rect 4907 -9378 4933 -9352
rect 5067 -9378 5093 -9352
rect 5227 -9378 5253 -9352
rect 5387 -9378 5413 -9352
rect 5547 -9378 5573 -9352
rect 5707 -9378 5733 -9352
rect 5867 -9378 5893 -9352
rect 6027 -9378 6053 -9352
rect 6187 -9378 6213 -9352
rect 6347 -9378 6373 -9352
rect 6507 -9378 6533 -9352
rect 6667 -9378 6693 -9352
rect 9307 -5650 9333 -5624
rect 9467 -5650 9493 -5624
rect 9627 -5650 9653 -5624
rect 9787 -5650 9813 -5624
rect 9947 -5650 9973 -5624
rect 10107 -5650 10133 -5624
rect 10267 -5650 10293 -5624
rect 10427 -5650 10453 -5624
rect 10587 -5650 10613 -5624
rect 10747 -5650 10773 -5624
rect 10907 -5650 10933 -5624
rect 11067 -5650 11093 -5624
rect 11227 -5650 11253 -5624
rect 11387 -5650 11413 -5624
rect 11547 -5650 11573 -5624
rect 11707 -5650 11733 -5624
rect 11867 -5650 11893 -5624
rect 12027 -5650 12053 -5624
rect 12187 -5650 12213 -5624
rect 12347 -5650 12373 -5624
rect 12507 -5650 12533 -5624
rect 12667 -5650 12693 -5624
rect 9122 -5753 9148 -5727
rect 12855 -5753 12881 -5727
rect 9122 -5913 9148 -5887
rect 9122 -6073 9148 -6047
rect 9122 -6233 9148 -6207
rect 9122 -6393 9148 -6367
rect 9122 -6553 9148 -6527
rect 9122 -6713 9148 -6687
rect 9122 -6873 9148 -6847
rect 9122 -7033 9148 -7007
rect 9122 -7193 9148 -7167
rect 9122 -7353 9148 -7327
rect 9122 -7513 9148 -7487
rect 9122 -7673 9148 -7647
rect 9122 -7833 9148 -7807
rect 9122 -7993 9148 -7967
rect 9122 -8153 9148 -8127
rect 9122 -8313 9148 -8287
rect 9122 -8473 9148 -8447
rect 9122 -8633 9148 -8607
rect 9122 -8793 9148 -8767
rect 9122 -8953 9148 -8927
rect 9122 -9113 9148 -9087
rect 12855 -5913 12881 -5887
rect 12855 -6073 12881 -6047
rect 12855 -6233 12881 -6207
rect 12855 -6393 12881 -6367
rect 12855 -6553 12881 -6527
rect 12855 -6713 12881 -6687
rect 12855 -6873 12881 -6847
rect 12855 -7033 12881 -7007
rect 12855 -7193 12881 -7167
rect 12855 -7353 12881 -7327
rect 12855 -7513 12881 -7487
rect 12855 -7673 12881 -7647
rect 12855 -7833 12881 -7807
rect 12855 -7993 12881 -7967
rect 12855 -8153 12881 -8127
rect 12855 -8313 12881 -8287
rect 12855 -8473 12881 -8447
rect 12855 -8633 12881 -8607
rect 12855 -8793 12881 -8767
rect 12855 -8953 12881 -8927
rect 12855 -9113 12881 -9087
rect 9122 -9273 9148 -9247
rect 12855 -9273 12881 -9247
rect 9307 -9378 9333 -9352
rect 9467 -9378 9493 -9352
rect 9627 -9378 9653 -9352
rect 9787 -9378 9813 -9352
rect 9947 -9378 9973 -9352
rect 10107 -9378 10133 -9352
rect 10267 -9378 10293 -9352
rect 10427 -9378 10453 -9352
rect 10587 -9378 10613 -9352
rect 10747 -9378 10773 -9352
rect 10907 -9378 10933 -9352
rect 11067 -9378 11093 -9352
rect 11227 -9378 11253 -9352
rect 11387 -9378 11413 -9352
rect 11547 -9378 11573 -9352
rect 11707 -9378 11733 -9352
rect 11867 -9378 11893 -9352
rect 12027 -9378 12053 -9352
rect 12187 -9378 12213 -9352
rect 12347 -9378 12373 -9352
rect 12507 -9378 12533 -9352
rect 12667 -9378 12693 -9352
rect 15307 -5650 15333 -5624
rect 15467 -5650 15493 -5624
rect 15627 -5650 15653 -5624
rect 15787 -5650 15813 -5624
rect 15947 -5650 15973 -5624
rect 16107 -5650 16133 -5624
rect 16267 -5650 16293 -5624
rect 16427 -5650 16453 -5624
rect 16587 -5650 16613 -5624
rect 16747 -5650 16773 -5624
rect 16907 -5650 16933 -5624
rect 17067 -5650 17093 -5624
rect 17227 -5650 17253 -5624
rect 17387 -5650 17413 -5624
rect 17547 -5650 17573 -5624
rect 17707 -5650 17733 -5624
rect 17867 -5650 17893 -5624
rect 18027 -5650 18053 -5624
rect 18187 -5650 18213 -5624
rect 18347 -5650 18373 -5624
rect 18507 -5650 18533 -5624
rect 18667 -5650 18693 -5624
rect 15122 -5753 15148 -5727
rect 18855 -5753 18881 -5727
rect 15122 -5913 15148 -5887
rect 15122 -6073 15148 -6047
rect 15122 -6233 15148 -6207
rect 15122 -6393 15148 -6367
rect 15122 -6553 15148 -6527
rect 15122 -6713 15148 -6687
rect 15122 -6873 15148 -6847
rect 15122 -7033 15148 -7007
rect 15122 -7193 15148 -7167
rect 15122 -7353 15148 -7327
rect 15122 -7513 15148 -7487
rect 15122 -7673 15148 -7647
rect 15122 -7833 15148 -7807
rect 15122 -7993 15148 -7967
rect 15122 -8153 15148 -8127
rect 15122 -8313 15148 -8287
rect 15122 -8473 15148 -8447
rect 15122 -8633 15148 -8607
rect 15122 -8793 15148 -8767
rect 15122 -8953 15148 -8927
rect 15122 -9113 15148 -9087
rect 18855 -5913 18881 -5887
rect 18855 -6073 18881 -6047
rect 18855 -6233 18881 -6207
rect 18855 -6393 18881 -6367
rect 18855 -6553 18881 -6527
rect 18855 -6713 18881 -6687
rect 18855 -6873 18881 -6847
rect 18855 -7033 18881 -7007
rect 18855 -7193 18881 -7167
rect 18855 -7353 18881 -7327
rect 18855 -7513 18881 -7487
rect 18855 -7673 18881 -7647
rect 18855 -7833 18881 -7807
rect 18855 -7993 18881 -7967
rect 18855 -8153 18881 -8127
rect 18855 -8313 18881 -8287
rect 18855 -8473 18881 -8447
rect 18855 -8633 18881 -8607
rect 18855 -8793 18881 -8767
rect 18855 -8953 18881 -8927
rect 18855 -9113 18881 -9087
rect 15122 -9273 15148 -9247
rect 18855 -9273 18881 -9247
rect 15307 -9378 15333 -9352
rect 15467 -9378 15493 -9352
rect 15627 -9378 15653 -9352
rect 15787 -9378 15813 -9352
rect 15947 -9378 15973 -9352
rect 16107 -9378 16133 -9352
rect 16267 -9378 16293 -9352
rect 16427 -9378 16453 -9352
rect 16587 -9378 16613 -9352
rect 16747 -9378 16773 -9352
rect 16907 -9378 16933 -9352
rect 17067 -9378 17093 -9352
rect 17227 -9378 17253 -9352
rect 17387 -9378 17413 -9352
rect 17547 -9378 17573 -9352
rect 17707 -9378 17733 -9352
rect 17867 -9378 17893 -9352
rect 18027 -9378 18053 -9352
rect 18187 -9378 18213 -9352
rect 18347 -9378 18373 -9352
rect 18507 -9378 18533 -9352
rect 18667 -9378 18693 -9352
rect 21307 -5650 21333 -5624
rect 21467 -5650 21493 -5624
rect 21627 -5650 21653 -5624
rect 21787 -5650 21813 -5624
rect 21947 -5650 21973 -5624
rect 22107 -5650 22133 -5624
rect 22267 -5650 22293 -5624
rect 22427 -5650 22453 -5624
rect 22587 -5650 22613 -5624
rect 22747 -5650 22773 -5624
rect 22907 -5650 22933 -5624
rect 23067 -5650 23093 -5624
rect 23227 -5650 23253 -5624
rect 23387 -5650 23413 -5624
rect 23547 -5650 23573 -5624
rect 23707 -5650 23733 -5624
rect 23867 -5650 23893 -5624
rect 24027 -5650 24053 -5624
rect 24187 -5650 24213 -5624
rect 24347 -5650 24373 -5624
rect 24507 -5650 24533 -5624
rect 24667 -5650 24693 -5624
rect 21122 -5753 21148 -5727
rect 24855 -5753 24881 -5727
rect 21122 -5913 21148 -5887
rect 21122 -6073 21148 -6047
rect 21122 -6233 21148 -6207
rect 21122 -6393 21148 -6367
rect 21122 -6553 21148 -6527
rect 21122 -6713 21148 -6687
rect 21122 -6873 21148 -6847
rect 21122 -7033 21148 -7007
rect 21122 -7193 21148 -7167
rect 21122 -7353 21148 -7327
rect 21122 -7513 21148 -7487
rect 21122 -7673 21148 -7647
rect 21122 -7833 21148 -7807
rect 21122 -7993 21148 -7967
rect 21122 -8153 21148 -8127
rect 21122 -8313 21148 -8287
rect 21122 -8473 21148 -8447
rect 21122 -8633 21148 -8607
rect 21122 -8793 21148 -8767
rect 21122 -8953 21148 -8927
rect 21122 -9113 21148 -9087
rect 24855 -5913 24881 -5887
rect 24855 -6073 24881 -6047
rect 24855 -6233 24881 -6207
rect 24855 -6393 24881 -6367
rect 24855 -6553 24881 -6527
rect 24855 -6713 24881 -6687
rect 24855 -6873 24881 -6847
rect 24855 -7033 24881 -7007
rect 24855 -7193 24881 -7167
rect 24855 -7353 24881 -7327
rect 24855 -7513 24881 -7487
rect 24855 -7673 24881 -7647
rect 24855 -7833 24881 -7807
rect 24855 -7993 24881 -7967
rect 24855 -8153 24881 -8127
rect 24855 -8313 24881 -8287
rect 24855 -8473 24881 -8447
rect 24855 -8633 24881 -8607
rect 24855 -8793 24881 -8767
rect 24855 -8953 24881 -8927
rect 24855 -9113 24881 -9087
rect 21122 -9273 21148 -9247
rect 24855 -9273 24881 -9247
rect 21307 -9378 21333 -9352
rect 21467 -9378 21493 -9352
rect 21627 -9378 21653 -9352
rect 21787 -9378 21813 -9352
rect 21947 -9378 21973 -9352
rect 22107 -9378 22133 -9352
rect 22267 -9378 22293 -9352
rect 22427 -9378 22453 -9352
rect 22587 -9378 22613 -9352
rect 22747 -9378 22773 -9352
rect 22907 -9378 22933 -9352
rect 23067 -9378 23093 -9352
rect 23227 -9378 23253 -9352
rect 23387 -9378 23413 -9352
rect 23547 -9378 23573 -9352
rect 23707 -9378 23733 -9352
rect 23867 -9378 23893 -9352
rect 24027 -9378 24053 -9352
rect 24187 -9378 24213 -9352
rect 24347 -9378 24373 -9352
rect 24507 -9378 24533 -9352
rect 24667 -9378 24693 -9352
rect 3307 -11650 3333 -11624
rect 3467 -11650 3493 -11624
rect 3627 -11650 3653 -11624
rect 3787 -11650 3813 -11624
rect 3947 -11650 3973 -11624
rect 4107 -11650 4133 -11624
rect 4267 -11650 4293 -11624
rect 4427 -11650 4453 -11624
rect 4587 -11650 4613 -11624
rect 4747 -11650 4773 -11624
rect 4907 -11650 4933 -11624
rect 5067 -11650 5093 -11624
rect 5227 -11650 5253 -11624
rect 5387 -11650 5413 -11624
rect 5547 -11650 5573 -11624
rect 5707 -11650 5733 -11624
rect 5867 -11650 5893 -11624
rect 6027 -11650 6053 -11624
rect 6187 -11650 6213 -11624
rect 6347 -11650 6373 -11624
rect 6507 -11650 6533 -11624
rect 6667 -11650 6693 -11624
rect 3122 -11753 3148 -11727
rect 6855 -11753 6881 -11727
rect 3122 -11913 3148 -11887
rect 3122 -12073 3148 -12047
rect 3122 -12233 3148 -12207
rect 3122 -12393 3148 -12367
rect 3122 -12553 3148 -12527
rect 3122 -12713 3148 -12687
rect 3122 -12873 3148 -12847
rect 3122 -13033 3148 -13007
rect 3122 -13193 3148 -13167
rect 3122 -13353 3148 -13327
rect 3122 -13513 3148 -13487
rect 3122 -13673 3148 -13647
rect 3122 -13833 3148 -13807
rect 3122 -13993 3148 -13967
rect 3122 -14153 3148 -14127
rect 3122 -14313 3148 -14287
rect 3122 -14473 3148 -14447
rect 3122 -14633 3148 -14607
rect 3122 -14793 3148 -14767
rect 3122 -14953 3148 -14927
rect 3122 -15113 3148 -15087
rect 6855 -11913 6881 -11887
rect 6855 -12073 6881 -12047
rect 6855 -12233 6881 -12207
rect 6855 -12393 6881 -12367
rect 6855 -12553 6881 -12527
rect 6855 -12713 6881 -12687
rect 6855 -12873 6881 -12847
rect 6855 -13033 6881 -13007
rect 6855 -13193 6881 -13167
rect 6855 -13353 6881 -13327
rect 6855 -13513 6881 -13487
rect 6855 -13673 6881 -13647
rect 6855 -13833 6881 -13807
rect 6855 -13993 6881 -13967
rect 6855 -14153 6881 -14127
rect 6855 -14313 6881 -14287
rect 6855 -14473 6881 -14447
rect 6855 -14633 6881 -14607
rect 6855 -14793 6881 -14767
rect 6855 -14953 6881 -14927
rect 6855 -15113 6881 -15087
rect 3122 -15273 3148 -15247
rect 6855 -15273 6881 -15247
rect 3307 -15378 3333 -15352
rect 3467 -15378 3493 -15352
rect 3627 -15378 3653 -15352
rect 3787 -15378 3813 -15352
rect 3947 -15378 3973 -15352
rect 4107 -15378 4133 -15352
rect 4267 -15378 4293 -15352
rect 4427 -15378 4453 -15352
rect 4587 -15378 4613 -15352
rect 4747 -15378 4773 -15352
rect 4907 -15378 4933 -15352
rect 5067 -15378 5093 -15352
rect 5227 -15378 5253 -15352
rect 5387 -15378 5413 -15352
rect 5547 -15378 5573 -15352
rect 5707 -15378 5733 -15352
rect 5867 -15378 5893 -15352
rect 6027 -15378 6053 -15352
rect 6187 -15378 6213 -15352
rect 6347 -15378 6373 -15352
rect 6507 -15378 6533 -15352
rect 6667 -15378 6693 -15352
rect 9307 -11650 9333 -11624
rect 9467 -11650 9493 -11624
rect 9627 -11650 9653 -11624
rect 9787 -11650 9813 -11624
rect 9947 -11650 9973 -11624
rect 10107 -11650 10133 -11624
rect 10267 -11650 10293 -11624
rect 10427 -11650 10453 -11624
rect 10587 -11650 10613 -11624
rect 10747 -11650 10773 -11624
rect 10907 -11650 10933 -11624
rect 11067 -11650 11093 -11624
rect 11227 -11650 11253 -11624
rect 11387 -11650 11413 -11624
rect 11547 -11650 11573 -11624
rect 11707 -11650 11733 -11624
rect 11867 -11650 11893 -11624
rect 12027 -11650 12053 -11624
rect 12187 -11650 12213 -11624
rect 12347 -11650 12373 -11624
rect 12507 -11650 12533 -11624
rect 12667 -11650 12693 -11624
rect 9122 -11753 9148 -11727
rect 12855 -11753 12881 -11727
rect 9122 -11913 9148 -11887
rect 9122 -12073 9148 -12047
rect 9122 -12233 9148 -12207
rect 9122 -12393 9148 -12367
rect 9122 -12553 9148 -12527
rect 9122 -12713 9148 -12687
rect 9122 -12873 9148 -12847
rect 9122 -13033 9148 -13007
rect 9122 -13193 9148 -13167
rect 9122 -13353 9148 -13327
rect 9122 -13513 9148 -13487
rect 9122 -13673 9148 -13647
rect 9122 -13833 9148 -13807
rect 9122 -13993 9148 -13967
rect 9122 -14153 9148 -14127
rect 9122 -14313 9148 -14287
rect 9122 -14473 9148 -14447
rect 9122 -14633 9148 -14607
rect 9122 -14793 9148 -14767
rect 9122 -14953 9148 -14927
rect 9122 -15113 9148 -15087
rect 12855 -11913 12881 -11887
rect 12855 -12073 12881 -12047
rect 12855 -12233 12881 -12207
rect 12855 -12393 12881 -12367
rect 12855 -12553 12881 -12527
rect 12855 -12713 12881 -12687
rect 12855 -12873 12881 -12847
rect 12855 -13033 12881 -13007
rect 12855 -13193 12881 -13167
rect 12855 -13353 12881 -13327
rect 12855 -13513 12881 -13487
rect 12855 -13673 12881 -13647
rect 12855 -13833 12881 -13807
rect 12855 -13993 12881 -13967
rect 12855 -14153 12881 -14127
rect 12855 -14313 12881 -14287
rect 12855 -14473 12881 -14447
rect 12855 -14633 12881 -14607
rect 12855 -14793 12881 -14767
rect 12855 -14953 12881 -14927
rect 12855 -15113 12881 -15087
rect 9122 -15273 9148 -15247
rect 12855 -15273 12881 -15247
rect 9307 -15378 9333 -15352
rect 9467 -15378 9493 -15352
rect 9627 -15378 9653 -15352
rect 9787 -15378 9813 -15352
rect 9947 -15378 9973 -15352
rect 10107 -15378 10133 -15352
rect 10267 -15378 10293 -15352
rect 10427 -15378 10453 -15352
rect 10587 -15378 10613 -15352
rect 10747 -15378 10773 -15352
rect 10907 -15378 10933 -15352
rect 11067 -15378 11093 -15352
rect 11227 -15378 11253 -15352
rect 11387 -15378 11413 -15352
rect 11547 -15378 11573 -15352
rect 11707 -15378 11733 -15352
rect 11867 -15378 11893 -15352
rect 12027 -15378 12053 -15352
rect 12187 -15378 12213 -15352
rect 12347 -15378 12373 -15352
rect 12507 -15378 12533 -15352
rect 12667 -15378 12693 -15352
rect 15307 -11650 15333 -11624
rect 15467 -11650 15493 -11624
rect 15627 -11650 15653 -11624
rect 15787 -11650 15813 -11624
rect 15947 -11650 15973 -11624
rect 16107 -11650 16133 -11624
rect 16267 -11650 16293 -11624
rect 16427 -11650 16453 -11624
rect 16587 -11650 16613 -11624
rect 16747 -11650 16773 -11624
rect 16907 -11650 16933 -11624
rect 17067 -11650 17093 -11624
rect 17227 -11650 17253 -11624
rect 17387 -11650 17413 -11624
rect 17547 -11650 17573 -11624
rect 17707 -11650 17733 -11624
rect 17867 -11650 17893 -11624
rect 18027 -11650 18053 -11624
rect 18187 -11650 18213 -11624
rect 18347 -11650 18373 -11624
rect 18507 -11650 18533 -11624
rect 18667 -11650 18693 -11624
rect 15122 -11753 15148 -11727
rect 18855 -11753 18881 -11727
rect 15122 -11913 15148 -11887
rect 15122 -12073 15148 -12047
rect 15122 -12233 15148 -12207
rect 15122 -12393 15148 -12367
rect 15122 -12553 15148 -12527
rect 15122 -12713 15148 -12687
rect 15122 -12873 15148 -12847
rect 15122 -13033 15148 -13007
rect 15122 -13193 15148 -13167
rect 15122 -13353 15148 -13327
rect 15122 -13513 15148 -13487
rect 15122 -13673 15148 -13647
rect 15122 -13833 15148 -13807
rect 15122 -13993 15148 -13967
rect 15122 -14153 15148 -14127
rect 15122 -14313 15148 -14287
rect 15122 -14473 15148 -14447
rect 15122 -14633 15148 -14607
rect 15122 -14793 15148 -14767
rect 15122 -14953 15148 -14927
rect 15122 -15113 15148 -15087
rect 18855 -11913 18881 -11887
rect 18855 -12073 18881 -12047
rect 18855 -12233 18881 -12207
rect 18855 -12393 18881 -12367
rect 18855 -12553 18881 -12527
rect 18855 -12713 18881 -12687
rect 18855 -12873 18881 -12847
rect 18855 -13033 18881 -13007
rect 18855 -13193 18881 -13167
rect 18855 -13353 18881 -13327
rect 18855 -13513 18881 -13487
rect 18855 -13673 18881 -13647
rect 18855 -13833 18881 -13807
rect 18855 -13993 18881 -13967
rect 18855 -14153 18881 -14127
rect 18855 -14313 18881 -14287
rect 18855 -14473 18881 -14447
rect 18855 -14633 18881 -14607
rect 18855 -14793 18881 -14767
rect 18855 -14953 18881 -14927
rect 18855 -15113 18881 -15087
rect 15122 -15273 15148 -15247
rect 18855 -15273 18881 -15247
rect 15307 -15378 15333 -15352
rect 15467 -15378 15493 -15352
rect 15627 -15378 15653 -15352
rect 15787 -15378 15813 -15352
rect 15947 -15378 15973 -15352
rect 16107 -15378 16133 -15352
rect 16267 -15378 16293 -15352
rect 16427 -15378 16453 -15352
rect 16587 -15378 16613 -15352
rect 16747 -15378 16773 -15352
rect 16907 -15378 16933 -15352
rect 17067 -15378 17093 -15352
rect 17227 -15378 17253 -15352
rect 17387 -15378 17413 -15352
rect 17547 -15378 17573 -15352
rect 17707 -15378 17733 -15352
rect 17867 -15378 17893 -15352
rect 18027 -15378 18053 -15352
rect 18187 -15378 18213 -15352
rect 18347 -15378 18373 -15352
rect 18507 -15378 18533 -15352
rect 18667 -15378 18693 -15352
rect 21307 -11650 21333 -11624
rect 21467 -11650 21493 -11624
rect 21627 -11650 21653 -11624
rect 21787 -11650 21813 -11624
rect 21947 -11650 21973 -11624
rect 22107 -11650 22133 -11624
rect 22267 -11650 22293 -11624
rect 22427 -11650 22453 -11624
rect 22587 -11650 22613 -11624
rect 22747 -11650 22773 -11624
rect 22907 -11650 22933 -11624
rect 23067 -11650 23093 -11624
rect 23227 -11650 23253 -11624
rect 23387 -11650 23413 -11624
rect 23547 -11650 23573 -11624
rect 23707 -11650 23733 -11624
rect 23867 -11650 23893 -11624
rect 24027 -11650 24053 -11624
rect 24187 -11650 24213 -11624
rect 24347 -11650 24373 -11624
rect 24507 -11650 24533 -11624
rect 24667 -11650 24693 -11624
rect 21122 -11753 21148 -11727
rect 24855 -11753 24881 -11727
rect 21122 -11913 21148 -11887
rect 21122 -12073 21148 -12047
rect 21122 -12233 21148 -12207
rect 21122 -12393 21148 -12367
rect 21122 -12553 21148 -12527
rect 21122 -12713 21148 -12687
rect 21122 -12873 21148 -12847
rect 21122 -13033 21148 -13007
rect 21122 -13193 21148 -13167
rect 21122 -13353 21148 -13327
rect 21122 -13513 21148 -13487
rect 21122 -13673 21148 -13647
rect 21122 -13833 21148 -13807
rect 21122 -13993 21148 -13967
rect 21122 -14153 21148 -14127
rect 21122 -14313 21148 -14287
rect 21122 -14473 21148 -14447
rect 21122 -14633 21148 -14607
rect 21122 -14793 21148 -14767
rect 21122 -14953 21148 -14927
rect 21122 -15113 21148 -15087
rect 24855 -11913 24881 -11887
rect 24855 -12073 24881 -12047
rect 24855 -12233 24881 -12207
rect 24855 -12393 24881 -12367
rect 24855 -12553 24881 -12527
rect 24855 -12713 24881 -12687
rect 24855 -12873 24881 -12847
rect 24855 -13033 24881 -13007
rect 24855 -13193 24881 -13167
rect 24855 -13353 24881 -13327
rect 24855 -13513 24881 -13487
rect 24855 -13673 24881 -13647
rect 24855 -13833 24881 -13807
rect 24855 -13993 24881 -13967
rect 24855 -14153 24881 -14127
rect 24855 -14313 24881 -14287
rect 24855 -14473 24881 -14447
rect 24855 -14633 24881 -14607
rect 24855 -14793 24881 -14767
rect 24855 -14953 24881 -14927
rect 24855 -15113 24881 -15087
rect 21122 -15273 21148 -15247
rect 24855 -15273 24881 -15247
rect 21307 -15378 21333 -15352
rect 21467 -15378 21493 -15352
rect 21627 -15378 21653 -15352
rect 21787 -15378 21813 -15352
rect 21947 -15378 21973 -15352
rect 22107 -15378 22133 -15352
rect 22267 -15378 22293 -15352
rect 22427 -15378 22453 -15352
rect 22587 -15378 22613 -15352
rect 22747 -15378 22773 -15352
rect 22907 -15378 22933 -15352
rect 23067 -15378 23093 -15352
rect 23227 -15378 23253 -15352
rect 23387 -15378 23413 -15352
rect 23547 -15378 23573 -15352
rect 23707 -15378 23733 -15352
rect 23867 -15378 23893 -15352
rect 24027 -15378 24053 -15352
rect 24187 -15378 24213 -15352
rect 24347 -15378 24373 -15352
rect 24507 -15378 24533 -15352
rect 24667 -15378 24693 -15352
<< metal2 >>
rect 3000 9379 7000 9500
rect 3000 9351 3306 9379
rect 3334 9351 3466 9379
rect 3494 9351 3626 9379
rect 3654 9351 3786 9379
rect 3814 9351 3946 9379
rect 3974 9351 4106 9379
rect 4134 9351 4266 9379
rect 4294 9351 4426 9379
rect 4454 9351 4586 9379
rect 4614 9351 4746 9379
rect 4774 9351 4906 9379
rect 4934 9351 5066 9379
rect 5094 9351 5226 9379
rect 5254 9351 5386 9379
rect 5414 9351 5546 9379
rect 5574 9351 5706 9379
rect 5734 9351 5866 9379
rect 5894 9351 6026 9379
rect 6054 9351 6186 9379
rect 6214 9351 6346 9379
rect 6374 9351 6506 9379
rect 6534 9351 6666 9379
rect 6694 9351 7000 9379
rect 3000 9274 7000 9351
rect 3000 9246 3118 9274
rect 3146 9246 6851 9274
rect 6879 9246 7000 9274
rect 3000 9230 7000 9246
rect 3000 9114 3270 9230
rect 3000 9086 3118 9114
rect 3146 9086 3270 9114
rect 3000 8954 3270 9086
rect 3000 8926 3118 8954
rect 3146 8926 3270 8954
rect 3000 8794 3270 8926
rect 3000 8766 3118 8794
rect 3146 8766 3270 8794
rect 3000 8634 3270 8766
rect 3000 8606 3118 8634
rect 3146 8606 3270 8634
rect 3000 8474 3270 8606
rect 3000 8446 3118 8474
rect 3146 8446 3270 8474
rect 3000 8314 3270 8446
rect 3000 8286 3118 8314
rect 3146 8286 3270 8314
rect 3000 8154 3270 8286
rect 3000 8126 3118 8154
rect 3146 8126 3270 8154
rect 3000 7994 3270 8126
rect 3000 7966 3118 7994
rect 3146 7966 3270 7994
rect 3000 7834 3270 7966
rect 3000 7806 3118 7834
rect 3146 7806 3270 7834
rect 3000 7674 3270 7806
rect 3000 7646 3118 7674
rect 3146 7646 3270 7674
rect 3000 7514 3270 7646
rect 3000 7486 3118 7514
rect 3146 7486 3270 7514
rect 3000 7354 3270 7486
rect 3000 7326 3118 7354
rect 3146 7326 3270 7354
rect 3000 7194 3270 7326
rect 3000 7166 3118 7194
rect 3146 7166 3270 7194
rect 3000 7034 3270 7166
rect 3000 7006 3118 7034
rect 3146 7006 3270 7034
rect 3000 6874 3270 7006
rect 3000 6846 3118 6874
rect 3146 6846 3270 6874
rect 3000 6714 3270 6846
rect 3000 6686 3118 6714
rect 3146 6686 3270 6714
rect 3000 6554 3270 6686
rect 3000 6526 3118 6554
rect 3146 6526 3270 6554
rect 3000 6394 3270 6526
rect 3000 6366 3118 6394
rect 3146 6366 3270 6394
rect 3000 6234 3270 6366
rect 3000 6206 3118 6234
rect 3146 6206 3270 6234
rect 3000 6074 3270 6206
rect 3000 6046 3118 6074
rect 3146 6046 3270 6074
rect 3000 5914 3270 6046
rect 3000 5886 3118 5914
rect 3146 5886 3270 5914
rect 3000 5770 3270 5886
rect 6730 9114 7000 9230
rect 6730 9086 6851 9114
rect 6879 9086 7000 9114
rect 6730 8954 7000 9086
rect 6730 8926 6851 8954
rect 6879 8926 7000 8954
rect 6730 8794 7000 8926
rect 6730 8766 6851 8794
rect 6879 8766 7000 8794
rect 6730 8634 7000 8766
rect 6730 8606 6851 8634
rect 6879 8606 7000 8634
rect 6730 8474 7000 8606
rect 6730 8446 6851 8474
rect 6879 8446 7000 8474
rect 6730 8314 7000 8446
rect 6730 8286 6851 8314
rect 6879 8286 7000 8314
rect 6730 8154 7000 8286
rect 6730 8126 6851 8154
rect 6879 8126 7000 8154
rect 6730 7994 7000 8126
rect 6730 7966 6851 7994
rect 6879 7966 7000 7994
rect 6730 7834 7000 7966
rect 6730 7806 6851 7834
rect 6879 7806 7000 7834
rect 6730 7674 7000 7806
rect 6730 7646 6851 7674
rect 6879 7646 7000 7674
rect 6730 7514 7000 7646
rect 6730 7486 6851 7514
rect 6879 7486 7000 7514
rect 6730 7354 7000 7486
rect 6730 7326 6851 7354
rect 6879 7326 7000 7354
rect 6730 7194 7000 7326
rect 6730 7166 6851 7194
rect 6879 7166 7000 7194
rect 6730 7034 7000 7166
rect 6730 7006 6851 7034
rect 6879 7006 7000 7034
rect 6730 6874 7000 7006
rect 6730 6846 6851 6874
rect 6879 6846 7000 6874
rect 6730 6714 7000 6846
rect 6730 6686 6851 6714
rect 6879 6686 7000 6714
rect 6730 6554 7000 6686
rect 6730 6526 6851 6554
rect 6879 6526 7000 6554
rect 6730 6394 7000 6526
rect 6730 6366 6851 6394
rect 6879 6366 7000 6394
rect 6730 6234 7000 6366
rect 6730 6206 6851 6234
rect 6879 6206 7000 6234
rect 6730 6074 7000 6206
rect 6730 6046 6851 6074
rect 6879 6046 7000 6074
rect 6730 5914 7000 6046
rect 6730 5886 6851 5914
rect 6879 5886 7000 5914
rect 6730 5770 7000 5886
rect 3000 5754 7000 5770
rect 3000 5726 3118 5754
rect 3146 5726 6851 5754
rect 6879 5726 7000 5754
rect 3000 5651 7000 5726
rect 3000 5623 3306 5651
rect 3334 5623 3466 5651
rect 3494 5623 3626 5651
rect 3654 5623 3786 5651
rect 3814 5623 3946 5651
rect 3974 5623 4106 5651
rect 4134 5623 4266 5651
rect 4294 5623 4426 5651
rect 4454 5623 4586 5651
rect 4614 5623 4746 5651
rect 4774 5623 4906 5651
rect 4934 5623 5066 5651
rect 5094 5623 5226 5651
rect 5254 5623 5386 5651
rect 5414 5623 5546 5651
rect 5574 5623 5706 5651
rect 5734 5623 5866 5651
rect 5894 5623 6026 5651
rect 6054 5623 6186 5651
rect 6214 5623 6346 5651
rect 6374 5623 6506 5651
rect 6534 5623 6666 5651
rect 6694 5623 7000 5651
rect 3000 5500 7000 5623
rect 9000 9379 13000 9500
rect 9000 9351 9306 9379
rect 9334 9351 9466 9379
rect 9494 9351 9626 9379
rect 9654 9351 9786 9379
rect 9814 9351 9946 9379
rect 9974 9351 10106 9379
rect 10134 9351 10266 9379
rect 10294 9351 10426 9379
rect 10454 9351 10586 9379
rect 10614 9351 10746 9379
rect 10774 9351 10906 9379
rect 10934 9351 11066 9379
rect 11094 9351 11226 9379
rect 11254 9351 11386 9379
rect 11414 9351 11546 9379
rect 11574 9351 11706 9379
rect 11734 9351 11866 9379
rect 11894 9351 12026 9379
rect 12054 9351 12186 9379
rect 12214 9351 12346 9379
rect 12374 9351 12506 9379
rect 12534 9351 12666 9379
rect 12694 9351 13000 9379
rect 9000 9274 13000 9351
rect 9000 9246 9118 9274
rect 9146 9246 12851 9274
rect 12879 9246 13000 9274
rect 9000 9230 13000 9246
rect 9000 9114 9270 9230
rect 9000 9086 9118 9114
rect 9146 9086 9270 9114
rect 9000 8954 9270 9086
rect 9000 8926 9118 8954
rect 9146 8926 9270 8954
rect 9000 8794 9270 8926
rect 9000 8766 9118 8794
rect 9146 8766 9270 8794
rect 9000 8634 9270 8766
rect 9000 8606 9118 8634
rect 9146 8606 9270 8634
rect 9000 8474 9270 8606
rect 9000 8446 9118 8474
rect 9146 8446 9270 8474
rect 9000 8314 9270 8446
rect 9000 8286 9118 8314
rect 9146 8286 9270 8314
rect 9000 8154 9270 8286
rect 9000 8126 9118 8154
rect 9146 8126 9270 8154
rect 9000 7994 9270 8126
rect 9000 7966 9118 7994
rect 9146 7966 9270 7994
rect 9000 7834 9270 7966
rect 9000 7806 9118 7834
rect 9146 7806 9270 7834
rect 9000 7674 9270 7806
rect 9000 7646 9118 7674
rect 9146 7646 9270 7674
rect 9000 7514 9270 7646
rect 9000 7486 9118 7514
rect 9146 7486 9270 7514
rect 9000 7354 9270 7486
rect 9000 7326 9118 7354
rect 9146 7326 9270 7354
rect 9000 7194 9270 7326
rect 9000 7166 9118 7194
rect 9146 7166 9270 7194
rect 9000 7034 9270 7166
rect 9000 7006 9118 7034
rect 9146 7006 9270 7034
rect 9000 6874 9270 7006
rect 9000 6846 9118 6874
rect 9146 6846 9270 6874
rect 9000 6714 9270 6846
rect 9000 6686 9118 6714
rect 9146 6686 9270 6714
rect 9000 6554 9270 6686
rect 9000 6526 9118 6554
rect 9146 6526 9270 6554
rect 9000 6394 9270 6526
rect 9000 6366 9118 6394
rect 9146 6366 9270 6394
rect 9000 6234 9270 6366
rect 9000 6206 9118 6234
rect 9146 6206 9270 6234
rect 9000 6074 9270 6206
rect 9000 6046 9118 6074
rect 9146 6046 9270 6074
rect 9000 5914 9270 6046
rect 9000 5886 9118 5914
rect 9146 5886 9270 5914
rect 9000 5770 9270 5886
rect 12730 9114 13000 9230
rect 12730 9086 12851 9114
rect 12879 9086 13000 9114
rect 12730 8954 13000 9086
rect 12730 8926 12851 8954
rect 12879 8926 13000 8954
rect 12730 8794 13000 8926
rect 12730 8766 12851 8794
rect 12879 8766 13000 8794
rect 12730 8634 13000 8766
rect 12730 8606 12851 8634
rect 12879 8606 13000 8634
rect 12730 8474 13000 8606
rect 12730 8446 12851 8474
rect 12879 8446 13000 8474
rect 12730 8314 13000 8446
rect 12730 8286 12851 8314
rect 12879 8286 13000 8314
rect 12730 8154 13000 8286
rect 12730 8126 12851 8154
rect 12879 8126 13000 8154
rect 12730 7994 13000 8126
rect 12730 7966 12851 7994
rect 12879 7966 13000 7994
rect 12730 7834 13000 7966
rect 12730 7806 12851 7834
rect 12879 7806 13000 7834
rect 12730 7674 13000 7806
rect 12730 7646 12851 7674
rect 12879 7646 13000 7674
rect 12730 7514 13000 7646
rect 12730 7486 12851 7514
rect 12879 7486 13000 7514
rect 12730 7354 13000 7486
rect 12730 7326 12851 7354
rect 12879 7326 13000 7354
rect 12730 7194 13000 7326
rect 12730 7166 12851 7194
rect 12879 7166 13000 7194
rect 12730 7034 13000 7166
rect 12730 7006 12851 7034
rect 12879 7006 13000 7034
rect 12730 6874 13000 7006
rect 12730 6846 12851 6874
rect 12879 6846 13000 6874
rect 12730 6714 13000 6846
rect 12730 6686 12851 6714
rect 12879 6686 13000 6714
rect 12730 6554 13000 6686
rect 12730 6526 12851 6554
rect 12879 6526 13000 6554
rect 12730 6394 13000 6526
rect 12730 6366 12851 6394
rect 12879 6366 13000 6394
rect 12730 6234 13000 6366
rect 12730 6206 12851 6234
rect 12879 6206 13000 6234
rect 12730 6074 13000 6206
rect 12730 6046 12851 6074
rect 12879 6046 13000 6074
rect 12730 5914 13000 6046
rect 12730 5886 12851 5914
rect 12879 5886 13000 5914
rect 12730 5770 13000 5886
rect 9000 5754 13000 5770
rect 9000 5726 9118 5754
rect 9146 5726 12851 5754
rect 12879 5726 13000 5754
rect 9000 5651 13000 5726
rect 9000 5623 9306 5651
rect 9334 5623 9466 5651
rect 9494 5623 9626 5651
rect 9654 5623 9786 5651
rect 9814 5623 9946 5651
rect 9974 5623 10106 5651
rect 10134 5623 10266 5651
rect 10294 5623 10426 5651
rect 10454 5623 10586 5651
rect 10614 5623 10746 5651
rect 10774 5623 10906 5651
rect 10934 5623 11066 5651
rect 11094 5623 11226 5651
rect 11254 5623 11386 5651
rect 11414 5623 11546 5651
rect 11574 5623 11706 5651
rect 11734 5623 11866 5651
rect 11894 5623 12026 5651
rect 12054 5623 12186 5651
rect 12214 5623 12346 5651
rect 12374 5623 12506 5651
rect 12534 5623 12666 5651
rect 12694 5623 13000 5651
rect 9000 5500 13000 5623
rect 15000 9379 19000 9500
rect 15000 9351 15306 9379
rect 15334 9351 15466 9379
rect 15494 9351 15626 9379
rect 15654 9351 15786 9379
rect 15814 9351 15946 9379
rect 15974 9351 16106 9379
rect 16134 9351 16266 9379
rect 16294 9351 16426 9379
rect 16454 9351 16586 9379
rect 16614 9351 16746 9379
rect 16774 9351 16906 9379
rect 16934 9351 17066 9379
rect 17094 9351 17226 9379
rect 17254 9351 17386 9379
rect 17414 9351 17546 9379
rect 17574 9351 17706 9379
rect 17734 9351 17866 9379
rect 17894 9351 18026 9379
rect 18054 9351 18186 9379
rect 18214 9351 18346 9379
rect 18374 9351 18506 9379
rect 18534 9351 18666 9379
rect 18694 9351 19000 9379
rect 15000 9274 19000 9351
rect 15000 9246 15118 9274
rect 15146 9246 18851 9274
rect 18879 9246 19000 9274
rect 15000 9230 19000 9246
rect 15000 9114 15270 9230
rect 15000 9086 15118 9114
rect 15146 9086 15270 9114
rect 15000 8954 15270 9086
rect 15000 8926 15118 8954
rect 15146 8926 15270 8954
rect 15000 8794 15270 8926
rect 15000 8766 15118 8794
rect 15146 8766 15270 8794
rect 15000 8634 15270 8766
rect 15000 8606 15118 8634
rect 15146 8606 15270 8634
rect 15000 8474 15270 8606
rect 15000 8446 15118 8474
rect 15146 8446 15270 8474
rect 15000 8314 15270 8446
rect 15000 8286 15118 8314
rect 15146 8286 15270 8314
rect 15000 8154 15270 8286
rect 15000 8126 15118 8154
rect 15146 8126 15270 8154
rect 15000 7994 15270 8126
rect 15000 7966 15118 7994
rect 15146 7966 15270 7994
rect 15000 7834 15270 7966
rect 15000 7806 15118 7834
rect 15146 7806 15270 7834
rect 15000 7674 15270 7806
rect 15000 7646 15118 7674
rect 15146 7646 15270 7674
rect 15000 7514 15270 7646
rect 15000 7486 15118 7514
rect 15146 7486 15270 7514
rect 15000 7354 15270 7486
rect 15000 7326 15118 7354
rect 15146 7326 15270 7354
rect 15000 7194 15270 7326
rect 15000 7166 15118 7194
rect 15146 7166 15270 7194
rect 15000 7034 15270 7166
rect 15000 7006 15118 7034
rect 15146 7006 15270 7034
rect 15000 6874 15270 7006
rect 15000 6846 15118 6874
rect 15146 6846 15270 6874
rect 15000 6714 15270 6846
rect 15000 6686 15118 6714
rect 15146 6686 15270 6714
rect 15000 6554 15270 6686
rect 15000 6526 15118 6554
rect 15146 6526 15270 6554
rect 15000 6394 15270 6526
rect 15000 6366 15118 6394
rect 15146 6366 15270 6394
rect 15000 6234 15270 6366
rect 15000 6206 15118 6234
rect 15146 6206 15270 6234
rect 15000 6074 15270 6206
rect 15000 6046 15118 6074
rect 15146 6046 15270 6074
rect 15000 5914 15270 6046
rect 15000 5886 15118 5914
rect 15146 5886 15270 5914
rect 15000 5770 15270 5886
rect 18730 9114 19000 9230
rect 18730 9086 18851 9114
rect 18879 9086 19000 9114
rect 18730 8954 19000 9086
rect 18730 8926 18851 8954
rect 18879 8926 19000 8954
rect 18730 8794 19000 8926
rect 18730 8766 18851 8794
rect 18879 8766 19000 8794
rect 18730 8634 19000 8766
rect 18730 8606 18851 8634
rect 18879 8606 19000 8634
rect 18730 8474 19000 8606
rect 18730 8446 18851 8474
rect 18879 8446 19000 8474
rect 18730 8314 19000 8446
rect 18730 8286 18851 8314
rect 18879 8286 19000 8314
rect 18730 8154 19000 8286
rect 18730 8126 18851 8154
rect 18879 8126 19000 8154
rect 18730 7994 19000 8126
rect 18730 7966 18851 7994
rect 18879 7966 19000 7994
rect 18730 7834 19000 7966
rect 18730 7806 18851 7834
rect 18879 7806 19000 7834
rect 18730 7674 19000 7806
rect 18730 7646 18851 7674
rect 18879 7646 19000 7674
rect 18730 7514 19000 7646
rect 18730 7486 18851 7514
rect 18879 7486 19000 7514
rect 18730 7354 19000 7486
rect 18730 7326 18851 7354
rect 18879 7326 19000 7354
rect 18730 7194 19000 7326
rect 18730 7166 18851 7194
rect 18879 7166 19000 7194
rect 18730 7034 19000 7166
rect 18730 7006 18851 7034
rect 18879 7006 19000 7034
rect 18730 6874 19000 7006
rect 18730 6846 18851 6874
rect 18879 6846 19000 6874
rect 18730 6714 19000 6846
rect 18730 6686 18851 6714
rect 18879 6686 19000 6714
rect 18730 6554 19000 6686
rect 18730 6526 18851 6554
rect 18879 6526 19000 6554
rect 18730 6394 19000 6526
rect 18730 6366 18851 6394
rect 18879 6366 19000 6394
rect 18730 6234 19000 6366
rect 18730 6206 18851 6234
rect 18879 6206 19000 6234
rect 18730 6074 19000 6206
rect 18730 6046 18851 6074
rect 18879 6046 19000 6074
rect 18730 5914 19000 6046
rect 18730 5886 18851 5914
rect 18879 5886 19000 5914
rect 18730 5770 19000 5886
rect 15000 5754 19000 5770
rect 15000 5726 15118 5754
rect 15146 5726 18851 5754
rect 18879 5726 19000 5754
rect 15000 5651 19000 5726
rect 15000 5623 15306 5651
rect 15334 5623 15466 5651
rect 15494 5623 15626 5651
rect 15654 5623 15786 5651
rect 15814 5623 15946 5651
rect 15974 5623 16106 5651
rect 16134 5623 16266 5651
rect 16294 5623 16426 5651
rect 16454 5623 16586 5651
rect 16614 5623 16746 5651
rect 16774 5623 16906 5651
rect 16934 5623 17066 5651
rect 17094 5623 17226 5651
rect 17254 5623 17386 5651
rect 17414 5623 17546 5651
rect 17574 5623 17706 5651
rect 17734 5623 17866 5651
rect 17894 5623 18026 5651
rect 18054 5623 18186 5651
rect 18214 5623 18346 5651
rect 18374 5623 18506 5651
rect 18534 5623 18666 5651
rect 18694 5623 19000 5651
rect 15000 5500 19000 5623
rect 21000 9379 25000 9500
rect 21000 9351 21306 9379
rect 21334 9351 21466 9379
rect 21494 9351 21626 9379
rect 21654 9351 21786 9379
rect 21814 9351 21946 9379
rect 21974 9351 22106 9379
rect 22134 9351 22266 9379
rect 22294 9351 22426 9379
rect 22454 9351 22586 9379
rect 22614 9351 22746 9379
rect 22774 9351 22906 9379
rect 22934 9351 23066 9379
rect 23094 9351 23226 9379
rect 23254 9351 23386 9379
rect 23414 9351 23546 9379
rect 23574 9351 23706 9379
rect 23734 9351 23866 9379
rect 23894 9351 24026 9379
rect 24054 9351 24186 9379
rect 24214 9351 24346 9379
rect 24374 9351 24506 9379
rect 24534 9351 24666 9379
rect 24694 9351 25000 9379
rect 21000 9274 25000 9351
rect 21000 9246 21118 9274
rect 21146 9246 24851 9274
rect 24879 9246 25000 9274
rect 21000 9230 25000 9246
rect 21000 9114 21270 9230
rect 21000 9086 21118 9114
rect 21146 9086 21270 9114
rect 21000 8954 21270 9086
rect 21000 8926 21118 8954
rect 21146 8926 21270 8954
rect 21000 8794 21270 8926
rect 21000 8766 21118 8794
rect 21146 8766 21270 8794
rect 21000 8634 21270 8766
rect 21000 8606 21118 8634
rect 21146 8606 21270 8634
rect 21000 8474 21270 8606
rect 21000 8446 21118 8474
rect 21146 8446 21270 8474
rect 21000 8314 21270 8446
rect 21000 8286 21118 8314
rect 21146 8286 21270 8314
rect 21000 8154 21270 8286
rect 21000 8126 21118 8154
rect 21146 8126 21270 8154
rect 21000 7994 21270 8126
rect 21000 7966 21118 7994
rect 21146 7966 21270 7994
rect 21000 7834 21270 7966
rect 21000 7806 21118 7834
rect 21146 7806 21270 7834
rect 21000 7674 21270 7806
rect 21000 7646 21118 7674
rect 21146 7646 21270 7674
rect 21000 7514 21270 7646
rect 21000 7486 21118 7514
rect 21146 7486 21270 7514
rect 21000 7354 21270 7486
rect 21000 7326 21118 7354
rect 21146 7326 21270 7354
rect 21000 7194 21270 7326
rect 21000 7166 21118 7194
rect 21146 7166 21270 7194
rect 21000 7034 21270 7166
rect 21000 7006 21118 7034
rect 21146 7006 21270 7034
rect 21000 6874 21270 7006
rect 21000 6846 21118 6874
rect 21146 6846 21270 6874
rect 21000 6714 21270 6846
rect 21000 6686 21118 6714
rect 21146 6686 21270 6714
rect 21000 6554 21270 6686
rect 21000 6526 21118 6554
rect 21146 6526 21270 6554
rect 21000 6394 21270 6526
rect 21000 6366 21118 6394
rect 21146 6366 21270 6394
rect 21000 6234 21270 6366
rect 21000 6206 21118 6234
rect 21146 6206 21270 6234
rect 21000 6074 21270 6206
rect 21000 6046 21118 6074
rect 21146 6046 21270 6074
rect 21000 5914 21270 6046
rect 21000 5886 21118 5914
rect 21146 5886 21270 5914
rect 21000 5770 21270 5886
rect 24730 9114 25000 9230
rect 24730 9086 24851 9114
rect 24879 9086 25000 9114
rect 24730 8954 25000 9086
rect 24730 8926 24851 8954
rect 24879 8926 25000 8954
rect 24730 8794 25000 8926
rect 24730 8766 24851 8794
rect 24879 8766 25000 8794
rect 24730 8634 25000 8766
rect 24730 8606 24851 8634
rect 24879 8606 25000 8634
rect 24730 8474 25000 8606
rect 24730 8446 24851 8474
rect 24879 8446 25000 8474
rect 24730 8314 25000 8446
rect 24730 8286 24851 8314
rect 24879 8286 25000 8314
rect 24730 8154 25000 8286
rect 24730 8126 24851 8154
rect 24879 8126 25000 8154
rect 24730 7994 25000 8126
rect 24730 7966 24851 7994
rect 24879 7966 25000 7994
rect 24730 7834 25000 7966
rect 24730 7806 24851 7834
rect 24879 7806 25000 7834
rect 24730 7674 25000 7806
rect 24730 7646 24851 7674
rect 24879 7646 25000 7674
rect 24730 7514 25000 7646
rect 24730 7486 24851 7514
rect 24879 7486 25000 7514
rect 24730 7354 25000 7486
rect 24730 7326 24851 7354
rect 24879 7326 25000 7354
rect 24730 7194 25000 7326
rect 24730 7166 24851 7194
rect 24879 7166 25000 7194
rect 24730 7034 25000 7166
rect 24730 7006 24851 7034
rect 24879 7006 25000 7034
rect 24730 6874 25000 7006
rect 24730 6846 24851 6874
rect 24879 6846 25000 6874
rect 24730 6714 25000 6846
rect 24730 6686 24851 6714
rect 24879 6686 25000 6714
rect 24730 6554 25000 6686
rect 24730 6526 24851 6554
rect 24879 6526 25000 6554
rect 24730 6394 25000 6526
rect 24730 6366 24851 6394
rect 24879 6366 25000 6394
rect 24730 6234 25000 6366
rect 24730 6206 24851 6234
rect 24879 6206 25000 6234
rect 24730 6074 25000 6206
rect 24730 6046 24851 6074
rect 24879 6046 25000 6074
rect 24730 5914 25000 6046
rect 24730 5886 24851 5914
rect 24879 5886 25000 5914
rect 24730 5770 25000 5886
rect 21000 5754 25000 5770
rect 21000 5726 21118 5754
rect 21146 5726 24851 5754
rect 24879 5726 25000 5754
rect 21000 5651 25000 5726
rect 21000 5623 21306 5651
rect 21334 5623 21466 5651
rect 21494 5623 21626 5651
rect 21654 5623 21786 5651
rect 21814 5623 21946 5651
rect 21974 5623 22106 5651
rect 22134 5623 22266 5651
rect 22294 5623 22426 5651
rect 22454 5623 22586 5651
rect 22614 5623 22746 5651
rect 22774 5623 22906 5651
rect 22934 5623 23066 5651
rect 23094 5623 23226 5651
rect 23254 5623 23386 5651
rect 23414 5623 23546 5651
rect 23574 5623 23706 5651
rect 23734 5623 23866 5651
rect 23894 5623 24026 5651
rect 24054 5623 24186 5651
rect 24214 5623 24346 5651
rect 24374 5623 24506 5651
rect 24534 5623 24666 5651
rect 24694 5623 25000 5651
rect 21000 5500 25000 5623
rect 3000 3379 7000 3500
rect 3000 3351 3306 3379
rect 3334 3351 3466 3379
rect 3494 3351 3626 3379
rect 3654 3351 3786 3379
rect 3814 3351 3946 3379
rect 3974 3351 4106 3379
rect 4134 3351 4266 3379
rect 4294 3351 4426 3379
rect 4454 3351 4586 3379
rect 4614 3351 4746 3379
rect 4774 3351 4906 3379
rect 4934 3351 5066 3379
rect 5094 3351 5226 3379
rect 5254 3351 5386 3379
rect 5414 3351 5546 3379
rect 5574 3351 5706 3379
rect 5734 3351 5866 3379
rect 5894 3351 6026 3379
rect 6054 3351 6186 3379
rect 6214 3351 6346 3379
rect 6374 3351 6506 3379
rect 6534 3351 6666 3379
rect 6694 3351 7000 3379
rect 3000 3274 7000 3351
rect 3000 3246 3118 3274
rect 3146 3246 6851 3274
rect 6879 3246 7000 3274
rect 3000 3230 7000 3246
rect 3000 3114 3270 3230
rect 3000 3086 3118 3114
rect 3146 3086 3270 3114
rect 3000 2954 3270 3086
rect 3000 2926 3118 2954
rect 3146 2926 3270 2954
rect 3000 2794 3270 2926
rect 3000 2766 3118 2794
rect 3146 2766 3270 2794
rect 3000 2634 3270 2766
rect 3000 2606 3118 2634
rect 3146 2606 3270 2634
rect 3000 2474 3270 2606
rect 3000 2446 3118 2474
rect 3146 2446 3270 2474
rect 3000 2314 3270 2446
rect 3000 2286 3118 2314
rect 3146 2286 3270 2314
rect 3000 2154 3270 2286
rect 3000 2126 3118 2154
rect 3146 2126 3270 2154
rect 3000 1994 3270 2126
rect 3000 1966 3118 1994
rect 3146 1966 3270 1994
rect 3000 1834 3270 1966
rect 3000 1806 3118 1834
rect 3146 1806 3270 1834
rect 3000 1674 3270 1806
rect 3000 1646 3118 1674
rect 3146 1646 3270 1674
rect 3000 1514 3270 1646
rect 3000 1486 3118 1514
rect 3146 1486 3270 1514
rect 3000 1354 3270 1486
rect 3000 1326 3118 1354
rect 3146 1326 3270 1354
rect 3000 1194 3270 1326
rect 3000 1166 3118 1194
rect 3146 1166 3270 1194
rect 3000 1034 3270 1166
rect 3000 1006 3118 1034
rect 3146 1006 3270 1034
rect 3000 874 3270 1006
rect 3000 846 3118 874
rect 3146 846 3270 874
rect 3000 714 3270 846
rect 3000 686 3118 714
rect 3146 686 3270 714
rect 3000 554 3270 686
rect 3000 526 3118 554
rect 3146 526 3270 554
rect 3000 394 3270 526
rect 3000 366 3118 394
rect 3146 366 3270 394
rect 3000 234 3270 366
rect 3000 206 3118 234
rect 3146 206 3270 234
rect 3000 74 3270 206
rect 3000 46 3118 74
rect 3146 46 3270 74
rect 3000 -86 3270 46
rect 3000 -114 3118 -86
rect 3146 -114 3270 -86
rect 3000 -230 3270 -114
rect 6730 3114 7000 3230
rect 6730 3086 6851 3114
rect 6879 3086 7000 3114
rect 6730 2954 7000 3086
rect 6730 2926 6851 2954
rect 6879 2926 7000 2954
rect 6730 2794 7000 2926
rect 6730 2766 6851 2794
rect 6879 2766 7000 2794
rect 6730 2634 7000 2766
rect 6730 2606 6851 2634
rect 6879 2606 7000 2634
rect 6730 2474 7000 2606
rect 6730 2446 6851 2474
rect 6879 2446 7000 2474
rect 6730 2314 7000 2446
rect 6730 2286 6851 2314
rect 6879 2286 7000 2314
rect 6730 2154 7000 2286
rect 6730 2126 6851 2154
rect 6879 2126 7000 2154
rect 6730 1994 7000 2126
rect 6730 1966 6851 1994
rect 6879 1966 7000 1994
rect 6730 1834 7000 1966
rect 6730 1806 6851 1834
rect 6879 1806 7000 1834
rect 6730 1674 7000 1806
rect 6730 1646 6851 1674
rect 6879 1646 7000 1674
rect 6730 1514 7000 1646
rect 6730 1486 6851 1514
rect 6879 1486 7000 1514
rect 6730 1354 7000 1486
rect 6730 1326 6851 1354
rect 6879 1326 7000 1354
rect 6730 1194 7000 1326
rect 6730 1166 6851 1194
rect 6879 1166 7000 1194
rect 6730 1034 7000 1166
rect 6730 1006 6851 1034
rect 6879 1006 7000 1034
rect 6730 874 7000 1006
rect 6730 846 6851 874
rect 6879 846 7000 874
rect 6730 714 7000 846
rect 6730 686 6851 714
rect 6879 686 7000 714
rect 6730 554 7000 686
rect 6730 526 6851 554
rect 6879 526 7000 554
rect 6730 394 7000 526
rect 6730 366 6851 394
rect 6879 366 7000 394
rect 6730 234 7000 366
rect 6730 206 6851 234
rect 6879 206 7000 234
rect 6730 74 7000 206
rect 6730 46 6851 74
rect 6879 46 7000 74
rect 6730 -86 7000 46
rect 6730 -114 6851 -86
rect 6879 -114 7000 -86
rect 6730 -230 7000 -114
rect 3000 -246 7000 -230
rect 3000 -274 3118 -246
rect 3146 -274 6851 -246
rect 6879 -274 7000 -246
rect 3000 -349 7000 -274
rect 3000 -377 3306 -349
rect 3334 -377 3466 -349
rect 3494 -377 3626 -349
rect 3654 -377 3786 -349
rect 3814 -377 3946 -349
rect 3974 -377 4106 -349
rect 4134 -377 4266 -349
rect 4294 -377 4426 -349
rect 4454 -377 4586 -349
rect 4614 -377 4746 -349
rect 4774 -377 4906 -349
rect 4934 -377 5066 -349
rect 5094 -377 5226 -349
rect 5254 -377 5386 -349
rect 5414 -377 5546 -349
rect 5574 -377 5706 -349
rect 5734 -377 5866 -349
rect 5894 -377 6026 -349
rect 6054 -377 6186 -349
rect 6214 -377 6346 -349
rect 6374 -377 6506 -349
rect 6534 -377 6666 -349
rect 6694 -377 7000 -349
rect 3000 -500 7000 -377
rect 9000 3379 13000 3500
rect 9000 3351 9306 3379
rect 9334 3351 9466 3379
rect 9494 3351 9626 3379
rect 9654 3351 9786 3379
rect 9814 3351 9946 3379
rect 9974 3351 10106 3379
rect 10134 3351 10266 3379
rect 10294 3351 10426 3379
rect 10454 3351 10586 3379
rect 10614 3351 10746 3379
rect 10774 3351 10906 3379
rect 10934 3351 11066 3379
rect 11094 3351 11226 3379
rect 11254 3351 11386 3379
rect 11414 3351 11546 3379
rect 11574 3351 11706 3379
rect 11734 3351 11866 3379
rect 11894 3351 12026 3379
rect 12054 3351 12186 3379
rect 12214 3351 12346 3379
rect 12374 3351 12506 3379
rect 12534 3351 12666 3379
rect 12694 3351 13000 3379
rect 9000 3274 13000 3351
rect 9000 3246 9118 3274
rect 9146 3246 12851 3274
rect 12879 3246 13000 3274
rect 9000 3230 13000 3246
rect 9000 3114 9270 3230
rect 9000 3086 9118 3114
rect 9146 3086 9270 3114
rect 9000 2954 9270 3086
rect 9000 2926 9118 2954
rect 9146 2926 9270 2954
rect 9000 2794 9270 2926
rect 9000 2766 9118 2794
rect 9146 2766 9270 2794
rect 9000 2634 9270 2766
rect 9000 2606 9118 2634
rect 9146 2606 9270 2634
rect 9000 2474 9270 2606
rect 9000 2446 9118 2474
rect 9146 2446 9270 2474
rect 9000 2314 9270 2446
rect 9000 2286 9118 2314
rect 9146 2286 9270 2314
rect 9000 2154 9270 2286
rect 9000 2126 9118 2154
rect 9146 2126 9270 2154
rect 9000 1994 9270 2126
rect 9000 1966 9118 1994
rect 9146 1966 9270 1994
rect 9000 1834 9270 1966
rect 9000 1806 9118 1834
rect 9146 1806 9270 1834
rect 9000 1674 9270 1806
rect 9000 1646 9118 1674
rect 9146 1646 9270 1674
rect 9000 1514 9270 1646
rect 9000 1486 9118 1514
rect 9146 1486 9270 1514
rect 9000 1354 9270 1486
rect 9000 1326 9118 1354
rect 9146 1326 9270 1354
rect 9000 1194 9270 1326
rect 9000 1166 9118 1194
rect 9146 1166 9270 1194
rect 9000 1034 9270 1166
rect 9000 1006 9118 1034
rect 9146 1006 9270 1034
rect 9000 874 9270 1006
rect 9000 846 9118 874
rect 9146 846 9270 874
rect 9000 714 9270 846
rect 9000 686 9118 714
rect 9146 686 9270 714
rect 9000 554 9270 686
rect 9000 526 9118 554
rect 9146 526 9270 554
rect 9000 394 9270 526
rect 9000 366 9118 394
rect 9146 366 9270 394
rect 9000 234 9270 366
rect 9000 206 9118 234
rect 9146 206 9270 234
rect 9000 74 9270 206
rect 9000 46 9118 74
rect 9146 46 9270 74
rect 9000 -86 9270 46
rect 9000 -114 9118 -86
rect 9146 -114 9270 -86
rect 9000 -230 9270 -114
rect 12730 3114 13000 3230
rect 12730 3086 12851 3114
rect 12879 3086 13000 3114
rect 12730 2954 13000 3086
rect 12730 2926 12851 2954
rect 12879 2926 13000 2954
rect 12730 2794 13000 2926
rect 12730 2766 12851 2794
rect 12879 2766 13000 2794
rect 12730 2634 13000 2766
rect 12730 2606 12851 2634
rect 12879 2606 13000 2634
rect 12730 2474 13000 2606
rect 12730 2446 12851 2474
rect 12879 2446 13000 2474
rect 12730 2314 13000 2446
rect 12730 2286 12851 2314
rect 12879 2286 13000 2314
rect 12730 2154 13000 2286
rect 12730 2126 12851 2154
rect 12879 2126 13000 2154
rect 12730 1994 13000 2126
rect 12730 1966 12851 1994
rect 12879 1966 13000 1994
rect 12730 1834 13000 1966
rect 12730 1806 12851 1834
rect 12879 1806 13000 1834
rect 12730 1674 13000 1806
rect 12730 1646 12851 1674
rect 12879 1646 13000 1674
rect 12730 1514 13000 1646
rect 12730 1486 12851 1514
rect 12879 1486 13000 1514
rect 12730 1354 13000 1486
rect 12730 1326 12851 1354
rect 12879 1326 13000 1354
rect 12730 1194 13000 1326
rect 12730 1166 12851 1194
rect 12879 1166 13000 1194
rect 12730 1034 13000 1166
rect 12730 1006 12851 1034
rect 12879 1006 13000 1034
rect 12730 874 13000 1006
rect 12730 846 12851 874
rect 12879 846 13000 874
rect 12730 714 13000 846
rect 12730 686 12851 714
rect 12879 686 13000 714
rect 12730 554 13000 686
rect 12730 526 12851 554
rect 12879 526 13000 554
rect 12730 394 13000 526
rect 12730 366 12851 394
rect 12879 366 13000 394
rect 12730 234 13000 366
rect 12730 206 12851 234
rect 12879 206 13000 234
rect 12730 74 13000 206
rect 12730 46 12851 74
rect 12879 46 13000 74
rect 12730 -86 13000 46
rect 12730 -114 12851 -86
rect 12879 -114 13000 -86
rect 12730 -230 13000 -114
rect 9000 -246 13000 -230
rect 9000 -274 9118 -246
rect 9146 -274 12851 -246
rect 12879 -274 13000 -246
rect 9000 -349 13000 -274
rect 9000 -377 9306 -349
rect 9334 -377 9466 -349
rect 9494 -377 9626 -349
rect 9654 -377 9786 -349
rect 9814 -377 9946 -349
rect 9974 -377 10106 -349
rect 10134 -377 10266 -349
rect 10294 -377 10426 -349
rect 10454 -377 10586 -349
rect 10614 -377 10746 -349
rect 10774 -377 10906 -349
rect 10934 -377 11066 -349
rect 11094 -377 11226 -349
rect 11254 -377 11386 -349
rect 11414 -377 11546 -349
rect 11574 -377 11706 -349
rect 11734 -377 11866 -349
rect 11894 -377 12026 -349
rect 12054 -377 12186 -349
rect 12214 -377 12346 -349
rect 12374 -377 12506 -349
rect 12534 -377 12666 -349
rect 12694 -377 13000 -349
rect 9000 -500 13000 -377
rect 15000 3379 19000 3500
rect 15000 3351 15306 3379
rect 15334 3351 15466 3379
rect 15494 3351 15626 3379
rect 15654 3351 15786 3379
rect 15814 3351 15946 3379
rect 15974 3351 16106 3379
rect 16134 3351 16266 3379
rect 16294 3351 16426 3379
rect 16454 3351 16586 3379
rect 16614 3351 16746 3379
rect 16774 3351 16906 3379
rect 16934 3351 17066 3379
rect 17094 3351 17226 3379
rect 17254 3351 17386 3379
rect 17414 3351 17546 3379
rect 17574 3351 17706 3379
rect 17734 3351 17866 3379
rect 17894 3351 18026 3379
rect 18054 3351 18186 3379
rect 18214 3351 18346 3379
rect 18374 3351 18506 3379
rect 18534 3351 18666 3379
rect 18694 3351 19000 3379
rect 15000 3274 19000 3351
rect 15000 3246 15118 3274
rect 15146 3246 18851 3274
rect 18879 3246 19000 3274
rect 15000 3230 19000 3246
rect 15000 3114 15270 3230
rect 15000 3086 15118 3114
rect 15146 3086 15270 3114
rect 15000 2954 15270 3086
rect 15000 2926 15118 2954
rect 15146 2926 15270 2954
rect 15000 2794 15270 2926
rect 15000 2766 15118 2794
rect 15146 2766 15270 2794
rect 15000 2634 15270 2766
rect 15000 2606 15118 2634
rect 15146 2606 15270 2634
rect 15000 2474 15270 2606
rect 15000 2446 15118 2474
rect 15146 2446 15270 2474
rect 15000 2314 15270 2446
rect 15000 2286 15118 2314
rect 15146 2286 15270 2314
rect 15000 2154 15270 2286
rect 15000 2126 15118 2154
rect 15146 2126 15270 2154
rect 15000 1994 15270 2126
rect 15000 1966 15118 1994
rect 15146 1966 15270 1994
rect 15000 1834 15270 1966
rect 15000 1806 15118 1834
rect 15146 1806 15270 1834
rect 15000 1674 15270 1806
rect 15000 1646 15118 1674
rect 15146 1646 15270 1674
rect 15000 1514 15270 1646
rect 15000 1486 15118 1514
rect 15146 1486 15270 1514
rect 15000 1354 15270 1486
rect 15000 1326 15118 1354
rect 15146 1326 15270 1354
rect 15000 1194 15270 1326
rect 15000 1166 15118 1194
rect 15146 1166 15270 1194
rect 15000 1034 15270 1166
rect 15000 1006 15118 1034
rect 15146 1006 15270 1034
rect 15000 874 15270 1006
rect 15000 846 15118 874
rect 15146 846 15270 874
rect 15000 714 15270 846
rect 15000 686 15118 714
rect 15146 686 15270 714
rect 15000 554 15270 686
rect 15000 526 15118 554
rect 15146 526 15270 554
rect 15000 394 15270 526
rect 15000 366 15118 394
rect 15146 366 15270 394
rect 15000 234 15270 366
rect 15000 206 15118 234
rect 15146 206 15270 234
rect 15000 74 15270 206
rect 15000 46 15118 74
rect 15146 46 15270 74
rect 15000 -86 15270 46
rect 15000 -114 15118 -86
rect 15146 -114 15270 -86
rect 15000 -230 15270 -114
rect 18730 3114 19000 3230
rect 18730 3086 18851 3114
rect 18879 3086 19000 3114
rect 18730 2954 19000 3086
rect 18730 2926 18851 2954
rect 18879 2926 19000 2954
rect 18730 2794 19000 2926
rect 18730 2766 18851 2794
rect 18879 2766 19000 2794
rect 18730 2634 19000 2766
rect 18730 2606 18851 2634
rect 18879 2606 19000 2634
rect 18730 2474 19000 2606
rect 18730 2446 18851 2474
rect 18879 2446 19000 2474
rect 18730 2314 19000 2446
rect 18730 2286 18851 2314
rect 18879 2286 19000 2314
rect 18730 2154 19000 2286
rect 18730 2126 18851 2154
rect 18879 2126 19000 2154
rect 18730 1994 19000 2126
rect 18730 1966 18851 1994
rect 18879 1966 19000 1994
rect 18730 1834 19000 1966
rect 18730 1806 18851 1834
rect 18879 1806 19000 1834
rect 18730 1674 19000 1806
rect 18730 1646 18851 1674
rect 18879 1646 19000 1674
rect 18730 1514 19000 1646
rect 18730 1486 18851 1514
rect 18879 1486 19000 1514
rect 18730 1354 19000 1486
rect 18730 1326 18851 1354
rect 18879 1326 19000 1354
rect 18730 1194 19000 1326
rect 18730 1166 18851 1194
rect 18879 1166 19000 1194
rect 18730 1034 19000 1166
rect 18730 1006 18851 1034
rect 18879 1006 19000 1034
rect 18730 874 19000 1006
rect 18730 846 18851 874
rect 18879 846 19000 874
rect 18730 714 19000 846
rect 18730 686 18851 714
rect 18879 686 19000 714
rect 18730 554 19000 686
rect 18730 526 18851 554
rect 18879 526 19000 554
rect 18730 394 19000 526
rect 18730 366 18851 394
rect 18879 366 19000 394
rect 18730 234 19000 366
rect 18730 206 18851 234
rect 18879 206 19000 234
rect 18730 74 19000 206
rect 18730 46 18851 74
rect 18879 46 19000 74
rect 18730 -86 19000 46
rect 18730 -114 18851 -86
rect 18879 -114 19000 -86
rect 18730 -230 19000 -114
rect 15000 -246 19000 -230
rect 15000 -274 15118 -246
rect 15146 -274 18851 -246
rect 18879 -274 19000 -246
rect 15000 -349 19000 -274
rect 21000 3379 25000 3500
rect 21000 3351 21306 3379
rect 21334 3351 21466 3379
rect 21494 3351 21626 3379
rect 21654 3351 21786 3379
rect 21814 3351 21946 3379
rect 21974 3351 22106 3379
rect 22134 3351 22266 3379
rect 22294 3351 22426 3379
rect 22454 3351 22586 3379
rect 22614 3351 22746 3379
rect 22774 3351 22906 3379
rect 22934 3351 23066 3379
rect 23094 3351 23226 3379
rect 23254 3351 23386 3379
rect 23414 3351 23546 3379
rect 23574 3351 23706 3379
rect 23734 3351 23866 3379
rect 23894 3351 24026 3379
rect 24054 3351 24186 3379
rect 24214 3351 24346 3379
rect 24374 3351 24506 3379
rect 24534 3351 24666 3379
rect 24694 3351 25000 3379
rect 21000 3274 25000 3351
rect 21000 3246 21118 3274
rect 21146 3246 24851 3274
rect 24879 3246 25000 3274
rect 21000 3230 25000 3246
rect 21000 3114 21270 3230
rect 21000 3086 21118 3114
rect 21146 3086 21270 3114
rect 21000 2954 21270 3086
rect 21000 2926 21118 2954
rect 21146 2926 21270 2954
rect 21000 2794 21270 2926
rect 21000 2766 21118 2794
rect 21146 2766 21270 2794
rect 21000 2634 21270 2766
rect 21000 2606 21118 2634
rect 21146 2606 21270 2634
rect 21000 2474 21270 2606
rect 21000 2446 21118 2474
rect 21146 2446 21270 2474
rect 21000 2314 21270 2446
rect 21000 2286 21118 2314
rect 21146 2286 21270 2314
rect 21000 2154 21270 2286
rect 21000 2126 21118 2154
rect 21146 2126 21270 2154
rect 21000 1994 21270 2126
rect 21000 1966 21118 1994
rect 21146 1966 21270 1994
rect 21000 1834 21270 1966
rect 21000 1806 21118 1834
rect 21146 1806 21270 1834
rect 21000 1674 21270 1806
rect 21000 1646 21118 1674
rect 21146 1646 21270 1674
rect 21000 1514 21270 1646
rect 21000 1486 21118 1514
rect 21146 1486 21270 1514
rect 21000 1354 21270 1486
rect 21000 1326 21118 1354
rect 21146 1326 21270 1354
rect 21000 1194 21270 1326
rect 21000 1166 21118 1194
rect 21146 1166 21270 1194
rect 21000 1034 21270 1166
rect 21000 1006 21118 1034
rect 21146 1006 21270 1034
rect 21000 874 21270 1006
rect 21000 846 21118 874
rect 21146 846 21270 874
rect 21000 714 21270 846
rect 21000 686 21118 714
rect 21146 686 21270 714
rect 21000 554 21270 686
rect 21000 526 21118 554
rect 21146 526 21270 554
rect 21000 394 21270 526
rect 21000 366 21118 394
rect 21146 366 21270 394
rect 21000 234 21270 366
rect 21000 206 21118 234
rect 21146 206 21270 234
rect 21000 74 21270 206
rect 21000 46 21118 74
rect 21146 46 21270 74
rect 21000 -86 21270 46
rect 21000 -114 21118 -86
rect 21146 -114 21270 -86
rect 21000 -230 21270 -114
rect 24730 3114 25000 3230
rect 24730 3086 24851 3114
rect 24879 3086 25000 3114
rect 24730 2954 25000 3086
rect 24730 2926 24851 2954
rect 24879 2926 25000 2954
rect 24730 2794 25000 2926
rect 24730 2766 24851 2794
rect 24879 2766 25000 2794
rect 24730 2634 25000 2766
rect 24730 2606 24851 2634
rect 24879 2606 25000 2634
rect 24730 2474 25000 2606
rect 24730 2446 24851 2474
rect 24879 2446 25000 2474
rect 24730 2314 25000 2446
rect 24730 2286 24851 2314
rect 24879 2286 25000 2314
rect 24730 2154 25000 2286
rect 24730 2126 24851 2154
rect 24879 2126 25000 2154
rect 24730 1994 25000 2126
rect 24730 1966 24851 1994
rect 24879 1966 25000 1994
rect 24730 1834 25000 1966
rect 24730 1806 24851 1834
rect 24879 1806 25000 1834
rect 24730 1674 25000 1806
rect 24730 1646 24851 1674
rect 24879 1646 25000 1674
rect 24730 1514 25000 1646
rect 24730 1486 24851 1514
rect 24879 1486 25000 1514
rect 24730 1354 25000 1486
rect 24730 1326 24851 1354
rect 24879 1326 25000 1354
rect 24730 1194 25000 1326
rect 24730 1166 24851 1194
rect 24879 1166 25000 1194
rect 24730 1034 25000 1166
rect 24730 1006 24851 1034
rect 24879 1006 25000 1034
rect 24730 874 25000 1006
rect 24730 846 24851 874
rect 24879 846 25000 874
rect 24730 714 25000 846
rect 24730 686 24851 714
rect 24879 686 25000 714
rect 24730 554 25000 686
rect 24730 526 24851 554
rect 24879 526 25000 554
rect 24730 394 25000 526
rect 24730 366 24851 394
rect 24879 366 25000 394
rect 24730 234 25000 366
rect 24730 206 24851 234
rect 24879 206 25000 234
rect 24730 74 25000 206
rect 24730 46 24851 74
rect 24879 46 25000 74
rect 24730 -86 25000 46
rect 24730 -114 24851 -86
rect 24879 -114 25000 -86
rect 24730 -230 25000 -114
rect 21000 -246 25000 -230
rect 21000 -274 21118 -246
rect 21146 -274 24851 -246
rect 24879 -274 25000 -246
rect 21000 -345 25000 -274
rect 15000 -377 15306 -349
rect 15334 -377 15466 -349
rect 15494 -377 15626 -349
rect 15654 -377 15786 -349
rect 15814 -377 15946 -349
rect 15974 -377 16106 -349
rect 16134 -377 16266 -349
rect 16294 -377 16426 -349
rect 16454 -377 16586 -349
rect 16614 -377 16746 -349
rect 16774 -377 16906 -349
rect 16934 -377 17066 -349
rect 17094 -377 17226 -349
rect 17254 -377 17386 -349
rect 17414 -377 17546 -349
rect 17574 -377 17706 -349
rect 17734 -377 17866 -349
rect 17894 -377 18026 -349
rect 18054 -377 18186 -349
rect 18214 -377 18346 -349
rect 18374 -377 18506 -349
rect 18534 -377 18666 -349
rect 18694 -377 19000 -349
rect 15000 -500 19000 -377
rect 19915 -349 25000 -345
rect 19915 -377 21306 -349
rect 21334 -377 21466 -349
rect 21494 -377 21626 -349
rect 21654 -377 21786 -349
rect 21814 -377 21946 -349
rect 21974 -377 22106 -349
rect 22134 -377 22266 -349
rect 22294 -377 22426 -349
rect 22454 -377 22586 -349
rect 22614 -377 22746 -349
rect 22774 -377 22906 -349
rect 22934 -377 23066 -349
rect 23094 -377 23226 -349
rect 23254 -377 23386 -349
rect 23414 -377 23546 -349
rect 23574 -377 23706 -349
rect 23734 -377 23866 -349
rect 23894 -377 24026 -349
rect 24054 -377 24186 -349
rect 24214 -377 24346 -349
rect 24374 -377 24506 -349
rect 24534 -377 24666 -349
rect 24694 -377 25000 -349
rect 19915 -445 25000 -377
rect 19915 -570 20025 -445
rect 21000 -500 25000 -445
rect 19240 -575 19295 -570
rect 19240 -745 19245 -575
rect 19290 -745 19295 -575
rect 19595 -575 20025 -570
rect 19430 -630 19490 -625
rect 19430 -690 19435 -630
rect 19485 -690 19490 -630
rect 19430 -695 19490 -690
rect 19240 -1250 19295 -745
rect 19595 -745 19600 -575
rect 19645 -745 20025 -575
rect 19595 -750 20025 -745
rect 20030 -1140 20070 -1135
rect 20030 -1170 20035 -1140
rect 20065 -1170 20070 -1140
rect 20030 -1175 20070 -1170
rect 20065 -1210 20105 -1205
rect 20065 -1240 20070 -1210
rect 20100 -1240 20105 -1210
rect 20065 -1245 20105 -1240
rect 10900 -1500 11700 -1400
rect 11600 -3600 11700 -1500
rect 16300 -1850 16950 -1750
rect 16300 -1950 16400 -1850
rect 16200 -2050 16250 -1950
rect 16350 -2050 16400 -1950
rect 16150 -2070 16230 -2065
rect 16150 -2100 16155 -2070
rect 16225 -2100 16230 -2070
rect 16150 -2140 16230 -2100
rect 16150 -2180 16155 -2140
rect 16225 -2180 16230 -2140
rect 16290 -2180 16295 -2140
rect 16365 -2180 16370 -2140
rect 16290 -2230 16370 -2180
rect 16290 -2260 16295 -2230
rect 16365 -2260 16370 -2230
rect 16290 -2265 16370 -2260
rect 16200 -2400 16250 -2300
rect 16350 -2400 16400 -2300
rect 11600 -3700 11650 -3600
rect 11750 -3700 11800 -3600
rect 11630 -3740 11710 -3735
rect 11630 -3770 11635 -3740
rect 11705 -3770 11710 -3740
rect 11630 -3820 11710 -3770
rect 11630 -3860 11635 -3820
rect 11705 -3860 11710 -3820
rect 11770 -3860 11775 -3820
rect 11845 -3860 11850 -3820
rect 11770 -3900 11850 -3860
rect 11770 -3930 11775 -3900
rect 11845 -3930 11850 -3900
rect 11770 -3935 11850 -3930
rect 11600 -4050 11650 -3950
rect 11750 -4050 11800 -3950
rect 11600 -4150 11700 -4050
rect 11050 -4250 11700 -4150
rect 16300 -4500 16400 -2400
rect 16300 -4600 17100 -4500
rect 8195 -4760 8235 -4755
rect 8195 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8195 -4795 8235 -4790
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 7975 -5255 8405 -5250
rect 7975 -5425 8355 -5255
rect 8400 -5425 8405 -5255
rect 8705 -5255 8760 -4750
rect 8510 -5310 8570 -5305
rect 8510 -5370 8515 -5310
rect 8565 -5370 8570 -5310
rect 8510 -5375 8570 -5370
rect 7975 -5430 8405 -5425
rect 8705 -5425 8710 -5255
rect 8755 -5425 8760 -5255
rect 8705 -5430 8760 -5425
rect 3000 -5555 7000 -5500
rect 7975 -5555 8085 -5430
rect 3000 -5623 8085 -5555
rect 3000 -5651 3306 -5623
rect 3334 -5651 3466 -5623
rect 3494 -5651 3626 -5623
rect 3654 -5651 3786 -5623
rect 3814 -5651 3946 -5623
rect 3974 -5651 4106 -5623
rect 4134 -5651 4266 -5623
rect 4294 -5651 4426 -5623
rect 4454 -5651 4586 -5623
rect 4614 -5651 4746 -5623
rect 4774 -5651 4906 -5623
rect 4934 -5651 5066 -5623
rect 5094 -5651 5226 -5623
rect 5254 -5651 5386 -5623
rect 5414 -5651 5546 -5623
rect 5574 -5651 5706 -5623
rect 5734 -5651 5866 -5623
rect 5894 -5651 6026 -5623
rect 6054 -5651 6186 -5623
rect 6214 -5651 6346 -5623
rect 6374 -5651 6506 -5623
rect 6534 -5651 6666 -5623
rect 6694 -5651 8085 -5623
rect 3000 -5655 8085 -5651
rect 9000 -5623 13000 -5500
rect 9000 -5651 9306 -5623
rect 9334 -5651 9466 -5623
rect 9494 -5651 9626 -5623
rect 9654 -5651 9786 -5623
rect 9814 -5651 9946 -5623
rect 9974 -5651 10106 -5623
rect 10134 -5651 10266 -5623
rect 10294 -5651 10426 -5623
rect 10454 -5651 10586 -5623
rect 10614 -5651 10746 -5623
rect 10774 -5651 10906 -5623
rect 10934 -5651 11066 -5623
rect 11094 -5651 11226 -5623
rect 11254 -5651 11386 -5623
rect 11414 -5651 11546 -5623
rect 11574 -5651 11706 -5623
rect 11734 -5651 11866 -5623
rect 11894 -5651 12026 -5623
rect 12054 -5651 12186 -5623
rect 12214 -5651 12346 -5623
rect 12374 -5651 12506 -5623
rect 12534 -5651 12666 -5623
rect 12694 -5651 13000 -5623
rect 3000 -5726 7000 -5655
rect 3000 -5754 3121 -5726
rect 3149 -5754 6854 -5726
rect 6882 -5754 7000 -5726
rect 3000 -5770 7000 -5754
rect 3000 -5886 3270 -5770
rect 3000 -5914 3121 -5886
rect 3149 -5914 3270 -5886
rect 3000 -6046 3270 -5914
rect 3000 -6074 3121 -6046
rect 3149 -6074 3270 -6046
rect 3000 -6206 3270 -6074
rect 3000 -6234 3121 -6206
rect 3149 -6234 3270 -6206
rect 3000 -6366 3270 -6234
rect 3000 -6394 3121 -6366
rect 3149 -6394 3270 -6366
rect 3000 -6526 3270 -6394
rect 3000 -6554 3121 -6526
rect 3149 -6554 3270 -6526
rect 3000 -6686 3270 -6554
rect 3000 -6714 3121 -6686
rect 3149 -6714 3270 -6686
rect 3000 -6846 3270 -6714
rect 3000 -6874 3121 -6846
rect 3149 -6874 3270 -6846
rect 3000 -7006 3270 -6874
rect 3000 -7034 3121 -7006
rect 3149 -7034 3270 -7006
rect 3000 -7166 3270 -7034
rect 3000 -7194 3121 -7166
rect 3149 -7194 3270 -7166
rect 3000 -7326 3270 -7194
rect 3000 -7354 3121 -7326
rect 3149 -7354 3270 -7326
rect 3000 -7486 3270 -7354
rect 3000 -7514 3121 -7486
rect 3149 -7514 3270 -7486
rect 3000 -7646 3270 -7514
rect 3000 -7674 3121 -7646
rect 3149 -7674 3270 -7646
rect 3000 -7806 3270 -7674
rect 3000 -7834 3121 -7806
rect 3149 -7834 3270 -7806
rect 3000 -7966 3270 -7834
rect 3000 -7994 3121 -7966
rect 3149 -7994 3270 -7966
rect 3000 -8126 3270 -7994
rect 3000 -8154 3121 -8126
rect 3149 -8154 3270 -8126
rect 3000 -8286 3270 -8154
rect 3000 -8314 3121 -8286
rect 3149 -8314 3270 -8286
rect 3000 -8446 3270 -8314
rect 3000 -8474 3121 -8446
rect 3149 -8474 3270 -8446
rect 3000 -8606 3270 -8474
rect 3000 -8634 3121 -8606
rect 3149 -8634 3270 -8606
rect 3000 -8766 3270 -8634
rect 3000 -8794 3121 -8766
rect 3149 -8794 3270 -8766
rect 3000 -8926 3270 -8794
rect 3000 -8954 3121 -8926
rect 3149 -8954 3270 -8926
rect 3000 -9086 3270 -8954
rect 3000 -9114 3121 -9086
rect 3149 -9114 3270 -9086
rect 3000 -9230 3270 -9114
rect 6730 -5886 7000 -5770
rect 6730 -5914 6854 -5886
rect 6882 -5914 7000 -5886
rect 6730 -6046 7000 -5914
rect 6730 -6074 6854 -6046
rect 6882 -6074 7000 -6046
rect 6730 -6206 7000 -6074
rect 6730 -6234 6854 -6206
rect 6882 -6234 7000 -6206
rect 6730 -6366 7000 -6234
rect 6730 -6394 6854 -6366
rect 6882 -6394 7000 -6366
rect 6730 -6526 7000 -6394
rect 6730 -6554 6854 -6526
rect 6882 -6554 7000 -6526
rect 6730 -6686 7000 -6554
rect 6730 -6714 6854 -6686
rect 6882 -6714 7000 -6686
rect 6730 -6846 7000 -6714
rect 6730 -6874 6854 -6846
rect 6882 -6874 7000 -6846
rect 6730 -7006 7000 -6874
rect 6730 -7034 6854 -7006
rect 6882 -7034 7000 -7006
rect 6730 -7166 7000 -7034
rect 6730 -7194 6854 -7166
rect 6882 -7194 7000 -7166
rect 6730 -7326 7000 -7194
rect 6730 -7354 6854 -7326
rect 6882 -7354 7000 -7326
rect 6730 -7486 7000 -7354
rect 6730 -7514 6854 -7486
rect 6882 -7514 7000 -7486
rect 6730 -7646 7000 -7514
rect 6730 -7674 6854 -7646
rect 6882 -7674 7000 -7646
rect 6730 -7806 7000 -7674
rect 6730 -7834 6854 -7806
rect 6882 -7834 7000 -7806
rect 6730 -7966 7000 -7834
rect 6730 -7994 6854 -7966
rect 6882 -7994 7000 -7966
rect 6730 -8126 7000 -7994
rect 6730 -8154 6854 -8126
rect 6882 -8154 7000 -8126
rect 6730 -8286 7000 -8154
rect 6730 -8314 6854 -8286
rect 6882 -8314 7000 -8286
rect 6730 -8446 7000 -8314
rect 6730 -8474 6854 -8446
rect 6882 -8474 7000 -8446
rect 6730 -8606 7000 -8474
rect 6730 -8634 6854 -8606
rect 6882 -8634 7000 -8606
rect 6730 -8766 7000 -8634
rect 6730 -8794 6854 -8766
rect 6882 -8794 7000 -8766
rect 6730 -8926 7000 -8794
rect 6730 -8954 6854 -8926
rect 6882 -8954 7000 -8926
rect 6730 -9086 7000 -8954
rect 6730 -9114 6854 -9086
rect 6882 -9114 7000 -9086
rect 6730 -9230 7000 -9114
rect 3000 -9246 7000 -9230
rect 3000 -9274 3121 -9246
rect 3149 -9274 6854 -9246
rect 6882 -9274 7000 -9246
rect 3000 -9351 7000 -9274
rect 3000 -9379 3306 -9351
rect 3334 -9379 3466 -9351
rect 3494 -9379 3626 -9351
rect 3654 -9379 3786 -9351
rect 3814 -9379 3946 -9351
rect 3974 -9379 4106 -9351
rect 4134 -9379 4266 -9351
rect 4294 -9379 4426 -9351
rect 4454 -9379 4586 -9351
rect 4614 -9379 4746 -9351
rect 4774 -9379 4906 -9351
rect 4934 -9379 5066 -9351
rect 5094 -9379 5226 -9351
rect 5254 -9379 5386 -9351
rect 5414 -9379 5546 -9351
rect 5574 -9379 5706 -9351
rect 5734 -9379 5866 -9351
rect 5894 -9379 6026 -9351
rect 6054 -9379 6186 -9351
rect 6214 -9379 6346 -9351
rect 6374 -9379 6506 -9351
rect 6534 -9379 6666 -9351
rect 6694 -9379 7000 -9351
rect 3000 -9500 7000 -9379
rect 9000 -5726 13000 -5651
rect 9000 -5754 9121 -5726
rect 9149 -5754 12854 -5726
rect 12882 -5754 13000 -5726
rect 9000 -5770 13000 -5754
rect 9000 -5886 9270 -5770
rect 9000 -5914 9121 -5886
rect 9149 -5914 9270 -5886
rect 9000 -6046 9270 -5914
rect 9000 -6074 9121 -6046
rect 9149 -6074 9270 -6046
rect 9000 -6206 9270 -6074
rect 9000 -6234 9121 -6206
rect 9149 -6234 9270 -6206
rect 9000 -6366 9270 -6234
rect 9000 -6394 9121 -6366
rect 9149 -6394 9270 -6366
rect 9000 -6526 9270 -6394
rect 9000 -6554 9121 -6526
rect 9149 -6554 9270 -6526
rect 9000 -6686 9270 -6554
rect 9000 -6714 9121 -6686
rect 9149 -6714 9270 -6686
rect 9000 -6846 9270 -6714
rect 9000 -6874 9121 -6846
rect 9149 -6874 9270 -6846
rect 9000 -7006 9270 -6874
rect 9000 -7034 9121 -7006
rect 9149 -7034 9270 -7006
rect 9000 -7166 9270 -7034
rect 9000 -7194 9121 -7166
rect 9149 -7194 9270 -7166
rect 9000 -7326 9270 -7194
rect 9000 -7354 9121 -7326
rect 9149 -7354 9270 -7326
rect 9000 -7486 9270 -7354
rect 9000 -7514 9121 -7486
rect 9149 -7514 9270 -7486
rect 9000 -7646 9270 -7514
rect 9000 -7674 9121 -7646
rect 9149 -7674 9270 -7646
rect 9000 -7806 9270 -7674
rect 9000 -7834 9121 -7806
rect 9149 -7834 9270 -7806
rect 9000 -7966 9270 -7834
rect 9000 -7994 9121 -7966
rect 9149 -7994 9270 -7966
rect 9000 -8126 9270 -7994
rect 9000 -8154 9121 -8126
rect 9149 -8154 9270 -8126
rect 9000 -8286 9270 -8154
rect 9000 -8314 9121 -8286
rect 9149 -8314 9270 -8286
rect 9000 -8446 9270 -8314
rect 9000 -8474 9121 -8446
rect 9149 -8474 9270 -8446
rect 9000 -8606 9270 -8474
rect 9000 -8634 9121 -8606
rect 9149 -8634 9270 -8606
rect 9000 -8766 9270 -8634
rect 9000 -8794 9121 -8766
rect 9149 -8794 9270 -8766
rect 9000 -8926 9270 -8794
rect 9000 -8954 9121 -8926
rect 9149 -8954 9270 -8926
rect 9000 -9086 9270 -8954
rect 9000 -9114 9121 -9086
rect 9149 -9114 9270 -9086
rect 9000 -9230 9270 -9114
rect 12730 -5886 13000 -5770
rect 12730 -5914 12854 -5886
rect 12882 -5914 13000 -5886
rect 12730 -6046 13000 -5914
rect 12730 -6074 12854 -6046
rect 12882 -6074 13000 -6046
rect 12730 -6206 13000 -6074
rect 12730 -6234 12854 -6206
rect 12882 -6234 13000 -6206
rect 12730 -6366 13000 -6234
rect 12730 -6394 12854 -6366
rect 12882 -6394 13000 -6366
rect 12730 -6526 13000 -6394
rect 12730 -6554 12854 -6526
rect 12882 -6554 13000 -6526
rect 12730 -6686 13000 -6554
rect 12730 -6714 12854 -6686
rect 12882 -6714 13000 -6686
rect 12730 -6846 13000 -6714
rect 12730 -6874 12854 -6846
rect 12882 -6874 13000 -6846
rect 12730 -7006 13000 -6874
rect 12730 -7034 12854 -7006
rect 12882 -7034 13000 -7006
rect 12730 -7166 13000 -7034
rect 12730 -7194 12854 -7166
rect 12882 -7194 13000 -7166
rect 12730 -7326 13000 -7194
rect 12730 -7354 12854 -7326
rect 12882 -7354 13000 -7326
rect 12730 -7486 13000 -7354
rect 12730 -7514 12854 -7486
rect 12882 -7514 13000 -7486
rect 12730 -7646 13000 -7514
rect 12730 -7674 12854 -7646
rect 12882 -7674 13000 -7646
rect 12730 -7806 13000 -7674
rect 12730 -7834 12854 -7806
rect 12882 -7834 13000 -7806
rect 12730 -7966 13000 -7834
rect 12730 -7994 12854 -7966
rect 12882 -7994 13000 -7966
rect 12730 -8126 13000 -7994
rect 12730 -8154 12854 -8126
rect 12882 -8154 13000 -8126
rect 12730 -8286 13000 -8154
rect 12730 -8314 12854 -8286
rect 12882 -8314 13000 -8286
rect 12730 -8446 13000 -8314
rect 12730 -8474 12854 -8446
rect 12882 -8474 13000 -8446
rect 12730 -8606 13000 -8474
rect 12730 -8634 12854 -8606
rect 12882 -8634 13000 -8606
rect 12730 -8766 13000 -8634
rect 12730 -8794 12854 -8766
rect 12882 -8794 13000 -8766
rect 12730 -8926 13000 -8794
rect 12730 -8954 12854 -8926
rect 12882 -8954 13000 -8926
rect 12730 -9086 13000 -8954
rect 12730 -9114 12854 -9086
rect 12882 -9114 13000 -9086
rect 12730 -9230 13000 -9114
rect 9000 -9246 13000 -9230
rect 9000 -9274 9121 -9246
rect 9149 -9274 12854 -9246
rect 12882 -9274 13000 -9246
rect 9000 -9351 13000 -9274
rect 9000 -9379 9306 -9351
rect 9334 -9379 9466 -9351
rect 9494 -9379 9626 -9351
rect 9654 -9379 9786 -9351
rect 9814 -9379 9946 -9351
rect 9974 -9379 10106 -9351
rect 10134 -9379 10266 -9351
rect 10294 -9379 10426 -9351
rect 10454 -9379 10586 -9351
rect 10614 -9379 10746 -9351
rect 10774 -9379 10906 -9351
rect 10934 -9379 11066 -9351
rect 11094 -9379 11226 -9351
rect 11254 -9379 11386 -9351
rect 11414 -9379 11546 -9351
rect 11574 -9379 11706 -9351
rect 11734 -9379 11866 -9351
rect 11894 -9379 12026 -9351
rect 12054 -9379 12186 -9351
rect 12214 -9379 12346 -9351
rect 12374 -9379 12506 -9351
rect 12534 -9379 12666 -9351
rect 12694 -9379 13000 -9351
rect 9000 -9500 13000 -9379
rect 15000 -5623 19000 -5500
rect 15000 -5651 15306 -5623
rect 15334 -5651 15466 -5623
rect 15494 -5651 15626 -5623
rect 15654 -5651 15786 -5623
rect 15814 -5651 15946 -5623
rect 15974 -5651 16106 -5623
rect 16134 -5651 16266 -5623
rect 16294 -5651 16426 -5623
rect 16454 -5651 16586 -5623
rect 16614 -5651 16746 -5623
rect 16774 -5651 16906 -5623
rect 16934 -5651 17066 -5623
rect 17094 -5651 17226 -5623
rect 17254 -5651 17386 -5623
rect 17414 -5651 17546 -5623
rect 17574 -5651 17706 -5623
rect 17734 -5651 17866 -5623
rect 17894 -5651 18026 -5623
rect 18054 -5651 18186 -5623
rect 18214 -5651 18346 -5623
rect 18374 -5651 18506 -5623
rect 18534 -5651 18666 -5623
rect 18694 -5651 19000 -5623
rect 15000 -5726 19000 -5651
rect 15000 -5754 15121 -5726
rect 15149 -5754 18854 -5726
rect 18882 -5754 19000 -5726
rect 15000 -5770 19000 -5754
rect 15000 -5886 15270 -5770
rect 15000 -5914 15121 -5886
rect 15149 -5914 15270 -5886
rect 15000 -6046 15270 -5914
rect 15000 -6074 15121 -6046
rect 15149 -6074 15270 -6046
rect 15000 -6206 15270 -6074
rect 15000 -6234 15121 -6206
rect 15149 -6234 15270 -6206
rect 15000 -6366 15270 -6234
rect 15000 -6394 15121 -6366
rect 15149 -6394 15270 -6366
rect 15000 -6526 15270 -6394
rect 15000 -6554 15121 -6526
rect 15149 -6554 15270 -6526
rect 15000 -6686 15270 -6554
rect 15000 -6714 15121 -6686
rect 15149 -6714 15270 -6686
rect 15000 -6846 15270 -6714
rect 15000 -6874 15121 -6846
rect 15149 -6874 15270 -6846
rect 15000 -7006 15270 -6874
rect 15000 -7034 15121 -7006
rect 15149 -7034 15270 -7006
rect 15000 -7166 15270 -7034
rect 15000 -7194 15121 -7166
rect 15149 -7194 15270 -7166
rect 15000 -7326 15270 -7194
rect 15000 -7354 15121 -7326
rect 15149 -7354 15270 -7326
rect 15000 -7486 15270 -7354
rect 15000 -7514 15121 -7486
rect 15149 -7514 15270 -7486
rect 15000 -7646 15270 -7514
rect 15000 -7674 15121 -7646
rect 15149 -7674 15270 -7646
rect 15000 -7806 15270 -7674
rect 15000 -7834 15121 -7806
rect 15149 -7834 15270 -7806
rect 15000 -7966 15270 -7834
rect 15000 -7994 15121 -7966
rect 15149 -7994 15270 -7966
rect 15000 -8126 15270 -7994
rect 15000 -8154 15121 -8126
rect 15149 -8154 15270 -8126
rect 15000 -8286 15270 -8154
rect 15000 -8314 15121 -8286
rect 15149 -8314 15270 -8286
rect 15000 -8446 15270 -8314
rect 15000 -8474 15121 -8446
rect 15149 -8474 15270 -8446
rect 15000 -8606 15270 -8474
rect 15000 -8634 15121 -8606
rect 15149 -8634 15270 -8606
rect 15000 -8766 15270 -8634
rect 15000 -8794 15121 -8766
rect 15149 -8794 15270 -8766
rect 15000 -8926 15270 -8794
rect 15000 -8954 15121 -8926
rect 15149 -8954 15270 -8926
rect 15000 -9086 15270 -8954
rect 15000 -9114 15121 -9086
rect 15149 -9114 15270 -9086
rect 15000 -9230 15270 -9114
rect 18730 -5886 19000 -5770
rect 18730 -5914 18854 -5886
rect 18882 -5914 19000 -5886
rect 18730 -6046 19000 -5914
rect 18730 -6074 18854 -6046
rect 18882 -6074 19000 -6046
rect 18730 -6206 19000 -6074
rect 18730 -6234 18854 -6206
rect 18882 -6234 19000 -6206
rect 18730 -6366 19000 -6234
rect 18730 -6394 18854 -6366
rect 18882 -6394 19000 -6366
rect 18730 -6526 19000 -6394
rect 18730 -6554 18854 -6526
rect 18882 -6554 19000 -6526
rect 18730 -6686 19000 -6554
rect 18730 -6714 18854 -6686
rect 18882 -6714 19000 -6686
rect 18730 -6846 19000 -6714
rect 18730 -6874 18854 -6846
rect 18882 -6874 19000 -6846
rect 18730 -7006 19000 -6874
rect 18730 -7034 18854 -7006
rect 18882 -7034 19000 -7006
rect 18730 -7166 19000 -7034
rect 18730 -7194 18854 -7166
rect 18882 -7194 19000 -7166
rect 18730 -7326 19000 -7194
rect 18730 -7354 18854 -7326
rect 18882 -7354 19000 -7326
rect 18730 -7486 19000 -7354
rect 18730 -7514 18854 -7486
rect 18882 -7514 19000 -7486
rect 18730 -7646 19000 -7514
rect 18730 -7674 18854 -7646
rect 18882 -7674 19000 -7646
rect 18730 -7806 19000 -7674
rect 18730 -7834 18854 -7806
rect 18882 -7834 19000 -7806
rect 18730 -7966 19000 -7834
rect 18730 -7994 18854 -7966
rect 18882 -7994 19000 -7966
rect 18730 -8126 19000 -7994
rect 18730 -8154 18854 -8126
rect 18882 -8154 19000 -8126
rect 18730 -8286 19000 -8154
rect 18730 -8314 18854 -8286
rect 18882 -8314 19000 -8286
rect 18730 -8446 19000 -8314
rect 18730 -8474 18854 -8446
rect 18882 -8474 19000 -8446
rect 18730 -8606 19000 -8474
rect 18730 -8634 18854 -8606
rect 18882 -8634 19000 -8606
rect 18730 -8766 19000 -8634
rect 18730 -8794 18854 -8766
rect 18882 -8794 19000 -8766
rect 18730 -8926 19000 -8794
rect 18730 -8954 18854 -8926
rect 18882 -8954 19000 -8926
rect 18730 -9086 19000 -8954
rect 18730 -9114 18854 -9086
rect 18882 -9114 19000 -9086
rect 18730 -9230 19000 -9114
rect 15000 -9246 19000 -9230
rect 15000 -9274 15121 -9246
rect 15149 -9274 18854 -9246
rect 18882 -9274 19000 -9246
rect 15000 -9351 19000 -9274
rect 15000 -9379 15306 -9351
rect 15334 -9379 15466 -9351
rect 15494 -9379 15626 -9351
rect 15654 -9379 15786 -9351
rect 15814 -9379 15946 -9351
rect 15974 -9379 16106 -9351
rect 16134 -9379 16266 -9351
rect 16294 -9379 16426 -9351
rect 16454 -9379 16586 -9351
rect 16614 -9379 16746 -9351
rect 16774 -9379 16906 -9351
rect 16934 -9379 17066 -9351
rect 17094 -9379 17226 -9351
rect 17254 -9379 17386 -9351
rect 17414 -9379 17546 -9351
rect 17574 -9379 17706 -9351
rect 17734 -9379 17866 -9351
rect 17894 -9379 18026 -9351
rect 18054 -9379 18186 -9351
rect 18214 -9379 18346 -9351
rect 18374 -9379 18506 -9351
rect 18534 -9379 18666 -9351
rect 18694 -9379 19000 -9351
rect 15000 -9500 19000 -9379
rect 21000 -5623 25000 -5500
rect 21000 -5651 21306 -5623
rect 21334 -5651 21466 -5623
rect 21494 -5651 21626 -5623
rect 21654 -5651 21786 -5623
rect 21814 -5651 21946 -5623
rect 21974 -5651 22106 -5623
rect 22134 -5651 22266 -5623
rect 22294 -5651 22426 -5623
rect 22454 -5651 22586 -5623
rect 22614 -5651 22746 -5623
rect 22774 -5651 22906 -5623
rect 22934 -5651 23066 -5623
rect 23094 -5651 23226 -5623
rect 23254 -5651 23386 -5623
rect 23414 -5651 23546 -5623
rect 23574 -5651 23706 -5623
rect 23734 -5651 23866 -5623
rect 23894 -5651 24026 -5623
rect 24054 -5651 24186 -5623
rect 24214 -5651 24346 -5623
rect 24374 -5651 24506 -5623
rect 24534 -5651 24666 -5623
rect 24694 -5651 25000 -5623
rect 21000 -5726 25000 -5651
rect 21000 -5754 21121 -5726
rect 21149 -5754 24854 -5726
rect 24882 -5754 25000 -5726
rect 21000 -5770 25000 -5754
rect 21000 -5886 21270 -5770
rect 21000 -5914 21121 -5886
rect 21149 -5914 21270 -5886
rect 21000 -6046 21270 -5914
rect 21000 -6074 21121 -6046
rect 21149 -6074 21270 -6046
rect 21000 -6206 21270 -6074
rect 21000 -6234 21121 -6206
rect 21149 -6234 21270 -6206
rect 21000 -6366 21270 -6234
rect 21000 -6394 21121 -6366
rect 21149 -6394 21270 -6366
rect 21000 -6526 21270 -6394
rect 21000 -6554 21121 -6526
rect 21149 -6554 21270 -6526
rect 21000 -6686 21270 -6554
rect 21000 -6714 21121 -6686
rect 21149 -6714 21270 -6686
rect 21000 -6846 21270 -6714
rect 21000 -6874 21121 -6846
rect 21149 -6874 21270 -6846
rect 21000 -7006 21270 -6874
rect 21000 -7034 21121 -7006
rect 21149 -7034 21270 -7006
rect 21000 -7166 21270 -7034
rect 21000 -7194 21121 -7166
rect 21149 -7194 21270 -7166
rect 21000 -7326 21270 -7194
rect 21000 -7354 21121 -7326
rect 21149 -7354 21270 -7326
rect 21000 -7486 21270 -7354
rect 21000 -7514 21121 -7486
rect 21149 -7514 21270 -7486
rect 21000 -7646 21270 -7514
rect 21000 -7674 21121 -7646
rect 21149 -7674 21270 -7646
rect 21000 -7806 21270 -7674
rect 21000 -7834 21121 -7806
rect 21149 -7834 21270 -7806
rect 21000 -7966 21270 -7834
rect 21000 -7994 21121 -7966
rect 21149 -7994 21270 -7966
rect 21000 -8126 21270 -7994
rect 21000 -8154 21121 -8126
rect 21149 -8154 21270 -8126
rect 21000 -8286 21270 -8154
rect 21000 -8314 21121 -8286
rect 21149 -8314 21270 -8286
rect 21000 -8446 21270 -8314
rect 21000 -8474 21121 -8446
rect 21149 -8474 21270 -8446
rect 21000 -8606 21270 -8474
rect 21000 -8634 21121 -8606
rect 21149 -8634 21270 -8606
rect 21000 -8766 21270 -8634
rect 21000 -8794 21121 -8766
rect 21149 -8794 21270 -8766
rect 21000 -8926 21270 -8794
rect 21000 -8954 21121 -8926
rect 21149 -8954 21270 -8926
rect 21000 -9086 21270 -8954
rect 21000 -9114 21121 -9086
rect 21149 -9114 21270 -9086
rect 21000 -9230 21270 -9114
rect 24730 -5886 25000 -5770
rect 24730 -5914 24854 -5886
rect 24882 -5914 25000 -5886
rect 24730 -6046 25000 -5914
rect 24730 -6074 24854 -6046
rect 24882 -6074 25000 -6046
rect 24730 -6206 25000 -6074
rect 24730 -6234 24854 -6206
rect 24882 -6234 25000 -6206
rect 24730 -6366 25000 -6234
rect 24730 -6394 24854 -6366
rect 24882 -6394 25000 -6366
rect 24730 -6526 25000 -6394
rect 24730 -6554 24854 -6526
rect 24882 -6554 25000 -6526
rect 24730 -6686 25000 -6554
rect 24730 -6714 24854 -6686
rect 24882 -6714 25000 -6686
rect 24730 -6846 25000 -6714
rect 24730 -6874 24854 -6846
rect 24882 -6874 25000 -6846
rect 24730 -7006 25000 -6874
rect 24730 -7034 24854 -7006
rect 24882 -7034 25000 -7006
rect 24730 -7166 25000 -7034
rect 24730 -7194 24854 -7166
rect 24882 -7194 25000 -7166
rect 24730 -7326 25000 -7194
rect 24730 -7354 24854 -7326
rect 24882 -7354 25000 -7326
rect 24730 -7486 25000 -7354
rect 24730 -7514 24854 -7486
rect 24882 -7514 25000 -7486
rect 24730 -7646 25000 -7514
rect 24730 -7674 24854 -7646
rect 24882 -7674 25000 -7646
rect 24730 -7806 25000 -7674
rect 24730 -7834 24854 -7806
rect 24882 -7834 25000 -7806
rect 24730 -7966 25000 -7834
rect 24730 -7994 24854 -7966
rect 24882 -7994 25000 -7966
rect 24730 -8126 25000 -7994
rect 24730 -8154 24854 -8126
rect 24882 -8154 25000 -8126
rect 24730 -8286 25000 -8154
rect 24730 -8314 24854 -8286
rect 24882 -8314 25000 -8286
rect 24730 -8446 25000 -8314
rect 24730 -8474 24854 -8446
rect 24882 -8474 25000 -8446
rect 24730 -8606 25000 -8474
rect 24730 -8634 24854 -8606
rect 24882 -8634 25000 -8606
rect 24730 -8766 25000 -8634
rect 24730 -8794 24854 -8766
rect 24882 -8794 25000 -8766
rect 24730 -8926 25000 -8794
rect 24730 -8954 24854 -8926
rect 24882 -8954 25000 -8926
rect 24730 -9086 25000 -8954
rect 24730 -9114 24854 -9086
rect 24882 -9114 25000 -9086
rect 24730 -9230 25000 -9114
rect 21000 -9246 25000 -9230
rect 21000 -9274 21121 -9246
rect 21149 -9274 24854 -9246
rect 24882 -9274 25000 -9246
rect 21000 -9351 25000 -9274
rect 21000 -9379 21306 -9351
rect 21334 -9379 21466 -9351
rect 21494 -9379 21626 -9351
rect 21654 -9379 21786 -9351
rect 21814 -9379 21946 -9351
rect 21974 -9379 22106 -9351
rect 22134 -9379 22266 -9351
rect 22294 -9379 22426 -9351
rect 22454 -9379 22586 -9351
rect 22614 -9379 22746 -9351
rect 22774 -9379 22906 -9351
rect 22934 -9379 23066 -9351
rect 23094 -9379 23226 -9351
rect 23254 -9379 23386 -9351
rect 23414 -9379 23546 -9351
rect 23574 -9379 23706 -9351
rect 23734 -9379 23866 -9351
rect 23894 -9379 24026 -9351
rect 24054 -9379 24186 -9351
rect 24214 -9379 24346 -9351
rect 24374 -9379 24506 -9351
rect 24534 -9379 24666 -9351
rect 24694 -9379 25000 -9351
rect 21000 -9500 25000 -9379
rect 3000 -11623 7000 -11500
rect 3000 -11651 3306 -11623
rect 3334 -11651 3466 -11623
rect 3494 -11651 3626 -11623
rect 3654 -11651 3786 -11623
rect 3814 -11651 3946 -11623
rect 3974 -11651 4106 -11623
rect 4134 -11651 4266 -11623
rect 4294 -11651 4426 -11623
rect 4454 -11651 4586 -11623
rect 4614 -11651 4746 -11623
rect 4774 -11651 4906 -11623
rect 4934 -11651 5066 -11623
rect 5094 -11651 5226 -11623
rect 5254 -11651 5386 -11623
rect 5414 -11651 5546 -11623
rect 5574 -11651 5706 -11623
rect 5734 -11651 5866 -11623
rect 5894 -11651 6026 -11623
rect 6054 -11651 6186 -11623
rect 6214 -11651 6346 -11623
rect 6374 -11651 6506 -11623
rect 6534 -11651 6666 -11623
rect 6694 -11651 7000 -11623
rect 3000 -11726 7000 -11651
rect 3000 -11754 3121 -11726
rect 3149 -11754 6854 -11726
rect 6882 -11754 7000 -11726
rect 3000 -11770 7000 -11754
rect 3000 -11886 3270 -11770
rect 3000 -11914 3121 -11886
rect 3149 -11914 3270 -11886
rect 3000 -12046 3270 -11914
rect 3000 -12074 3121 -12046
rect 3149 -12074 3270 -12046
rect 3000 -12206 3270 -12074
rect 3000 -12234 3121 -12206
rect 3149 -12234 3270 -12206
rect 3000 -12366 3270 -12234
rect 3000 -12394 3121 -12366
rect 3149 -12394 3270 -12366
rect 3000 -12526 3270 -12394
rect 3000 -12554 3121 -12526
rect 3149 -12554 3270 -12526
rect 3000 -12686 3270 -12554
rect 3000 -12714 3121 -12686
rect 3149 -12714 3270 -12686
rect 3000 -12846 3270 -12714
rect 3000 -12874 3121 -12846
rect 3149 -12874 3270 -12846
rect 3000 -13006 3270 -12874
rect 3000 -13034 3121 -13006
rect 3149 -13034 3270 -13006
rect 3000 -13166 3270 -13034
rect 3000 -13194 3121 -13166
rect 3149 -13194 3270 -13166
rect 3000 -13326 3270 -13194
rect 3000 -13354 3121 -13326
rect 3149 -13354 3270 -13326
rect 3000 -13486 3270 -13354
rect 3000 -13514 3121 -13486
rect 3149 -13514 3270 -13486
rect 3000 -13646 3270 -13514
rect 3000 -13674 3121 -13646
rect 3149 -13674 3270 -13646
rect 3000 -13806 3270 -13674
rect 3000 -13834 3121 -13806
rect 3149 -13834 3270 -13806
rect 3000 -13966 3270 -13834
rect 3000 -13994 3121 -13966
rect 3149 -13994 3270 -13966
rect 3000 -14126 3270 -13994
rect 3000 -14154 3121 -14126
rect 3149 -14154 3270 -14126
rect 3000 -14286 3270 -14154
rect 3000 -14314 3121 -14286
rect 3149 -14314 3270 -14286
rect 3000 -14446 3270 -14314
rect 3000 -14474 3121 -14446
rect 3149 -14474 3270 -14446
rect 3000 -14606 3270 -14474
rect 3000 -14634 3121 -14606
rect 3149 -14634 3270 -14606
rect 3000 -14766 3270 -14634
rect 3000 -14794 3121 -14766
rect 3149 -14794 3270 -14766
rect 3000 -14926 3270 -14794
rect 3000 -14954 3121 -14926
rect 3149 -14954 3270 -14926
rect 3000 -15086 3270 -14954
rect 3000 -15114 3121 -15086
rect 3149 -15114 3270 -15086
rect 3000 -15230 3270 -15114
rect 6730 -11886 7000 -11770
rect 6730 -11914 6854 -11886
rect 6882 -11914 7000 -11886
rect 6730 -12046 7000 -11914
rect 6730 -12074 6854 -12046
rect 6882 -12074 7000 -12046
rect 6730 -12206 7000 -12074
rect 6730 -12234 6854 -12206
rect 6882 -12234 7000 -12206
rect 6730 -12366 7000 -12234
rect 6730 -12394 6854 -12366
rect 6882 -12394 7000 -12366
rect 6730 -12526 7000 -12394
rect 6730 -12554 6854 -12526
rect 6882 -12554 7000 -12526
rect 6730 -12686 7000 -12554
rect 6730 -12714 6854 -12686
rect 6882 -12714 7000 -12686
rect 6730 -12846 7000 -12714
rect 6730 -12874 6854 -12846
rect 6882 -12874 7000 -12846
rect 6730 -13006 7000 -12874
rect 6730 -13034 6854 -13006
rect 6882 -13034 7000 -13006
rect 6730 -13166 7000 -13034
rect 6730 -13194 6854 -13166
rect 6882 -13194 7000 -13166
rect 6730 -13326 7000 -13194
rect 6730 -13354 6854 -13326
rect 6882 -13354 7000 -13326
rect 6730 -13486 7000 -13354
rect 6730 -13514 6854 -13486
rect 6882 -13514 7000 -13486
rect 6730 -13646 7000 -13514
rect 6730 -13674 6854 -13646
rect 6882 -13674 7000 -13646
rect 6730 -13806 7000 -13674
rect 6730 -13834 6854 -13806
rect 6882 -13834 7000 -13806
rect 6730 -13966 7000 -13834
rect 6730 -13994 6854 -13966
rect 6882 -13994 7000 -13966
rect 6730 -14126 7000 -13994
rect 6730 -14154 6854 -14126
rect 6882 -14154 7000 -14126
rect 6730 -14286 7000 -14154
rect 6730 -14314 6854 -14286
rect 6882 -14314 7000 -14286
rect 6730 -14446 7000 -14314
rect 6730 -14474 6854 -14446
rect 6882 -14474 7000 -14446
rect 6730 -14606 7000 -14474
rect 6730 -14634 6854 -14606
rect 6882 -14634 7000 -14606
rect 6730 -14766 7000 -14634
rect 6730 -14794 6854 -14766
rect 6882 -14794 7000 -14766
rect 6730 -14926 7000 -14794
rect 6730 -14954 6854 -14926
rect 6882 -14954 7000 -14926
rect 6730 -15086 7000 -14954
rect 6730 -15114 6854 -15086
rect 6882 -15114 7000 -15086
rect 6730 -15230 7000 -15114
rect 3000 -15246 7000 -15230
rect 3000 -15274 3121 -15246
rect 3149 -15274 6854 -15246
rect 6882 -15274 7000 -15246
rect 3000 -15351 7000 -15274
rect 3000 -15379 3306 -15351
rect 3334 -15379 3466 -15351
rect 3494 -15379 3626 -15351
rect 3654 -15379 3786 -15351
rect 3814 -15379 3946 -15351
rect 3974 -15379 4106 -15351
rect 4134 -15379 4266 -15351
rect 4294 -15379 4426 -15351
rect 4454 -15379 4586 -15351
rect 4614 -15379 4746 -15351
rect 4774 -15379 4906 -15351
rect 4934 -15379 5066 -15351
rect 5094 -15379 5226 -15351
rect 5254 -15379 5386 -15351
rect 5414 -15379 5546 -15351
rect 5574 -15379 5706 -15351
rect 5734 -15379 5866 -15351
rect 5894 -15379 6026 -15351
rect 6054 -15379 6186 -15351
rect 6214 -15379 6346 -15351
rect 6374 -15379 6506 -15351
rect 6534 -15379 6666 -15351
rect 6694 -15379 7000 -15351
rect 3000 -15500 7000 -15379
rect 9000 -11623 13000 -11500
rect 9000 -11651 9306 -11623
rect 9334 -11651 9466 -11623
rect 9494 -11651 9626 -11623
rect 9654 -11651 9786 -11623
rect 9814 -11651 9946 -11623
rect 9974 -11651 10106 -11623
rect 10134 -11651 10266 -11623
rect 10294 -11651 10426 -11623
rect 10454 -11651 10586 -11623
rect 10614 -11651 10746 -11623
rect 10774 -11651 10906 -11623
rect 10934 -11651 11066 -11623
rect 11094 -11651 11226 -11623
rect 11254 -11651 11386 -11623
rect 11414 -11651 11546 -11623
rect 11574 -11651 11706 -11623
rect 11734 -11651 11866 -11623
rect 11894 -11651 12026 -11623
rect 12054 -11651 12186 -11623
rect 12214 -11651 12346 -11623
rect 12374 -11651 12506 -11623
rect 12534 -11651 12666 -11623
rect 12694 -11651 13000 -11623
rect 9000 -11726 13000 -11651
rect 9000 -11754 9121 -11726
rect 9149 -11754 12854 -11726
rect 12882 -11754 13000 -11726
rect 9000 -11770 13000 -11754
rect 9000 -11886 9270 -11770
rect 9000 -11914 9121 -11886
rect 9149 -11914 9270 -11886
rect 9000 -12046 9270 -11914
rect 9000 -12074 9121 -12046
rect 9149 -12074 9270 -12046
rect 9000 -12206 9270 -12074
rect 9000 -12234 9121 -12206
rect 9149 -12234 9270 -12206
rect 9000 -12366 9270 -12234
rect 9000 -12394 9121 -12366
rect 9149 -12394 9270 -12366
rect 9000 -12526 9270 -12394
rect 9000 -12554 9121 -12526
rect 9149 -12554 9270 -12526
rect 9000 -12686 9270 -12554
rect 9000 -12714 9121 -12686
rect 9149 -12714 9270 -12686
rect 9000 -12846 9270 -12714
rect 9000 -12874 9121 -12846
rect 9149 -12874 9270 -12846
rect 9000 -13006 9270 -12874
rect 9000 -13034 9121 -13006
rect 9149 -13034 9270 -13006
rect 9000 -13166 9270 -13034
rect 9000 -13194 9121 -13166
rect 9149 -13194 9270 -13166
rect 9000 -13326 9270 -13194
rect 9000 -13354 9121 -13326
rect 9149 -13354 9270 -13326
rect 9000 -13486 9270 -13354
rect 9000 -13514 9121 -13486
rect 9149 -13514 9270 -13486
rect 9000 -13646 9270 -13514
rect 9000 -13674 9121 -13646
rect 9149 -13674 9270 -13646
rect 9000 -13806 9270 -13674
rect 9000 -13834 9121 -13806
rect 9149 -13834 9270 -13806
rect 9000 -13966 9270 -13834
rect 9000 -13994 9121 -13966
rect 9149 -13994 9270 -13966
rect 9000 -14126 9270 -13994
rect 9000 -14154 9121 -14126
rect 9149 -14154 9270 -14126
rect 9000 -14286 9270 -14154
rect 9000 -14314 9121 -14286
rect 9149 -14314 9270 -14286
rect 9000 -14446 9270 -14314
rect 9000 -14474 9121 -14446
rect 9149 -14474 9270 -14446
rect 9000 -14606 9270 -14474
rect 9000 -14634 9121 -14606
rect 9149 -14634 9270 -14606
rect 9000 -14766 9270 -14634
rect 9000 -14794 9121 -14766
rect 9149 -14794 9270 -14766
rect 9000 -14926 9270 -14794
rect 9000 -14954 9121 -14926
rect 9149 -14954 9270 -14926
rect 9000 -15086 9270 -14954
rect 9000 -15114 9121 -15086
rect 9149 -15114 9270 -15086
rect 9000 -15230 9270 -15114
rect 12730 -11886 13000 -11770
rect 12730 -11914 12854 -11886
rect 12882 -11914 13000 -11886
rect 12730 -12046 13000 -11914
rect 12730 -12074 12854 -12046
rect 12882 -12074 13000 -12046
rect 12730 -12206 13000 -12074
rect 12730 -12234 12854 -12206
rect 12882 -12234 13000 -12206
rect 12730 -12366 13000 -12234
rect 12730 -12394 12854 -12366
rect 12882 -12394 13000 -12366
rect 12730 -12526 13000 -12394
rect 12730 -12554 12854 -12526
rect 12882 -12554 13000 -12526
rect 12730 -12686 13000 -12554
rect 12730 -12714 12854 -12686
rect 12882 -12714 13000 -12686
rect 12730 -12846 13000 -12714
rect 12730 -12874 12854 -12846
rect 12882 -12874 13000 -12846
rect 12730 -13006 13000 -12874
rect 12730 -13034 12854 -13006
rect 12882 -13034 13000 -13006
rect 12730 -13166 13000 -13034
rect 12730 -13194 12854 -13166
rect 12882 -13194 13000 -13166
rect 12730 -13326 13000 -13194
rect 12730 -13354 12854 -13326
rect 12882 -13354 13000 -13326
rect 12730 -13486 13000 -13354
rect 12730 -13514 12854 -13486
rect 12882 -13514 13000 -13486
rect 12730 -13646 13000 -13514
rect 12730 -13674 12854 -13646
rect 12882 -13674 13000 -13646
rect 12730 -13806 13000 -13674
rect 12730 -13834 12854 -13806
rect 12882 -13834 13000 -13806
rect 12730 -13966 13000 -13834
rect 12730 -13994 12854 -13966
rect 12882 -13994 13000 -13966
rect 12730 -14126 13000 -13994
rect 12730 -14154 12854 -14126
rect 12882 -14154 13000 -14126
rect 12730 -14286 13000 -14154
rect 12730 -14314 12854 -14286
rect 12882 -14314 13000 -14286
rect 12730 -14446 13000 -14314
rect 12730 -14474 12854 -14446
rect 12882 -14474 13000 -14446
rect 12730 -14606 13000 -14474
rect 12730 -14634 12854 -14606
rect 12882 -14634 13000 -14606
rect 12730 -14766 13000 -14634
rect 12730 -14794 12854 -14766
rect 12882 -14794 13000 -14766
rect 12730 -14926 13000 -14794
rect 12730 -14954 12854 -14926
rect 12882 -14954 13000 -14926
rect 12730 -15086 13000 -14954
rect 12730 -15114 12854 -15086
rect 12882 -15114 13000 -15086
rect 12730 -15230 13000 -15114
rect 9000 -15246 13000 -15230
rect 9000 -15274 9121 -15246
rect 9149 -15274 12854 -15246
rect 12882 -15274 13000 -15246
rect 9000 -15351 13000 -15274
rect 9000 -15379 9306 -15351
rect 9334 -15379 9466 -15351
rect 9494 -15379 9626 -15351
rect 9654 -15379 9786 -15351
rect 9814 -15379 9946 -15351
rect 9974 -15379 10106 -15351
rect 10134 -15379 10266 -15351
rect 10294 -15379 10426 -15351
rect 10454 -15379 10586 -15351
rect 10614 -15379 10746 -15351
rect 10774 -15379 10906 -15351
rect 10934 -15379 11066 -15351
rect 11094 -15379 11226 -15351
rect 11254 -15379 11386 -15351
rect 11414 -15379 11546 -15351
rect 11574 -15379 11706 -15351
rect 11734 -15379 11866 -15351
rect 11894 -15379 12026 -15351
rect 12054 -15379 12186 -15351
rect 12214 -15379 12346 -15351
rect 12374 -15379 12506 -15351
rect 12534 -15379 12666 -15351
rect 12694 -15379 13000 -15351
rect 9000 -15500 13000 -15379
rect 15000 -11623 19000 -11500
rect 15000 -11651 15306 -11623
rect 15334 -11651 15466 -11623
rect 15494 -11651 15626 -11623
rect 15654 -11651 15786 -11623
rect 15814 -11651 15946 -11623
rect 15974 -11651 16106 -11623
rect 16134 -11651 16266 -11623
rect 16294 -11651 16426 -11623
rect 16454 -11651 16586 -11623
rect 16614 -11651 16746 -11623
rect 16774 -11651 16906 -11623
rect 16934 -11651 17066 -11623
rect 17094 -11651 17226 -11623
rect 17254 -11651 17386 -11623
rect 17414 -11651 17546 -11623
rect 17574 -11651 17706 -11623
rect 17734 -11651 17866 -11623
rect 17894 -11651 18026 -11623
rect 18054 -11651 18186 -11623
rect 18214 -11651 18346 -11623
rect 18374 -11651 18506 -11623
rect 18534 -11651 18666 -11623
rect 18694 -11651 19000 -11623
rect 15000 -11726 19000 -11651
rect 15000 -11754 15121 -11726
rect 15149 -11754 18854 -11726
rect 18882 -11754 19000 -11726
rect 15000 -11770 19000 -11754
rect 15000 -11886 15270 -11770
rect 15000 -11914 15121 -11886
rect 15149 -11914 15270 -11886
rect 15000 -12046 15270 -11914
rect 15000 -12074 15121 -12046
rect 15149 -12074 15270 -12046
rect 15000 -12206 15270 -12074
rect 15000 -12234 15121 -12206
rect 15149 -12234 15270 -12206
rect 15000 -12366 15270 -12234
rect 15000 -12394 15121 -12366
rect 15149 -12394 15270 -12366
rect 15000 -12526 15270 -12394
rect 15000 -12554 15121 -12526
rect 15149 -12554 15270 -12526
rect 15000 -12686 15270 -12554
rect 15000 -12714 15121 -12686
rect 15149 -12714 15270 -12686
rect 15000 -12846 15270 -12714
rect 15000 -12874 15121 -12846
rect 15149 -12874 15270 -12846
rect 15000 -13006 15270 -12874
rect 15000 -13034 15121 -13006
rect 15149 -13034 15270 -13006
rect 15000 -13166 15270 -13034
rect 15000 -13194 15121 -13166
rect 15149 -13194 15270 -13166
rect 15000 -13326 15270 -13194
rect 15000 -13354 15121 -13326
rect 15149 -13354 15270 -13326
rect 15000 -13486 15270 -13354
rect 15000 -13514 15121 -13486
rect 15149 -13514 15270 -13486
rect 15000 -13646 15270 -13514
rect 15000 -13674 15121 -13646
rect 15149 -13674 15270 -13646
rect 15000 -13806 15270 -13674
rect 15000 -13834 15121 -13806
rect 15149 -13834 15270 -13806
rect 15000 -13966 15270 -13834
rect 15000 -13994 15121 -13966
rect 15149 -13994 15270 -13966
rect 15000 -14126 15270 -13994
rect 15000 -14154 15121 -14126
rect 15149 -14154 15270 -14126
rect 15000 -14286 15270 -14154
rect 15000 -14314 15121 -14286
rect 15149 -14314 15270 -14286
rect 15000 -14446 15270 -14314
rect 15000 -14474 15121 -14446
rect 15149 -14474 15270 -14446
rect 15000 -14606 15270 -14474
rect 15000 -14634 15121 -14606
rect 15149 -14634 15270 -14606
rect 15000 -14766 15270 -14634
rect 15000 -14794 15121 -14766
rect 15149 -14794 15270 -14766
rect 15000 -14926 15270 -14794
rect 15000 -14954 15121 -14926
rect 15149 -14954 15270 -14926
rect 15000 -15086 15270 -14954
rect 15000 -15114 15121 -15086
rect 15149 -15114 15270 -15086
rect 15000 -15230 15270 -15114
rect 18730 -11886 19000 -11770
rect 18730 -11914 18854 -11886
rect 18882 -11914 19000 -11886
rect 18730 -12046 19000 -11914
rect 18730 -12074 18854 -12046
rect 18882 -12074 19000 -12046
rect 18730 -12206 19000 -12074
rect 18730 -12234 18854 -12206
rect 18882 -12234 19000 -12206
rect 18730 -12366 19000 -12234
rect 18730 -12394 18854 -12366
rect 18882 -12394 19000 -12366
rect 18730 -12526 19000 -12394
rect 18730 -12554 18854 -12526
rect 18882 -12554 19000 -12526
rect 18730 -12686 19000 -12554
rect 18730 -12714 18854 -12686
rect 18882 -12714 19000 -12686
rect 18730 -12846 19000 -12714
rect 18730 -12874 18854 -12846
rect 18882 -12874 19000 -12846
rect 18730 -13006 19000 -12874
rect 18730 -13034 18854 -13006
rect 18882 -13034 19000 -13006
rect 18730 -13166 19000 -13034
rect 18730 -13194 18854 -13166
rect 18882 -13194 19000 -13166
rect 18730 -13326 19000 -13194
rect 18730 -13354 18854 -13326
rect 18882 -13354 19000 -13326
rect 18730 -13486 19000 -13354
rect 18730 -13514 18854 -13486
rect 18882 -13514 19000 -13486
rect 18730 -13646 19000 -13514
rect 18730 -13674 18854 -13646
rect 18882 -13674 19000 -13646
rect 18730 -13806 19000 -13674
rect 18730 -13834 18854 -13806
rect 18882 -13834 19000 -13806
rect 18730 -13966 19000 -13834
rect 18730 -13994 18854 -13966
rect 18882 -13994 19000 -13966
rect 18730 -14126 19000 -13994
rect 18730 -14154 18854 -14126
rect 18882 -14154 19000 -14126
rect 18730 -14286 19000 -14154
rect 18730 -14314 18854 -14286
rect 18882 -14314 19000 -14286
rect 18730 -14446 19000 -14314
rect 18730 -14474 18854 -14446
rect 18882 -14474 19000 -14446
rect 18730 -14606 19000 -14474
rect 18730 -14634 18854 -14606
rect 18882 -14634 19000 -14606
rect 18730 -14766 19000 -14634
rect 18730 -14794 18854 -14766
rect 18882 -14794 19000 -14766
rect 18730 -14926 19000 -14794
rect 18730 -14954 18854 -14926
rect 18882 -14954 19000 -14926
rect 18730 -15086 19000 -14954
rect 18730 -15114 18854 -15086
rect 18882 -15114 19000 -15086
rect 18730 -15230 19000 -15114
rect 15000 -15246 19000 -15230
rect 15000 -15274 15121 -15246
rect 15149 -15274 18854 -15246
rect 18882 -15274 19000 -15246
rect 15000 -15351 19000 -15274
rect 15000 -15379 15306 -15351
rect 15334 -15379 15466 -15351
rect 15494 -15379 15626 -15351
rect 15654 -15379 15786 -15351
rect 15814 -15379 15946 -15351
rect 15974 -15379 16106 -15351
rect 16134 -15379 16266 -15351
rect 16294 -15379 16426 -15351
rect 16454 -15379 16586 -15351
rect 16614 -15379 16746 -15351
rect 16774 -15379 16906 -15351
rect 16934 -15379 17066 -15351
rect 17094 -15379 17226 -15351
rect 17254 -15379 17386 -15351
rect 17414 -15379 17546 -15351
rect 17574 -15379 17706 -15351
rect 17734 -15379 17866 -15351
rect 17894 -15379 18026 -15351
rect 18054 -15379 18186 -15351
rect 18214 -15379 18346 -15351
rect 18374 -15379 18506 -15351
rect 18534 -15379 18666 -15351
rect 18694 -15379 19000 -15351
rect 15000 -15500 19000 -15379
rect 21000 -11623 25000 -11500
rect 21000 -11651 21306 -11623
rect 21334 -11651 21466 -11623
rect 21494 -11651 21626 -11623
rect 21654 -11651 21786 -11623
rect 21814 -11651 21946 -11623
rect 21974 -11651 22106 -11623
rect 22134 -11651 22266 -11623
rect 22294 -11651 22426 -11623
rect 22454 -11651 22586 -11623
rect 22614 -11651 22746 -11623
rect 22774 -11651 22906 -11623
rect 22934 -11651 23066 -11623
rect 23094 -11651 23226 -11623
rect 23254 -11651 23386 -11623
rect 23414 -11651 23546 -11623
rect 23574 -11651 23706 -11623
rect 23734 -11651 23866 -11623
rect 23894 -11651 24026 -11623
rect 24054 -11651 24186 -11623
rect 24214 -11651 24346 -11623
rect 24374 -11651 24506 -11623
rect 24534 -11651 24666 -11623
rect 24694 -11651 25000 -11623
rect 21000 -11726 25000 -11651
rect 21000 -11754 21121 -11726
rect 21149 -11754 24854 -11726
rect 24882 -11754 25000 -11726
rect 21000 -11770 25000 -11754
rect 21000 -11886 21270 -11770
rect 21000 -11914 21121 -11886
rect 21149 -11914 21270 -11886
rect 21000 -12046 21270 -11914
rect 21000 -12074 21121 -12046
rect 21149 -12074 21270 -12046
rect 21000 -12206 21270 -12074
rect 21000 -12234 21121 -12206
rect 21149 -12234 21270 -12206
rect 21000 -12366 21270 -12234
rect 21000 -12394 21121 -12366
rect 21149 -12394 21270 -12366
rect 21000 -12526 21270 -12394
rect 21000 -12554 21121 -12526
rect 21149 -12554 21270 -12526
rect 21000 -12686 21270 -12554
rect 21000 -12714 21121 -12686
rect 21149 -12714 21270 -12686
rect 21000 -12846 21270 -12714
rect 21000 -12874 21121 -12846
rect 21149 -12874 21270 -12846
rect 21000 -13006 21270 -12874
rect 21000 -13034 21121 -13006
rect 21149 -13034 21270 -13006
rect 21000 -13166 21270 -13034
rect 21000 -13194 21121 -13166
rect 21149 -13194 21270 -13166
rect 21000 -13326 21270 -13194
rect 21000 -13354 21121 -13326
rect 21149 -13354 21270 -13326
rect 21000 -13486 21270 -13354
rect 21000 -13514 21121 -13486
rect 21149 -13514 21270 -13486
rect 21000 -13646 21270 -13514
rect 21000 -13674 21121 -13646
rect 21149 -13674 21270 -13646
rect 21000 -13806 21270 -13674
rect 21000 -13834 21121 -13806
rect 21149 -13834 21270 -13806
rect 21000 -13966 21270 -13834
rect 21000 -13994 21121 -13966
rect 21149 -13994 21270 -13966
rect 21000 -14126 21270 -13994
rect 21000 -14154 21121 -14126
rect 21149 -14154 21270 -14126
rect 21000 -14286 21270 -14154
rect 21000 -14314 21121 -14286
rect 21149 -14314 21270 -14286
rect 21000 -14446 21270 -14314
rect 21000 -14474 21121 -14446
rect 21149 -14474 21270 -14446
rect 21000 -14606 21270 -14474
rect 21000 -14634 21121 -14606
rect 21149 -14634 21270 -14606
rect 21000 -14766 21270 -14634
rect 21000 -14794 21121 -14766
rect 21149 -14794 21270 -14766
rect 21000 -14926 21270 -14794
rect 21000 -14954 21121 -14926
rect 21149 -14954 21270 -14926
rect 21000 -15086 21270 -14954
rect 21000 -15114 21121 -15086
rect 21149 -15114 21270 -15086
rect 21000 -15230 21270 -15114
rect 24730 -11886 25000 -11770
rect 24730 -11914 24854 -11886
rect 24882 -11914 25000 -11886
rect 24730 -12046 25000 -11914
rect 24730 -12074 24854 -12046
rect 24882 -12074 25000 -12046
rect 24730 -12206 25000 -12074
rect 24730 -12234 24854 -12206
rect 24882 -12234 25000 -12206
rect 24730 -12366 25000 -12234
rect 24730 -12394 24854 -12366
rect 24882 -12394 25000 -12366
rect 24730 -12526 25000 -12394
rect 24730 -12554 24854 -12526
rect 24882 -12554 25000 -12526
rect 24730 -12686 25000 -12554
rect 24730 -12714 24854 -12686
rect 24882 -12714 25000 -12686
rect 24730 -12846 25000 -12714
rect 24730 -12874 24854 -12846
rect 24882 -12874 25000 -12846
rect 24730 -13006 25000 -12874
rect 24730 -13034 24854 -13006
rect 24882 -13034 25000 -13006
rect 24730 -13166 25000 -13034
rect 24730 -13194 24854 -13166
rect 24882 -13194 25000 -13166
rect 24730 -13326 25000 -13194
rect 24730 -13354 24854 -13326
rect 24882 -13354 25000 -13326
rect 24730 -13486 25000 -13354
rect 24730 -13514 24854 -13486
rect 24882 -13514 25000 -13486
rect 24730 -13646 25000 -13514
rect 24730 -13674 24854 -13646
rect 24882 -13674 25000 -13646
rect 24730 -13806 25000 -13674
rect 24730 -13834 24854 -13806
rect 24882 -13834 25000 -13806
rect 24730 -13966 25000 -13834
rect 24730 -13994 24854 -13966
rect 24882 -13994 25000 -13966
rect 24730 -14126 25000 -13994
rect 24730 -14154 24854 -14126
rect 24882 -14154 25000 -14126
rect 24730 -14286 25000 -14154
rect 24730 -14314 24854 -14286
rect 24882 -14314 25000 -14286
rect 24730 -14446 25000 -14314
rect 24730 -14474 24854 -14446
rect 24882 -14474 25000 -14446
rect 24730 -14606 25000 -14474
rect 24730 -14634 24854 -14606
rect 24882 -14634 25000 -14606
rect 24730 -14766 25000 -14634
rect 24730 -14794 24854 -14766
rect 24882 -14794 25000 -14766
rect 24730 -14926 25000 -14794
rect 24730 -14954 24854 -14926
rect 24882 -14954 25000 -14926
rect 24730 -15086 25000 -14954
rect 24730 -15114 24854 -15086
rect 24882 -15114 25000 -15086
rect 24730 -15230 25000 -15114
rect 21000 -15246 25000 -15230
rect 21000 -15274 21121 -15246
rect 21149 -15274 24854 -15246
rect 24882 -15274 25000 -15246
rect 21000 -15351 25000 -15274
rect 21000 -15379 21306 -15351
rect 21334 -15379 21466 -15351
rect 21494 -15379 21626 -15351
rect 21654 -15379 21786 -15351
rect 21814 -15379 21946 -15351
rect 21974 -15379 22106 -15351
rect 22134 -15379 22266 -15351
rect 22294 -15379 22426 -15351
rect 22454 -15379 22586 -15351
rect 22614 -15379 22746 -15351
rect 22774 -15379 22906 -15351
rect 22934 -15379 23066 -15351
rect 23094 -15379 23226 -15351
rect 23254 -15379 23386 -15351
rect 23414 -15379 23546 -15351
rect 23574 -15379 23706 -15351
rect 23734 -15379 23866 -15351
rect 23894 -15379 24026 -15351
rect 24054 -15379 24186 -15351
rect 24214 -15379 24346 -15351
rect 24374 -15379 24506 -15351
rect 24534 -15379 24666 -15351
rect 24694 -15379 25000 -15351
rect 21000 -15500 25000 -15379
<< via2 >>
rect 3306 9378 3334 9379
rect 3306 9352 3307 9378
rect 3307 9352 3333 9378
rect 3333 9352 3334 9378
rect 3306 9351 3334 9352
rect 3466 9378 3494 9379
rect 3466 9352 3467 9378
rect 3467 9352 3493 9378
rect 3493 9352 3494 9378
rect 3466 9351 3494 9352
rect 3626 9378 3654 9379
rect 3626 9352 3627 9378
rect 3627 9352 3653 9378
rect 3653 9352 3654 9378
rect 3626 9351 3654 9352
rect 3786 9378 3814 9379
rect 3786 9352 3787 9378
rect 3787 9352 3813 9378
rect 3813 9352 3814 9378
rect 3786 9351 3814 9352
rect 3946 9378 3974 9379
rect 3946 9352 3947 9378
rect 3947 9352 3973 9378
rect 3973 9352 3974 9378
rect 3946 9351 3974 9352
rect 4106 9378 4134 9379
rect 4106 9352 4107 9378
rect 4107 9352 4133 9378
rect 4133 9352 4134 9378
rect 4106 9351 4134 9352
rect 4266 9378 4294 9379
rect 4266 9352 4267 9378
rect 4267 9352 4293 9378
rect 4293 9352 4294 9378
rect 4266 9351 4294 9352
rect 4426 9378 4454 9379
rect 4426 9352 4427 9378
rect 4427 9352 4453 9378
rect 4453 9352 4454 9378
rect 4426 9351 4454 9352
rect 4586 9378 4614 9379
rect 4586 9352 4587 9378
rect 4587 9352 4613 9378
rect 4613 9352 4614 9378
rect 4586 9351 4614 9352
rect 4746 9378 4774 9379
rect 4746 9352 4747 9378
rect 4747 9352 4773 9378
rect 4773 9352 4774 9378
rect 4746 9351 4774 9352
rect 4906 9378 4934 9379
rect 4906 9352 4907 9378
rect 4907 9352 4933 9378
rect 4933 9352 4934 9378
rect 4906 9351 4934 9352
rect 5066 9378 5094 9379
rect 5066 9352 5067 9378
rect 5067 9352 5093 9378
rect 5093 9352 5094 9378
rect 5066 9351 5094 9352
rect 5226 9378 5254 9379
rect 5226 9352 5227 9378
rect 5227 9352 5253 9378
rect 5253 9352 5254 9378
rect 5226 9351 5254 9352
rect 5386 9378 5414 9379
rect 5386 9352 5387 9378
rect 5387 9352 5413 9378
rect 5413 9352 5414 9378
rect 5386 9351 5414 9352
rect 5546 9378 5574 9379
rect 5546 9352 5547 9378
rect 5547 9352 5573 9378
rect 5573 9352 5574 9378
rect 5546 9351 5574 9352
rect 5706 9378 5734 9379
rect 5706 9352 5707 9378
rect 5707 9352 5733 9378
rect 5733 9352 5734 9378
rect 5706 9351 5734 9352
rect 5866 9378 5894 9379
rect 5866 9352 5867 9378
rect 5867 9352 5893 9378
rect 5893 9352 5894 9378
rect 5866 9351 5894 9352
rect 6026 9378 6054 9379
rect 6026 9352 6027 9378
rect 6027 9352 6053 9378
rect 6053 9352 6054 9378
rect 6026 9351 6054 9352
rect 6186 9378 6214 9379
rect 6186 9352 6187 9378
rect 6187 9352 6213 9378
rect 6213 9352 6214 9378
rect 6186 9351 6214 9352
rect 6346 9378 6374 9379
rect 6346 9352 6347 9378
rect 6347 9352 6373 9378
rect 6373 9352 6374 9378
rect 6346 9351 6374 9352
rect 6506 9378 6534 9379
rect 6506 9352 6507 9378
rect 6507 9352 6533 9378
rect 6533 9352 6534 9378
rect 6506 9351 6534 9352
rect 6666 9378 6694 9379
rect 6666 9352 6667 9378
rect 6667 9352 6693 9378
rect 6693 9352 6694 9378
rect 6666 9351 6694 9352
rect 3118 9273 3146 9274
rect 3118 9247 3119 9273
rect 3119 9247 3145 9273
rect 3145 9247 3146 9273
rect 3118 9246 3146 9247
rect 6851 9273 6879 9274
rect 6851 9247 6852 9273
rect 6852 9247 6878 9273
rect 6878 9247 6879 9273
rect 6851 9246 6879 9247
rect 3118 9113 3146 9114
rect 3118 9087 3119 9113
rect 3119 9087 3145 9113
rect 3145 9087 3146 9113
rect 3118 9086 3146 9087
rect 3118 8953 3146 8954
rect 3118 8927 3119 8953
rect 3119 8927 3145 8953
rect 3145 8927 3146 8953
rect 3118 8926 3146 8927
rect 3118 8793 3146 8794
rect 3118 8767 3119 8793
rect 3119 8767 3145 8793
rect 3145 8767 3146 8793
rect 3118 8766 3146 8767
rect 3118 8633 3146 8634
rect 3118 8607 3119 8633
rect 3119 8607 3145 8633
rect 3145 8607 3146 8633
rect 3118 8606 3146 8607
rect 3118 8473 3146 8474
rect 3118 8447 3119 8473
rect 3119 8447 3145 8473
rect 3145 8447 3146 8473
rect 3118 8446 3146 8447
rect 3118 8313 3146 8314
rect 3118 8287 3119 8313
rect 3119 8287 3145 8313
rect 3145 8287 3146 8313
rect 3118 8286 3146 8287
rect 3118 8153 3146 8154
rect 3118 8127 3119 8153
rect 3119 8127 3145 8153
rect 3145 8127 3146 8153
rect 3118 8126 3146 8127
rect 3118 7993 3146 7994
rect 3118 7967 3119 7993
rect 3119 7967 3145 7993
rect 3145 7967 3146 7993
rect 3118 7966 3146 7967
rect 3118 7833 3146 7834
rect 3118 7807 3119 7833
rect 3119 7807 3145 7833
rect 3145 7807 3146 7833
rect 3118 7806 3146 7807
rect 3118 7673 3146 7674
rect 3118 7647 3119 7673
rect 3119 7647 3145 7673
rect 3145 7647 3146 7673
rect 3118 7646 3146 7647
rect 3118 7513 3146 7514
rect 3118 7487 3119 7513
rect 3119 7487 3145 7513
rect 3145 7487 3146 7513
rect 3118 7486 3146 7487
rect 3118 7353 3146 7354
rect 3118 7327 3119 7353
rect 3119 7327 3145 7353
rect 3145 7327 3146 7353
rect 3118 7326 3146 7327
rect 3118 7193 3146 7194
rect 3118 7167 3119 7193
rect 3119 7167 3145 7193
rect 3145 7167 3146 7193
rect 3118 7166 3146 7167
rect 3118 7033 3146 7034
rect 3118 7007 3119 7033
rect 3119 7007 3145 7033
rect 3145 7007 3146 7033
rect 3118 7006 3146 7007
rect 3118 6873 3146 6874
rect 3118 6847 3119 6873
rect 3119 6847 3145 6873
rect 3145 6847 3146 6873
rect 3118 6846 3146 6847
rect 3118 6713 3146 6714
rect 3118 6687 3119 6713
rect 3119 6687 3145 6713
rect 3145 6687 3146 6713
rect 3118 6686 3146 6687
rect 3118 6553 3146 6554
rect 3118 6527 3119 6553
rect 3119 6527 3145 6553
rect 3145 6527 3146 6553
rect 3118 6526 3146 6527
rect 3118 6393 3146 6394
rect 3118 6367 3119 6393
rect 3119 6367 3145 6393
rect 3145 6367 3146 6393
rect 3118 6366 3146 6367
rect 3118 6233 3146 6234
rect 3118 6207 3119 6233
rect 3119 6207 3145 6233
rect 3145 6207 3146 6233
rect 3118 6206 3146 6207
rect 3118 6073 3146 6074
rect 3118 6047 3119 6073
rect 3119 6047 3145 6073
rect 3145 6047 3146 6073
rect 3118 6046 3146 6047
rect 3118 5913 3146 5914
rect 3118 5887 3119 5913
rect 3119 5887 3145 5913
rect 3145 5887 3146 5913
rect 3118 5886 3146 5887
rect 6851 9113 6879 9114
rect 6851 9087 6852 9113
rect 6852 9087 6878 9113
rect 6878 9087 6879 9113
rect 6851 9086 6879 9087
rect 6851 8953 6879 8954
rect 6851 8927 6852 8953
rect 6852 8927 6878 8953
rect 6878 8927 6879 8953
rect 6851 8926 6879 8927
rect 6851 8793 6879 8794
rect 6851 8767 6852 8793
rect 6852 8767 6878 8793
rect 6878 8767 6879 8793
rect 6851 8766 6879 8767
rect 6851 8633 6879 8634
rect 6851 8607 6852 8633
rect 6852 8607 6878 8633
rect 6878 8607 6879 8633
rect 6851 8606 6879 8607
rect 6851 8473 6879 8474
rect 6851 8447 6852 8473
rect 6852 8447 6878 8473
rect 6878 8447 6879 8473
rect 6851 8446 6879 8447
rect 6851 8313 6879 8314
rect 6851 8287 6852 8313
rect 6852 8287 6878 8313
rect 6878 8287 6879 8313
rect 6851 8286 6879 8287
rect 6851 8153 6879 8154
rect 6851 8127 6852 8153
rect 6852 8127 6878 8153
rect 6878 8127 6879 8153
rect 6851 8126 6879 8127
rect 6851 7993 6879 7994
rect 6851 7967 6852 7993
rect 6852 7967 6878 7993
rect 6878 7967 6879 7993
rect 6851 7966 6879 7967
rect 6851 7833 6879 7834
rect 6851 7807 6852 7833
rect 6852 7807 6878 7833
rect 6878 7807 6879 7833
rect 6851 7806 6879 7807
rect 6851 7673 6879 7674
rect 6851 7647 6852 7673
rect 6852 7647 6878 7673
rect 6878 7647 6879 7673
rect 6851 7646 6879 7647
rect 6851 7513 6879 7514
rect 6851 7487 6852 7513
rect 6852 7487 6878 7513
rect 6878 7487 6879 7513
rect 6851 7486 6879 7487
rect 6851 7353 6879 7354
rect 6851 7327 6852 7353
rect 6852 7327 6878 7353
rect 6878 7327 6879 7353
rect 6851 7326 6879 7327
rect 6851 7193 6879 7194
rect 6851 7167 6852 7193
rect 6852 7167 6878 7193
rect 6878 7167 6879 7193
rect 6851 7166 6879 7167
rect 6851 7033 6879 7034
rect 6851 7007 6852 7033
rect 6852 7007 6878 7033
rect 6878 7007 6879 7033
rect 6851 7006 6879 7007
rect 6851 6873 6879 6874
rect 6851 6847 6852 6873
rect 6852 6847 6878 6873
rect 6878 6847 6879 6873
rect 6851 6846 6879 6847
rect 6851 6713 6879 6714
rect 6851 6687 6852 6713
rect 6852 6687 6878 6713
rect 6878 6687 6879 6713
rect 6851 6686 6879 6687
rect 6851 6553 6879 6554
rect 6851 6527 6852 6553
rect 6852 6527 6878 6553
rect 6878 6527 6879 6553
rect 6851 6526 6879 6527
rect 6851 6393 6879 6394
rect 6851 6367 6852 6393
rect 6852 6367 6878 6393
rect 6878 6367 6879 6393
rect 6851 6366 6879 6367
rect 6851 6233 6879 6234
rect 6851 6207 6852 6233
rect 6852 6207 6878 6233
rect 6878 6207 6879 6233
rect 6851 6206 6879 6207
rect 6851 6073 6879 6074
rect 6851 6047 6852 6073
rect 6852 6047 6878 6073
rect 6878 6047 6879 6073
rect 6851 6046 6879 6047
rect 6851 5913 6879 5914
rect 6851 5887 6852 5913
rect 6852 5887 6878 5913
rect 6878 5887 6879 5913
rect 6851 5886 6879 5887
rect 3118 5753 3146 5754
rect 3118 5727 3119 5753
rect 3119 5727 3145 5753
rect 3145 5727 3146 5753
rect 3118 5726 3146 5727
rect 6851 5753 6879 5754
rect 6851 5727 6852 5753
rect 6852 5727 6878 5753
rect 6878 5727 6879 5753
rect 6851 5726 6879 5727
rect 3306 5650 3334 5651
rect 3306 5624 3307 5650
rect 3307 5624 3333 5650
rect 3333 5624 3334 5650
rect 3306 5623 3334 5624
rect 3466 5650 3494 5651
rect 3466 5624 3467 5650
rect 3467 5624 3493 5650
rect 3493 5624 3494 5650
rect 3466 5623 3494 5624
rect 3626 5650 3654 5651
rect 3626 5624 3627 5650
rect 3627 5624 3653 5650
rect 3653 5624 3654 5650
rect 3626 5623 3654 5624
rect 3786 5650 3814 5651
rect 3786 5624 3787 5650
rect 3787 5624 3813 5650
rect 3813 5624 3814 5650
rect 3786 5623 3814 5624
rect 3946 5650 3974 5651
rect 3946 5624 3947 5650
rect 3947 5624 3973 5650
rect 3973 5624 3974 5650
rect 3946 5623 3974 5624
rect 4106 5650 4134 5651
rect 4106 5624 4107 5650
rect 4107 5624 4133 5650
rect 4133 5624 4134 5650
rect 4106 5623 4134 5624
rect 4266 5650 4294 5651
rect 4266 5624 4267 5650
rect 4267 5624 4293 5650
rect 4293 5624 4294 5650
rect 4266 5623 4294 5624
rect 4426 5650 4454 5651
rect 4426 5624 4427 5650
rect 4427 5624 4453 5650
rect 4453 5624 4454 5650
rect 4426 5623 4454 5624
rect 4586 5650 4614 5651
rect 4586 5624 4587 5650
rect 4587 5624 4613 5650
rect 4613 5624 4614 5650
rect 4586 5623 4614 5624
rect 4746 5650 4774 5651
rect 4746 5624 4747 5650
rect 4747 5624 4773 5650
rect 4773 5624 4774 5650
rect 4746 5623 4774 5624
rect 4906 5650 4934 5651
rect 4906 5624 4907 5650
rect 4907 5624 4933 5650
rect 4933 5624 4934 5650
rect 4906 5623 4934 5624
rect 5066 5650 5094 5651
rect 5066 5624 5067 5650
rect 5067 5624 5093 5650
rect 5093 5624 5094 5650
rect 5066 5623 5094 5624
rect 5226 5650 5254 5651
rect 5226 5624 5227 5650
rect 5227 5624 5253 5650
rect 5253 5624 5254 5650
rect 5226 5623 5254 5624
rect 5386 5650 5414 5651
rect 5386 5624 5387 5650
rect 5387 5624 5413 5650
rect 5413 5624 5414 5650
rect 5386 5623 5414 5624
rect 5546 5650 5574 5651
rect 5546 5624 5547 5650
rect 5547 5624 5573 5650
rect 5573 5624 5574 5650
rect 5546 5623 5574 5624
rect 5706 5650 5734 5651
rect 5706 5624 5707 5650
rect 5707 5624 5733 5650
rect 5733 5624 5734 5650
rect 5706 5623 5734 5624
rect 5866 5650 5894 5651
rect 5866 5624 5867 5650
rect 5867 5624 5893 5650
rect 5893 5624 5894 5650
rect 5866 5623 5894 5624
rect 6026 5650 6054 5651
rect 6026 5624 6027 5650
rect 6027 5624 6053 5650
rect 6053 5624 6054 5650
rect 6026 5623 6054 5624
rect 6186 5650 6214 5651
rect 6186 5624 6187 5650
rect 6187 5624 6213 5650
rect 6213 5624 6214 5650
rect 6186 5623 6214 5624
rect 6346 5650 6374 5651
rect 6346 5624 6347 5650
rect 6347 5624 6373 5650
rect 6373 5624 6374 5650
rect 6346 5623 6374 5624
rect 6506 5650 6534 5651
rect 6506 5624 6507 5650
rect 6507 5624 6533 5650
rect 6533 5624 6534 5650
rect 6506 5623 6534 5624
rect 6666 5650 6694 5651
rect 6666 5624 6667 5650
rect 6667 5624 6693 5650
rect 6693 5624 6694 5650
rect 6666 5623 6694 5624
rect 9306 9378 9334 9379
rect 9306 9352 9307 9378
rect 9307 9352 9333 9378
rect 9333 9352 9334 9378
rect 9306 9351 9334 9352
rect 9466 9378 9494 9379
rect 9466 9352 9467 9378
rect 9467 9352 9493 9378
rect 9493 9352 9494 9378
rect 9466 9351 9494 9352
rect 9626 9378 9654 9379
rect 9626 9352 9627 9378
rect 9627 9352 9653 9378
rect 9653 9352 9654 9378
rect 9626 9351 9654 9352
rect 9786 9378 9814 9379
rect 9786 9352 9787 9378
rect 9787 9352 9813 9378
rect 9813 9352 9814 9378
rect 9786 9351 9814 9352
rect 9946 9378 9974 9379
rect 9946 9352 9947 9378
rect 9947 9352 9973 9378
rect 9973 9352 9974 9378
rect 9946 9351 9974 9352
rect 10106 9378 10134 9379
rect 10106 9352 10107 9378
rect 10107 9352 10133 9378
rect 10133 9352 10134 9378
rect 10106 9351 10134 9352
rect 10266 9378 10294 9379
rect 10266 9352 10267 9378
rect 10267 9352 10293 9378
rect 10293 9352 10294 9378
rect 10266 9351 10294 9352
rect 10426 9378 10454 9379
rect 10426 9352 10427 9378
rect 10427 9352 10453 9378
rect 10453 9352 10454 9378
rect 10426 9351 10454 9352
rect 10586 9378 10614 9379
rect 10586 9352 10587 9378
rect 10587 9352 10613 9378
rect 10613 9352 10614 9378
rect 10586 9351 10614 9352
rect 10746 9378 10774 9379
rect 10746 9352 10747 9378
rect 10747 9352 10773 9378
rect 10773 9352 10774 9378
rect 10746 9351 10774 9352
rect 10906 9378 10934 9379
rect 10906 9352 10907 9378
rect 10907 9352 10933 9378
rect 10933 9352 10934 9378
rect 10906 9351 10934 9352
rect 11066 9378 11094 9379
rect 11066 9352 11067 9378
rect 11067 9352 11093 9378
rect 11093 9352 11094 9378
rect 11066 9351 11094 9352
rect 11226 9378 11254 9379
rect 11226 9352 11227 9378
rect 11227 9352 11253 9378
rect 11253 9352 11254 9378
rect 11226 9351 11254 9352
rect 11386 9378 11414 9379
rect 11386 9352 11387 9378
rect 11387 9352 11413 9378
rect 11413 9352 11414 9378
rect 11386 9351 11414 9352
rect 11546 9378 11574 9379
rect 11546 9352 11547 9378
rect 11547 9352 11573 9378
rect 11573 9352 11574 9378
rect 11546 9351 11574 9352
rect 11706 9378 11734 9379
rect 11706 9352 11707 9378
rect 11707 9352 11733 9378
rect 11733 9352 11734 9378
rect 11706 9351 11734 9352
rect 11866 9378 11894 9379
rect 11866 9352 11867 9378
rect 11867 9352 11893 9378
rect 11893 9352 11894 9378
rect 11866 9351 11894 9352
rect 12026 9378 12054 9379
rect 12026 9352 12027 9378
rect 12027 9352 12053 9378
rect 12053 9352 12054 9378
rect 12026 9351 12054 9352
rect 12186 9378 12214 9379
rect 12186 9352 12187 9378
rect 12187 9352 12213 9378
rect 12213 9352 12214 9378
rect 12186 9351 12214 9352
rect 12346 9378 12374 9379
rect 12346 9352 12347 9378
rect 12347 9352 12373 9378
rect 12373 9352 12374 9378
rect 12346 9351 12374 9352
rect 12506 9378 12534 9379
rect 12506 9352 12507 9378
rect 12507 9352 12533 9378
rect 12533 9352 12534 9378
rect 12506 9351 12534 9352
rect 12666 9378 12694 9379
rect 12666 9352 12667 9378
rect 12667 9352 12693 9378
rect 12693 9352 12694 9378
rect 12666 9351 12694 9352
rect 9118 9273 9146 9274
rect 9118 9247 9119 9273
rect 9119 9247 9145 9273
rect 9145 9247 9146 9273
rect 9118 9246 9146 9247
rect 12851 9273 12879 9274
rect 12851 9247 12852 9273
rect 12852 9247 12878 9273
rect 12878 9247 12879 9273
rect 12851 9246 12879 9247
rect 9118 9113 9146 9114
rect 9118 9087 9119 9113
rect 9119 9087 9145 9113
rect 9145 9087 9146 9113
rect 9118 9086 9146 9087
rect 9118 8953 9146 8954
rect 9118 8927 9119 8953
rect 9119 8927 9145 8953
rect 9145 8927 9146 8953
rect 9118 8926 9146 8927
rect 9118 8793 9146 8794
rect 9118 8767 9119 8793
rect 9119 8767 9145 8793
rect 9145 8767 9146 8793
rect 9118 8766 9146 8767
rect 9118 8633 9146 8634
rect 9118 8607 9119 8633
rect 9119 8607 9145 8633
rect 9145 8607 9146 8633
rect 9118 8606 9146 8607
rect 9118 8473 9146 8474
rect 9118 8447 9119 8473
rect 9119 8447 9145 8473
rect 9145 8447 9146 8473
rect 9118 8446 9146 8447
rect 9118 8313 9146 8314
rect 9118 8287 9119 8313
rect 9119 8287 9145 8313
rect 9145 8287 9146 8313
rect 9118 8286 9146 8287
rect 9118 8153 9146 8154
rect 9118 8127 9119 8153
rect 9119 8127 9145 8153
rect 9145 8127 9146 8153
rect 9118 8126 9146 8127
rect 9118 7993 9146 7994
rect 9118 7967 9119 7993
rect 9119 7967 9145 7993
rect 9145 7967 9146 7993
rect 9118 7966 9146 7967
rect 9118 7833 9146 7834
rect 9118 7807 9119 7833
rect 9119 7807 9145 7833
rect 9145 7807 9146 7833
rect 9118 7806 9146 7807
rect 9118 7673 9146 7674
rect 9118 7647 9119 7673
rect 9119 7647 9145 7673
rect 9145 7647 9146 7673
rect 9118 7646 9146 7647
rect 9118 7513 9146 7514
rect 9118 7487 9119 7513
rect 9119 7487 9145 7513
rect 9145 7487 9146 7513
rect 9118 7486 9146 7487
rect 9118 7353 9146 7354
rect 9118 7327 9119 7353
rect 9119 7327 9145 7353
rect 9145 7327 9146 7353
rect 9118 7326 9146 7327
rect 9118 7193 9146 7194
rect 9118 7167 9119 7193
rect 9119 7167 9145 7193
rect 9145 7167 9146 7193
rect 9118 7166 9146 7167
rect 9118 7033 9146 7034
rect 9118 7007 9119 7033
rect 9119 7007 9145 7033
rect 9145 7007 9146 7033
rect 9118 7006 9146 7007
rect 9118 6873 9146 6874
rect 9118 6847 9119 6873
rect 9119 6847 9145 6873
rect 9145 6847 9146 6873
rect 9118 6846 9146 6847
rect 9118 6713 9146 6714
rect 9118 6687 9119 6713
rect 9119 6687 9145 6713
rect 9145 6687 9146 6713
rect 9118 6686 9146 6687
rect 9118 6553 9146 6554
rect 9118 6527 9119 6553
rect 9119 6527 9145 6553
rect 9145 6527 9146 6553
rect 9118 6526 9146 6527
rect 9118 6393 9146 6394
rect 9118 6367 9119 6393
rect 9119 6367 9145 6393
rect 9145 6367 9146 6393
rect 9118 6366 9146 6367
rect 9118 6233 9146 6234
rect 9118 6207 9119 6233
rect 9119 6207 9145 6233
rect 9145 6207 9146 6233
rect 9118 6206 9146 6207
rect 9118 6073 9146 6074
rect 9118 6047 9119 6073
rect 9119 6047 9145 6073
rect 9145 6047 9146 6073
rect 9118 6046 9146 6047
rect 9118 5913 9146 5914
rect 9118 5887 9119 5913
rect 9119 5887 9145 5913
rect 9145 5887 9146 5913
rect 9118 5886 9146 5887
rect 12851 9113 12879 9114
rect 12851 9087 12852 9113
rect 12852 9087 12878 9113
rect 12878 9087 12879 9113
rect 12851 9086 12879 9087
rect 12851 8953 12879 8954
rect 12851 8927 12852 8953
rect 12852 8927 12878 8953
rect 12878 8927 12879 8953
rect 12851 8926 12879 8927
rect 12851 8793 12879 8794
rect 12851 8767 12852 8793
rect 12852 8767 12878 8793
rect 12878 8767 12879 8793
rect 12851 8766 12879 8767
rect 12851 8633 12879 8634
rect 12851 8607 12852 8633
rect 12852 8607 12878 8633
rect 12878 8607 12879 8633
rect 12851 8606 12879 8607
rect 12851 8473 12879 8474
rect 12851 8447 12852 8473
rect 12852 8447 12878 8473
rect 12878 8447 12879 8473
rect 12851 8446 12879 8447
rect 12851 8313 12879 8314
rect 12851 8287 12852 8313
rect 12852 8287 12878 8313
rect 12878 8287 12879 8313
rect 12851 8286 12879 8287
rect 12851 8153 12879 8154
rect 12851 8127 12852 8153
rect 12852 8127 12878 8153
rect 12878 8127 12879 8153
rect 12851 8126 12879 8127
rect 12851 7993 12879 7994
rect 12851 7967 12852 7993
rect 12852 7967 12878 7993
rect 12878 7967 12879 7993
rect 12851 7966 12879 7967
rect 12851 7833 12879 7834
rect 12851 7807 12852 7833
rect 12852 7807 12878 7833
rect 12878 7807 12879 7833
rect 12851 7806 12879 7807
rect 12851 7673 12879 7674
rect 12851 7647 12852 7673
rect 12852 7647 12878 7673
rect 12878 7647 12879 7673
rect 12851 7646 12879 7647
rect 12851 7513 12879 7514
rect 12851 7487 12852 7513
rect 12852 7487 12878 7513
rect 12878 7487 12879 7513
rect 12851 7486 12879 7487
rect 12851 7353 12879 7354
rect 12851 7327 12852 7353
rect 12852 7327 12878 7353
rect 12878 7327 12879 7353
rect 12851 7326 12879 7327
rect 12851 7193 12879 7194
rect 12851 7167 12852 7193
rect 12852 7167 12878 7193
rect 12878 7167 12879 7193
rect 12851 7166 12879 7167
rect 12851 7033 12879 7034
rect 12851 7007 12852 7033
rect 12852 7007 12878 7033
rect 12878 7007 12879 7033
rect 12851 7006 12879 7007
rect 12851 6873 12879 6874
rect 12851 6847 12852 6873
rect 12852 6847 12878 6873
rect 12878 6847 12879 6873
rect 12851 6846 12879 6847
rect 12851 6713 12879 6714
rect 12851 6687 12852 6713
rect 12852 6687 12878 6713
rect 12878 6687 12879 6713
rect 12851 6686 12879 6687
rect 12851 6553 12879 6554
rect 12851 6527 12852 6553
rect 12852 6527 12878 6553
rect 12878 6527 12879 6553
rect 12851 6526 12879 6527
rect 12851 6393 12879 6394
rect 12851 6367 12852 6393
rect 12852 6367 12878 6393
rect 12878 6367 12879 6393
rect 12851 6366 12879 6367
rect 12851 6233 12879 6234
rect 12851 6207 12852 6233
rect 12852 6207 12878 6233
rect 12878 6207 12879 6233
rect 12851 6206 12879 6207
rect 12851 6073 12879 6074
rect 12851 6047 12852 6073
rect 12852 6047 12878 6073
rect 12878 6047 12879 6073
rect 12851 6046 12879 6047
rect 12851 5913 12879 5914
rect 12851 5887 12852 5913
rect 12852 5887 12878 5913
rect 12878 5887 12879 5913
rect 12851 5886 12879 5887
rect 9118 5753 9146 5754
rect 9118 5727 9119 5753
rect 9119 5727 9145 5753
rect 9145 5727 9146 5753
rect 9118 5726 9146 5727
rect 12851 5753 12879 5754
rect 12851 5727 12852 5753
rect 12852 5727 12878 5753
rect 12878 5727 12879 5753
rect 12851 5726 12879 5727
rect 9306 5650 9334 5651
rect 9306 5624 9307 5650
rect 9307 5624 9333 5650
rect 9333 5624 9334 5650
rect 9306 5623 9334 5624
rect 9466 5650 9494 5651
rect 9466 5624 9467 5650
rect 9467 5624 9493 5650
rect 9493 5624 9494 5650
rect 9466 5623 9494 5624
rect 9626 5650 9654 5651
rect 9626 5624 9627 5650
rect 9627 5624 9653 5650
rect 9653 5624 9654 5650
rect 9626 5623 9654 5624
rect 9786 5650 9814 5651
rect 9786 5624 9787 5650
rect 9787 5624 9813 5650
rect 9813 5624 9814 5650
rect 9786 5623 9814 5624
rect 9946 5650 9974 5651
rect 9946 5624 9947 5650
rect 9947 5624 9973 5650
rect 9973 5624 9974 5650
rect 9946 5623 9974 5624
rect 10106 5650 10134 5651
rect 10106 5624 10107 5650
rect 10107 5624 10133 5650
rect 10133 5624 10134 5650
rect 10106 5623 10134 5624
rect 10266 5650 10294 5651
rect 10266 5624 10267 5650
rect 10267 5624 10293 5650
rect 10293 5624 10294 5650
rect 10266 5623 10294 5624
rect 10426 5650 10454 5651
rect 10426 5624 10427 5650
rect 10427 5624 10453 5650
rect 10453 5624 10454 5650
rect 10426 5623 10454 5624
rect 10586 5650 10614 5651
rect 10586 5624 10587 5650
rect 10587 5624 10613 5650
rect 10613 5624 10614 5650
rect 10586 5623 10614 5624
rect 10746 5650 10774 5651
rect 10746 5624 10747 5650
rect 10747 5624 10773 5650
rect 10773 5624 10774 5650
rect 10746 5623 10774 5624
rect 10906 5650 10934 5651
rect 10906 5624 10907 5650
rect 10907 5624 10933 5650
rect 10933 5624 10934 5650
rect 10906 5623 10934 5624
rect 11066 5650 11094 5651
rect 11066 5624 11067 5650
rect 11067 5624 11093 5650
rect 11093 5624 11094 5650
rect 11066 5623 11094 5624
rect 11226 5650 11254 5651
rect 11226 5624 11227 5650
rect 11227 5624 11253 5650
rect 11253 5624 11254 5650
rect 11226 5623 11254 5624
rect 11386 5650 11414 5651
rect 11386 5624 11387 5650
rect 11387 5624 11413 5650
rect 11413 5624 11414 5650
rect 11386 5623 11414 5624
rect 11546 5650 11574 5651
rect 11546 5624 11547 5650
rect 11547 5624 11573 5650
rect 11573 5624 11574 5650
rect 11546 5623 11574 5624
rect 11706 5650 11734 5651
rect 11706 5624 11707 5650
rect 11707 5624 11733 5650
rect 11733 5624 11734 5650
rect 11706 5623 11734 5624
rect 11866 5650 11894 5651
rect 11866 5624 11867 5650
rect 11867 5624 11893 5650
rect 11893 5624 11894 5650
rect 11866 5623 11894 5624
rect 12026 5650 12054 5651
rect 12026 5624 12027 5650
rect 12027 5624 12053 5650
rect 12053 5624 12054 5650
rect 12026 5623 12054 5624
rect 12186 5650 12214 5651
rect 12186 5624 12187 5650
rect 12187 5624 12213 5650
rect 12213 5624 12214 5650
rect 12186 5623 12214 5624
rect 12346 5650 12374 5651
rect 12346 5624 12347 5650
rect 12347 5624 12373 5650
rect 12373 5624 12374 5650
rect 12346 5623 12374 5624
rect 12506 5650 12534 5651
rect 12506 5624 12507 5650
rect 12507 5624 12533 5650
rect 12533 5624 12534 5650
rect 12506 5623 12534 5624
rect 12666 5650 12694 5651
rect 12666 5624 12667 5650
rect 12667 5624 12693 5650
rect 12693 5624 12694 5650
rect 12666 5623 12694 5624
rect 15306 9378 15334 9379
rect 15306 9352 15307 9378
rect 15307 9352 15333 9378
rect 15333 9352 15334 9378
rect 15306 9351 15334 9352
rect 15466 9378 15494 9379
rect 15466 9352 15467 9378
rect 15467 9352 15493 9378
rect 15493 9352 15494 9378
rect 15466 9351 15494 9352
rect 15626 9378 15654 9379
rect 15626 9352 15627 9378
rect 15627 9352 15653 9378
rect 15653 9352 15654 9378
rect 15626 9351 15654 9352
rect 15786 9378 15814 9379
rect 15786 9352 15787 9378
rect 15787 9352 15813 9378
rect 15813 9352 15814 9378
rect 15786 9351 15814 9352
rect 15946 9378 15974 9379
rect 15946 9352 15947 9378
rect 15947 9352 15973 9378
rect 15973 9352 15974 9378
rect 15946 9351 15974 9352
rect 16106 9378 16134 9379
rect 16106 9352 16107 9378
rect 16107 9352 16133 9378
rect 16133 9352 16134 9378
rect 16106 9351 16134 9352
rect 16266 9378 16294 9379
rect 16266 9352 16267 9378
rect 16267 9352 16293 9378
rect 16293 9352 16294 9378
rect 16266 9351 16294 9352
rect 16426 9378 16454 9379
rect 16426 9352 16427 9378
rect 16427 9352 16453 9378
rect 16453 9352 16454 9378
rect 16426 9351 16454 9352
rect 16586 9378 16614 9379
rect 16586 9352 16587 9378
rect 16587 9352 16613 9378
rect 16613 9352 16614 9378
rect 16586 9351 16614 9352
rect 16746 9378 16774 9379
rect 16746 9352 16747 9378
rect 16747 9352 16773 9378
rect 16773 9352 16774 9378
rect 16746 9351 16774 9352
rect 16906 9378 16934 9379
rect 16906 9352 16907 9378
rect 16907 9352 16933 9378
rect 16933 9352 16934 9378
rect 16906 9351 16934 9352
rect 17066 9378 17094 9379
rect 17066 9352 17067 9378
rect 17067 9352 17093 9378
rect 17093 9352 17094 9378
rect 17066 9351 17094 9352
rect 17226 9378 17254 9379
rect 17226 9352 17227 9378
rect 17227 9352 17253 9378
rect 17253 9352 17254 9378
rect 17226 9351 17254 9352
rect 17386 9378 17414 9379
rect 17386 9352 17387 9378
rect 17387 9352 17413 9378
rect 17413 9352 17414 9378
rect 17386 9351 17414 9352
rect 17546 9378 17574 9379
rect 17546 9352 17547 9378
rect 17547 9352 17573 9378
rect 17573 9352 17574 9378
rect 17546 9351 17574 9352
rect 17706 9378 17734 9379
rect 17706 9352 17707 9378
rect 17707 9352 17733 9378
rect 17733 9352 17734 9378
rect 17706 9351 17734 9352
rect 17866 9378 17894 9379
rect 17866 9352 17867 9378
rect 17867 9352 17893 9378
rect 17893 9352 17894 9378
rect 17866 9351 17894 9352
rect 18026 9378 18054 9379
rect 18026 9352 18027 9378
rect 18027 9352 18053 9378
rect 18053 9352 18054 9378
rect 18026 9351 18054 9352
rect 18186 9378 18214 9379
rect 18186 9352 18187 9378
rect 18187 9352 18213 9378
rect 18213 9352 18214 9378
rect 18186 9351 18214 9352
rect 18346 9378 18374 9379
rect 18346 9352 18347 9378
rect 18347 9352 18373 9378
rect 18373 9352 18374 9378
rect 18346 9351 18374 9352
rect 18506 9378 18534 9379
rect 18506 9352 18507 9378
rect 18507 9352 18533 9378
rect 18533 9352 18534 9378
rect 18506 9351 18534 9352
rect 18666 9378 18694 9379
rect 18666 9352 18667 9378
rect 18667 9352 18693 9378
rect 18693 9352 18694 9378
rect 18666 9351 18694 9352
rect 15118 9273 15146 9274
rect 15118 9247 15119 9273
rect 15119 9247 15145 9273
rect 15145 9247 15146 9273
rect 15118 9246 15146 9247
rect 18851 9273 18879 9274
rect 18851 9247 18852 9273
rect 18852 9247 18878 9273
rect 18878 9247 18879 9273
rect 18851 9246 18879 9247
rect 15118 9113 15146 9114
rect 15118 9087 15119 9113
rect 15119 9087 15145 9113
rect 15145 9087 15146 9113
rect 15118 9086 15146 9087
rect 15118 8953 15146 8954
rect 15118 8927 15119 8953
rect 15119 8927 15145 8953
rect 15145 8927 15146 8953
rect 15118 8926 15146 8927
rect 15118 8793 15146 8794
rect 15118 8767 15119 8793
rect 15119 8767 15145 8793
rect 15145 8767 15146 8793
rect 15118 8766 15146 8767
rect 15118 8633 15146 8634
rect 15118 8607 15119 8633
rect 15119 8607 15145 8633
rect 15145 8607 15146 8633
rect 15118 8606 15146 8607
rect 15118 8473 15146 8474
rect 15118 8447 15119 8473
rect 15119 8447 15145 8473
rect 15145 8447 15146 8473
rect 15118 8446 15146 8447
rect 15118 8313 15146 8314
rect 15118 8287 15119 8313
rect 15119 8287 15145 8313
rect 15145 8287 15146 8313
rect 15118 8286 15146 8287
rect 15118 8153 15146 8154
rect 15118 8127 15119 8153
rect 15119 8127 15145 8153
rect 15145 8127 15146 8153
rect 15118 8126 15146 8127
rect 15118 7993 15146 7994
rect 15118 7967 15119 7993
rect 15119 7967 15145 7993
rect 15145 7967 15146 7993
rect 15118 7966 15146 7967
rect 15118 7833 15146 7834
rect 15118 7807 15119 7833
rect 15119 7807 15145 7833
rect 15145 7807 15146 7833
rect 15118 7806 15146 7807
rect 15118 7673 15146 7674
rect 15118 7647 15119 7673
rect 15119 7647 15145 7673
rect 15145 7647 15146 7673
rect 15118 7646 15146 7647
rect 15118 7513 15146 7514
rect 15118 7487 15119 7513
rect 15119 7487 15145 7513
rect 15145 7487 15146 7513
rect 15118 7486 15146 7487
rect 15118 7353 15146 7354
rect 15118 7327 15119 7353
rect 15119 7327 15145 7353
rect 15145 7327 15146 7353
rect 15118 7326 15146 7327
rect 15118 7193 15146 7194
rect 15118 7167 15119 7193
rect 15119 7167 15145 7193
rect 15145 7167 15146 7193
rect 15118 7166 15146 7167
rect 15118 7033 15146 7034
rect 15118 7007 15119 7033
rect 15119 7007 15145 7033
rect 15145 7007 15146 7033
rect 15118 7006 15146 7007
rect 15118 6873 15146 6874
rect 15118 6847 15119 6873
rect 15119 6847 15145 6873
rect 15145 6847 15146 6873
rect 15118 6846 15146 6847
rect 15118 6713 15146 6714
rect 15118 6687 15119 6713
rect 15119 6687 15145 6713
rect 15145 6687 15146 6713
rect 15118 6686 15146 6687
rect 15118 6553 15146 6554
rect 15118 6527 15119 6553
rect 15119 6527 15145 6553
rect 15145 6527 15146 6553
rect 15118 6526 15146 6527
rect 15118 6393 15146 6394
rect 15118 6367 15119 6393
rect 15119 6367 15145 6393
rect 15145 6367 15146 6393
rect 15118 6366 15146 6367
rect 15118 6233 15146 6234
rect 15118 6207 15119 6233
rect 15119 6207 15145 6233
rect 15145 6207 15146 6233
rect 15118 6206 15146 6207
rect 15118 6073 15146 6074
rect 15118 6047 15119 6073
rect 15119 6047 15145 6073
rect 15145 6047 15146 6073
rect 15118 6046 15146 6047
rect 15118 5913 15146 5914
rect 15118 5887 15119 5913
rect 15119 5887 15145 5913
rect 15145 5887 15146 5913
rect 15118 5886 15146 5887
rect 18851 9113 18879 9114
rect 18851 9087 18852 9113
rect 18852 9087 18878 9113
rect 18878 9087 18879 9113
rect 18851 9086 18879 9087
rect 18851 8953 18879 8954
rect 18851 8927 18852 8953
rect 18852 8927 18878 8953
rect 18878 8927 18879 8953
rect 18851 8926 18879 8927
rect 18851 8793 18879 8794
rect 18851 8767 18852 8793
rect 18852 8767 18878 8793
rect 18878 8767 18879 8793
rect 18851 8766 18879 8767
rect 18851 8633 18879 8634
rect 18851 8607 18852 8633
rect 18852 8607 18878 8633
rect 18878 8607 18879 8633
rect 18851 8606 18879 8607
rect 18851 8473 18879 8474
rect 18851 8447 18852 8473
rect 18852 8447 18878 8473
rect 18878 8447 18879 8473
rect 18851 8446 18879 8447
rect 18851 8313 18879 8314
rect 18851 8287 18852 8313
rect 18852 8287 18878 8313
rect 18878 8287 18879 8313
rect 18851 8286 18879 8287
rect 18851 8153 18879 8154
rect 18851 8127 18852 8153
rect 18852 8127 18878 8153
rect 18878 8127 18879 8153
rect 18851 8126 18879 8127
rect 18851 7993 18879 7994
rect 18851 7967 18852 7993
rect 18852 7967 18878 7993
rect 18878 7967 18879 7993
rect 18851 7966 18879 7967
rect 18851 7833 18879 7834
rect 18851 7807 18852 7833
rect 18852 7807 18878 7833
rect 18878 7807 18879 7833
rect 18851 7806 18879 7807
rect 18851 7673 18879 7674
rect 18851 7647 18852 7673
rect 18852 7647 18878 7673
rect 18878 7647 18879 7673
rect 18851 7646 18879 7647
rect 18851 7513 18879 7514
rect 18851 7487 18852 7513
rect 18852 7487 18878 7513
rect 18878 7487 18879 7513
rect 18851 7486 18879 7487
rect 18851 7353 18879 7354
rect 18851 7327 18852 7353
rect 18852 7327 18878 7353
rect 18878 7327 18879 7353
rect 18851 7326 18879 7327
rect 18851 7193 18879 7194
rect 18851 7167 18852 7193
rect 18852 7167 18878 7193
rect 18878 7167 18879 7193
rect 18851 7166 18879 7167
rect 18851 7033 18879 7034
rect 18851 7007 18852 7033
rect 18852 7007 18878 7033
rect 18878 7007 18879 7033
rect 18851 7006 18879 7007
rect 18851 6873 18879 6874
rect 18851 6847 18852 6873
rect 18852 6847 18878 6873
rect 18878 6847 18879 6873
rect 18851 6846 18879 6847
rect 18851 6713 18879 6714
rect 18851 6687 18852 6713
rect 18852 6687 18878 6713
rect 18878 6687 18879 6713
rect 18851 6686 18879 6687
rect 18851 6553 18879 6554
rect 18851 6527 18852 6553
rect 18852 6527 18878 6553
rect 18878 6527 18879 6553
rect 18851 6526 18879 6527
rect 18851 6393 18879 6394
rect 18851 6367 18852 6393
rect 18852 6367 18878 6393
rect 18878 6367 18879 6393
rect 18851 6366 18879 6367
rect 18851 6233 18879 6234
rect 18851 6207 18852 6233
rect 18852 6207 18878 6233
rect 18878 6207 18879 6233
rect 18851 6206 18879 6207
rect 18851 6073 18879 6074
rect 18851 6047 18852 6073
rect 18852 6047 18878 6073
rect 18878 6047 18879 6073
rect 18851 6046 18879 6047
rect 18851 5913 18879 5914
rect 18851 5887 18852 5913
rect 18852 5887 18878 5913
rect 18878 5887 18879 5913
rect 18851 5886 18879 5887
rect 15118 5753 15146 5754
rect 15118 5727 15119 5753
rect 15119 5727 15145 5753
rect 15145 5727 15146 5753
rect 15118 5726 15146 5727
rect 18851 5753 18879 5754
rect 18851 5727 18852 5753
rect 18852 5727 18878 5753
rect 18878 5727 18879 5753
rect 18851 5726 18879 5727
rect 15306 5650 15334 5651
rect 15306 5624 15307 5650
rect 15307 5624 15333 5650
rect 15333 5624 15334 5650
rect 15306 5623 15334 5624
rect 15466 5650 15494 5651
rect 15466 5624 15467 5650
rect 15467 5624 15493 5650
rect 15493 5624 15494 5650
rect 15466 5623 15494 5624
rect 15626 5650 15654 5651
rect 15626 5624 15627 5650
rect 15627 5624 15653 5650
rect 15653 5624 15654 5650
rect 15626 5623 15654 5624
rect 15786 5650 15814 5651
rect 15786 5624 15787 5650
rect 15787 5624 15813 5650
rect 15813 5624 15814 5650
rect 15786 5623 15814 5624
rect 15946 5650 15974 5651
rect 15946 5624 15947 5650
rect 15947 5624 15973 5650
rect 15973 5624 15974 5650
rect 15946 5623 15974 5624
rect 16106 5650 16134 5651
rect 16106 5624 16107 5650
rect 16107 5624 16133 5650
rect 16133 5624 16134 5650
rect 16106 5623 16134 5624
rect 16266 5650 16294 5651
rect 16266 5624 16267 5650
rect 16267 5624 16293 5650
rect 16293 5624 16294 5650
rect 16266 5623 16294 5624
rect 16426 5650 16454 5651
rect 16426 5624 16427 5650
rect 16427 5624 16453 5650
rect 16453 5624 16454 5650
rect 16426 5623 16454 5624
rect 16586 5650 16614 5651
rect 16586 5624 16587 5650
rect 16587 5624 16613 5650
rect 16613 5624 16614 5650
rect 16586 5623 16614 5624
rect 16746 5650 16774 5651
rect 16746 5624 16747 5650
rect 16747 5624 16773 5650
rect 16773 5624 16774 5650
rect 16746 5623 16774 5624
rect 16906 5650 16934 5651
rect 16906 5624 16907 5650
rect 16907 5624 16933 5650
rect 16933 5624 16934 5650
rect 16906 5623 16934 5624
rect 17066 5650 17094 5651
rect 17066 5624 17067 5650
rect 17067 5624 17093 5650
rect 17093 5624 17094 5650
rect 17066 5623 17094 5624
rect 17226 5650 17254 5651
rect 17226 5624 17227 5650
rect 17227 5624 17253 5650
rect 17253 5624 17254 5650
rect 17226 5623 17254 5624
rect 17386 5650 17414 5651
rect 17386 5624 17387 5650
rect 17387 5624 17413 5650
rect 17413 5624 17414 5650
rect 17386 5623 17414 5624
rect 17546 5650 17574 5651
rect 17546 5624 17547 5650
rect 17547 5624 17573 5650
rect 17573 5624 17574 5650
rect 17546 5623 17574 5624
rect 17706 5650 17734 5651
rect 17706 5624 17707 5650
rect 17707 5624 17733 5650
rect 17733 5624 17734 5650
rect 17706 5623 17734 5624
rect 17866 5650 17894 5651
rect 17866 5624 17867 5650
rect 17867 5624 17893 5650
rect 17893 5624 17894 5650
rect 17866 5623 17894 5624
rect 18026 5650 18054 5651
rect 18026 5624 18027 5650
rect 18027 5624 18053 5650
rect 18053 5624 18054 5650
rect 18026 5623 18054 5624
rect 18186 5650 18214 5651
rect 18186 5624 18187 5650
rect 18187 5624 18213 5650
rect 18213 5624 18214 5650
rect 18186 5623 18214 5624
rect 18346 5650 18374 5651
rect 18346 5624 18347 5650
rect 18347 5624 18373 5650
rect 18373 5624 18374 5650
rect 18346 5623 18374 5624
rect 18506 5650 18534 5651
rect 18506 5624 18507 5650
rect 18507 5624 18533 5650
rect 18533 5624 18534 5650
rect 18506 5623 18534 5624
rect 18666 5650 18694 5651
rect 18666 5624 18667 5650
rect 18667 5624 18693 5650
rect 18693 5624 18694 5650
rect 18666 5623 18694 5624
rect 21306 9378 21334 9379
rect 21306 9352 21307 9378
rect 21307 9352 21333 9378
rect 21333 9352 21334 9378
rect 21306 9351 21334 9352
rect 21466 9378 21494 9379
rect 21466 9352 21467 9378
rect 21467 9352 21493 9378
rect 21493 9352 21494 9378
rect 21466 9351 21494 9352
rect 21626 9378 21654 9379
rect 21626 9352 21627 9378
rect 21627 9352 21653 9378
rect 21653 9352 21654 9378
rect 21626 9351 21654 9352
rect 21786 9378 21814 9379
rect 21786 9352 21787 9378
rect 21787 9352 21813 9378
rect 21813 9352 21814 9378
rect 21786 9351 21814 9352
rect 21946 9378 21974 9379
rect 21946 9352 21947 9378
rect 21947 9352 21973 9378
rect 21973 9352 21974 9378
rect 21946 9351 21974 9352
rect 22106 9378 22134 9379
rect 22106 9352 22107 9378
rect 22107 9352 22133 9378
rect 22133 9352 22134 9378
rect 22106 9351 22134 9352
rect 22266 9378 22294 9379
rect 22266 9352 22267 9378
rect 22267 9352 22293 9378
rect 22293 9352 22294 9378
rect 22266 9351 22294 9352
rect 22426 9378 22454 9379
rect 22426 9352 22427 9378
rect 22427 9352 22453 9378
rect 22453 9352 22454 9378
rect 22426 9351 22454 9352
rect 22586 9378 22614 9379
rect 22586 9352 22587 9378
rect 22587 9352 22613 9378
rect 22613 9352 22614 9378
rect 22586 9351 22614 9352
rect 22746 9378 22774 9379
rect 22746 9352 22747 9378
rect 22747 9352 22773 9378
rect 22773 9352 22774 9378
rect 22746 9351 22774 9352
rect 22906 9378 22934 9379
rect 22906 9352 22907 9378
rect 22907 9352 22933 9378
rect 22933 9352 22934 9378
rect 22906 9351 22934 9352
rect 23066 9378 23094 9379
rect 23066 9352 23067 9378
rect 23067 9352 23093 9378
rect 23093 9352 23094 9378
rect 23066 9351 23094 9352
rect 23226 9378 23254 9379
rect 23226 9352 23227 9378
rect 23227 9352 23253 9378
rect 23253 9352 23254 9378
rect 23226 9351 23254 9352
rect 23386 9378 23414 9379
rect 23386 9352 23387 9378
rect 23387 9352 23413 9378
rect 23413 9352 23414 9378
rect 23386 9351 23414 9352
rect 23546 9378 23574 9379
rect 23546 9352 23547 9378
rect 23547 9352 23573 9378
rect 23573 9352 23574 9378
rect 23546 9351 23574 9352
rect 23706 9378 23734 9379
rect 23706 9352 23707 9378
rect 23707 9352 23733 9378
rect 23733 9352 23734 9378
rect 23706 9351 23734 9352
rect 23866 9378 23894 9379
rect 23866 9352 23867 9378
rect 23867 9352 23893 9378
rect 23893 9352 23894 9378
rect 23866 9351 23894 9352
rect 24026 9378 24054 9379
rect 24026 9352 24027 9378
rect 24027 9352 24053 9378
rect 24053 9352 24054 9378
rect 24026 9351 24054 9352
rect 24186 9378 24214 9379
rect 24186 9352 24187 9378
rect 24187 9352 24213 9378
rect 24213 9352 24214 9378
rect 24186 9351 24214 9352
rect 24346 9378 24374 9379
rect 24346 9352 24347 9378
rect 24347 9352 24373 9378
rect 24373 9352 24374 9378
rect 24346 9351 24374 9352
rect 24506 9378 24534 9379
rect 24506 9352 24507 9378
rect 24507 9352 24533 9378
rect 24533 9352 24534 9378
rect 24506 9351 24534 9352
rect 24666 9378 24694 9379
rect 24666 9352 24667 9378
rect 24667 9352 24693 9378
rect 24693 9352 24694 9378
rect 24666 9351 24694 9352
rect 21118 9273 21146 9274
rect 21118 9247 21119 9273
rect 21119 9247 21145 9273
rect 21145 9247 21146 9273
rect 21118 9246 21146 9247
rect 24851 9273 24879 9274
rect 24851 9247 24852 9273
rect 24852 9247 24878 9273
rect 24878 9247 24879 9273
rect 24851 9246 24879 9247
rect 21118 9113 21146 9114
rect 21118 9087 21119 9113
rect 21119 9087 21145 9113
rect 21145 9087 21146 9113
rect 21118 9086 21146 9087
rect 21118 8953 21146 8954
rect 21118 8927 21119 8953
rect 21119 8927 21145 8953
rect 21145 8927 21146 8953
rect 21118 8926 21146 8927
rect 21118 8793 21146 8794
rect 21118 8767 21119 8793
rect 21119 8767 21145 8793
rect 21145 8767 21146 8793
rect 21118 8766 21146 8767
rect 21118 8633 21146 8634
rect 21118 8607 21119 8633
rect 21119 8607 21145 8633
rect 21145 8607 21146 8633
rect 21118 8606 21146 8607
rect 21118 8473 21146 8474
rect 21118 8447 21119 8473
rect 21119 8447 21145 8473
rect 21145 8447 21146 8473
rect 21118 8446 21146 8447
rect 21118 8313 21146 8314
rect 21118 8287 21119 8313
rect 21119 8287 21145 8313
rect 21145 8287 21146 8313
rect 21118 8286 21146 8287
rect 21118 8153 21146 8154
rect 21118 8127 21119 8153
rect 21119 8127 21145 8153
rect 21145 8127 21146 8153
rect 21118 8126 21146 8127
rect 21118 7993 21146 7994
rect 21118 7967 21119 7993
rect 21119 7967 21145 7993
rect 21145 7967 21146 7993
rect 21118 7966 21146 7967
rect 21118 7833 21146 7834
rect 21118 7807 21119 7833
rect 21119 7807 21145 7833
rect 21145 7807 21146 7833
rect 21118 7806 21146 7807
rect 21118 7673 21146 7674
rect 21118 7647 21119 7673
rect 21119 7647 21145 7673
rect 21145 7647 21146 7673
rect 21118 7646 21146 7647
rect 21118 7513 21146 7514
rect 21118 7487 21119 7513
rect 21119 7487 21145 7513
rect 21145 7487 21146 7513
rect 21118 7486 21146 7487
rect 21118 7353 21146 7354
rect 21118 7327 21119 7353
rect 21119 7327 21145 7353
rect 21145 7327 21146 7353
rect 21118 7326 21146 7327
rect 21118 7193 21146 7194
rect 21118 7167 21119 7193
rect 21119 7167 21145 7193
rect 21145 7167 21146 7193
rect 21118 7166 21146 7167
rect 21118 7033 21146 7034
rect 21118 7007 21119 7033
rect 21119 7007 21145 7033
rect 21145 7007 21146 7033
rect 21118 7006 21146 7007
rect 21118 6873 21146 6874
rect 21118 6847 21119 6873
rect 21119 6847 21145 6873
rect 21145 6847 21146 6873
rect 21118 6846 21146 6847
rect 21118 6713 21146 6714
rect 21118 6687 21119 6713
rect 21119 6687 21145 6713
rect 21145 6687 21146 6713
rect 21118 6686 21146 6687
rect 21118 6553 21146 6554
rect 21118 6527 21119 6553
rect 21119 6527 21145 6553
rect 21145 6527 21146 6553
rect 21118 6526 21146 6527
rect 21118 6393 21146 6394
rect 21118 6367 21119 6393
rect 21119 6367 21145 6393
rect 21145 6367 21146 6393
rect 21118 6366 21146 6367
rect 21118 6233 21146 6234
rect 21118 6207 21119 6233
rect 21119 6207 21145 6233
rect 21145 6207 21146 6233
rect 21118 6206 21146 6207
rect 21118 6073 21146 6074
rect 21118 6047 21119 6073
rect 21119 6047 21145 6073
rect 21145 6047 21146 6073
rect 21118 6046 21146 6047
rect 21118 5913 21146 5914
rect 21118 5887 21119 5913
rect 21119 5887 21145 5913
rect 21145 5887 21146 5913
rect 21118 5886 21146 5887
rect 24851 9113 24879 9114
rect 24851 9087 24852 9113
rect 24852 9087 24878 9113
rect 24878 9087 24879 9113
rect 24851 9086 24879 9087
rect 24851 8953 24879 8954
rect 24851 8927 24852 8953
rect 24852 8927 24878 8953
rect 24878 8927 24879 8953
rect 24851 8926 24879 8927
rect 24851 8793 24879 8794
rect 24851 8767 24852 8793
rect 24852 8767 24878 8793
rect 24878 8767 24879 8793
rect 24851 8766 24879 8767
rect 24851 8633 24879 8634
rect 24851 8607 24852 8633
rect 24852 8607 24878 8633
rect 24878 8607 24879 8633
rect 24851 8606 24879 8607
rect 24851 8473 24879 8474
rect 24851 8447 24852 8473
rect 24852 8447 24878 8473
rect 24878 8447 24879 8473
rect 24851 8446 24879 8447
rect 24851 8313 24879 8314
rect 24851 8287 24852 8313
rect 24852 8287 24878 8313
rect 24878 8287 24879 8313
rect 24851 8286 24879 8287
rect 24851 8153 24879 8154
rect 24851 8127 24852 8153
rect 24852 8127 24878 8153
rect 24878 8127 24879 8153
rect 24851 8126 24879 8127
rect 24851 7993 24879 7994
rect 24851 7967 24852 7993
rect 24852 7967 24878 7993
rect 24878 7967 24879 7993
rect 24851 7966 24879 7967
rect 24851 7833 24879 7834
rect 24851 7807 24852 7833
rect 24852 7807 24878 7833
rect 24878 7807 24879 7833
rect 24851 7806 24879 7807
rect 24851 7673 24879 7674
rect 24851 7647 24852 7673
rect 24852 7647 24878 7673
rect 24878 7647 24879 7673
rect 24851 7646 24879 7647
rect 24851 7513 24879 7514
rect 24851 7487 24852 7513
rect 24852 7487 24878 7513
rect 24878 7487 24879 7513
rect 24851 7486 24879 7487
rect 24851 7353 24879 7354
rect 24851 7327 24852 7353
rect 24852 7327 24878 7353
rect 24878 7327 24879 7353
rect 24851 7326 24879 7327
rect 24851 7193 24879 7194
rect 24851 7167 24852 7193
rect 24852 7167 24878 7193
rect 24878 7167 24879 7193
rect 24851 7166 24879 7167
rect 24851 7033 24879 7034
rect 24851 7007 24852 7033
rect 24852 7007 24878 7033
rect 24878 7007 24879 7033
rect 24851 7006 24879 7007
rect 24851 6873 24879 6874
rect 24851 6847 24852 6873
rect 24852 6847 24878 6873
rect 24878 6847 24879 6873
rect 24851 6846 24879 6847
rect 24851 6713 24879 6714
rect 24851 6687 24852 6713
rect 24852 6687 24878 6713
rect 24878 6687 24879 6713
rect 24851 6686 24879 6687
rect 24851 6553 24879 6554
rect 24851 6527 24852 6553
rect 24852 6527 24878 6553
rect 24878 6527 24879 6553
rect 24851 6526 24879 6527
rect 24851 6393 24879 6394
rect 24851 6367 24852 6393
rect 24852 6367 24878 6393
rect 24878 6367 24879 6393
rect 24851 6366 24879 6367
rect 24851 6233 24879 6234
rect 24851 6207 24852 6233
rect 24852 6207 24878 6233
rect 24878 6207 24879 6233
rect 24851 6206 24879 6207
rect 24851 6073 24879 6074
rect 24851 6047 24852 6073
rect 24852 6047 24878 6073
rect 24878 6047 24879 6073
rect 24851 6046 24879 6047
rect 24851 5913 24879 5914
rect 24851 5887 24852 5913
rect 24852 5887 24878 5913
rect 24878 5887 24879 5913
rect 24851 5886 24879 5887
rect 21118 5753 21146 5754
rect 21118 5727 21119 5753
rect 21119 5727 21145 5753
rect 21145 5727 21146 5753
rect 21118 5726 21146 5727
rect 24851 5753 24879 5754
rect 24851 5727 24852 5753
rect 24852 5727 24878 5753
rect 24878 5727 24879 5753
rect 24851 5726 24879 5727
rect 21306 5650 21334 5651
rect 21306 5624 21307 5650
rect 21307 5624 21333 5650
rect 21333 5624 21334 5650
rect 21306 5623 21334 5624
rect 21466 5650 21494 5651
rect 21466 5624 21467 5650
rect 21467 5624 21493 5650
rect 21493 5624 21494 5650
rect 21466 5623 21494 5624
rect 21626 5650 21654 5651
rect 21626 5624 21627 5650
rect 21627 5624 21653 5650
rect 21653 5624 21654 5650
rect 21626 5623 21654 5624
rect 21786 5650 21814 5651
rect 21786 5624 21787 5650
rect 21787 5624 21813 5650
rect 21813 5624 21814 5650
rect 21786 5623 21814 5624
rect 21946 5650 21974 5651
rect 21946 5624 21947 5650
rect 21947 5624 21973 5650
rect 21973 5624 21974 5650
rect 21946 5623 21974 5624
rect 22106 5650 22134 5651
rect 22106 5624 22107 5650
rect 22107 5624 22133 5650
rect 22133 5624 22134 5650
rect 22106 5623 22134 5624
rect 22266 5650 22294 5651
rect 22266 5624 22267 5650
rect 22267 5624 22293 5650
rect 22293 5624 22294 5650
rect 22266 5623 22294 5624
rect 22426 5650 22454 5651
rect 22426 5624 22427 5650
rect 22427 5624 22453 5650
rect 22453 5624 22454 5650
rect 22426 5623 22454 5624
rect 22586 5650 22614 5651
rect 22586 5624 22587 5650
rect 22587 5624 22613 5650
rect 22613 5624 22614 5650
rect 22586 5623 22614 5624
rect 22746 5650 22774 5651
rect 22746 5624 22747 5650
rect 22747 5624 22773 5650
rect 22773 5624 22774 5650
rect 22746 5623 22774 5624
rect 22906 5650 22934 5651
rect 22906 5624 22907 5650
rect 22907 5624 22933 5650
rect 22933 5624 22934 5650
rect 22906 5623 22934 5624
rect 23066 5650 23094 5651
rect 23066 5624 23067 5650
rect 23067 5624 23093 5650
rect 23093 5624 23094 5650
rect 23066 5623 23094 5624
rect 23226 5650 23254 5651
rect 23226 5624 23227 5650
rect 23227 5624 23253 5650
rect 23253 5624 23254 5650
rect 23226 5623 23254 5624
rect 23386 5650 23414 5651
rect 23386 5624 23387 5650
rect 23387 5624 23413 5650
rect 23413 5624 23414 5650
rect 23386 5623 23414 5624
rect 23546 5650 23574 5651
rect 23546 5624 23547 5650
rect 23547 5624 23573 5650
rect 23573 5624 23574 5650
rect 23546 5623 23574 5624
rect 23706 5650 23734 5651
rect 23706 5624 23707 5650
rect 23707 5624 23733 5650
rect 23733 5624 23734 5650
rect 23706 5623 23734 5624
rect 23866 5650 23894 5651
rect 23866 5624 23867 5650
rect 23867 5624 23893 5650
rect 23893 5624 23894 5650
rect 23866 5623 23894 5624
rect 24026 5650 24054 5651
rect 24026 5624 24027 5650
rect 24027 5624 24053 5650
rect 24053 5624 24054 5650
rect 24026 5623 24054 5624
rect 24186 5650 24214 5651
rect 24186 5624 24187 5650
rect 24187 5624 24213 5650
rect 24213 5624 24214 5650
rect 24186 5623 24214 5624
rect 24346 5650 24374 5651
rect 24346 5624 24347 5650
rect 24347 5624 24373 5650
rect 24373 5624 24374 5650
rect 24346 5623 24374 5624
rect 24506 5650 24534 5651
rect 24506 5624 24507 5650
rect 24507 5624 24533 5650
rect 24533 5624 24534 5650
rect 24506 5623 24534 5624
rect 24666 5650 24694 5651
rect 24666 5624 24667 5650
rect 24667 5624 24693 5650
rect 24693 5624 24694 5650
rect 24666 5623 24694 5624
rect 3306 3378 3334 3379
rect 3306 3352 3307 3378
rect 3307 3352 3333 3378
rect 3333 3352 3334 3378
rect 3306 3351 3334 3352
rect 3466 3378 3494 3379
rect 3466 3352 3467 3378
rect 3467 3352 3493 3378
rect 3493 3352 3494 3378
rect 3466 3351 3494 3352
rect 3626 3378 3654 3379
rect 3626 3352 3627 3378
rect 3627 3352 3653 3378
rect 3653 3352 3654 3378
rect 3626 3351 3654 3352
rect 3786 3378 3814 3379
rect 3786 3352 3787 3378
rect 3787 3352 3813 3378
rect 3813 3352 3814 3378
rect 3786 3351 3814 3352
rect 3946 3378 3974 3379
rect 3946 3352 3947 3378
rect 3947 3352 3973 3378
rect 3973 3352 3974 3378
rect 3946 3351 3974 3352
rect 4106 3378 4134 3379
rect 4106 3352 4107 3378
rect 4107 3352 4133 3378
rect 4133 3352 4134 3378
rect 4106 3351 4134 3352
rect 4266 3378 4294 3379
rect 4266 3352 4267 3378
rect 4267 3352 4293 3378
rect 4293 3352 4294 3378
rect 4266 3351 4294 3352
rect 4426 3378 4454 3379
rect 4426 3352 4427 3378
rect 4427 3352 4453 3378
rect 4453 3352 4454 3378
rect 4426 3351 4454 3352
rect 4586 3378 4614 3379
rect 4586 3352 4587 3378
rect 4587 3352 4613 3378
rect 4613 3352 4614 3378
rect 4586 3351 4614 3352
rect 4746 3378 4774 3379
rect 4746 3352 4747 3378
rect 4747 3352 4773 3378
rect 4773 3352 4774 3378
rect 4746 3351 4774 3352
rect 4906 3378 4934 3379
rect 4906 3352 4907 3378
rect 4907 3352 4933 3378
rect 4933 3352 4934 3378
rect 4906 3351 4934 3352
rect 5066 3378 5094 3379
rect 5066 3352 5067 3378
rect 5067 3352 5093 3378
rect 5093 3352 5094 3378
rect 5066 3351 5094 3352
rect 5226 3378 5254 3379
rect 5226 3352 5227 3378
rect 5227 3352 5253 3378
rect 5253 3352 5254 3378
rect 5226 3351 5254 3352
rect 5386 3378 5414 3379
rect 5386 3352 5387 3378
rect 5387 3352 5413 3378
rect 5413 3352 5414 3378
rect 5386 3351 5414 3352
rect 5546 3378 5574 3379
rect 5546 3352 5547 3378
rect 5547 3352 5573 3378
rect 5573 3352 5574 3378
rect 5546 3351 5574 3352
rect 5706 3378 5734 3379
rect 5706 3352 5707 3378
rect 5707 3352 5733 3378
rect 5733 3352 5734 3378
rect 5706 3351 5734 3352
rect 5866 3378 5894 3379
rect 5866 3352 5867 3378
rect 5867 3352 5893 3378
rect 5893 3352 5894 3378
rect 5866 3351 5894 3352
rect 6026 3378 6054 3379
rect 6026 3352 6027 3378
rect 6027 3352 6053 3378
rect 6053 3352 6054 3378
rect 6026 3351 6054 3352
rect 6186 3378 6214 3379
rect 6186 3352 6187 3378
rect 6187 3352 6213 3378
rect 6213 3352 6214 3378
rect 6186 3351 6214 3352
rect 6346 3378 6374 3379
rect 6346 3352 6347 3378
rect 6347 3352 6373 3378
rect 6373 3352 6374 3378
rect 6346 3351 6374 3352
rect 6506 3378 6534 3379
rect 6506 3352 6507 3378
rect 6507 3352 6533 3378
rect 6533 3352 6534 3378
rect 6506 3351 6534 3352
rect 6666 3378 6694 3379
rect 6666 3352 6667 3378
rect 6667 3352 6693 3378
rect 6693 3352 6694 3378
rect 6666 3351 6694 3352
rect 3118 3273 3146 3274
rect 3118 3247 3119 3273
rect 3119 3247 3145 3273
rect 3145 3247 3146 3273
rect 3118 3246 3146 3247
rect 6851 3273 6879 3274
rect 6851 3247 6852 3273
rect 6852 3247 6878 3273
rect 6878 3247 6879 3273
rect 6851 3246 6879 3247
rect 3118 3113 3146 3114
rect 3118 3087 3119 3113
rect 3119 3087 3145 3113
rect 3145 3087 3146 3113
rect 3118 3086 3146 3087
rect 3118 2953 3146 2954
rect 3118 2927 3119 2953
rect 3119 2927 3145 2953
rect 3145 2927 3146 2953
rect 3118 2926 3146 2927
rect 3118 2793 3146 2794
rect 3118 2767 3119 2793
rect 3119 2767 3145 2793
rect 3145 2767 3146 2793
rect 3118 2766 3146 2767
rect 3118 2633 3146 2634
rect 3118 2607 3119 2633
rect 3119 2607 3145 2633
rect 3145 2607 3146 2633
rect 3118 2606 3146 2607
rect 3118 2473 3146 2474
rect 3118 2447 3119 2473
rect 3119 2447 3145 2473
rect 3145 2447 3146 2473
rect 3118 2446 3146 2447
rect 3118 2313 3146 2314
rect 3118 2287 3119 2313
rect 3119 2287 3145 2313
rect 3145 2287 3146 2313
rect 3118 2286 3146 2287
rect 3118 2153 3146 2154
rect 3118 2127 3119 2153
rect 3119 2127 3145 2153
rect 3145 2127 3146 2153
rect 3118 2126 3146 2127
rect 3118 1993 3146 1994
rect 3118 1967 3119 1993
rect 3119 1967 3145 1993
rect 3145 1967 3146 1993
rect 3118 1966 3146 1967
rect 3118 1833 3146 1834
rect 3118 1807 3119 1833
rect 3119 1807 3145 1833
rect 3145 1807 3146 1833
rect 3118 1806 3146 1807
rect 3118 1673 3146 1674
rect 3118 1647 3119 1673
rect 3119 1647 3145 1673
rect 3145 1647 3146 1673
rect 3118 1646 3146 1647
rect 3118 1513 3146 1514
rect 3118 1487 3119 1513
rect 3119 1487 3145 1513
rect 3145 1487 3146 1513
rect 3118 1486 3146 1487
rect 3118 1353 3146 1354
rect 3118 1327 3119 1353
rect 3119 1327 3145 1353
rect 3145 1327 3146 1353
rect 3118 1326 3146 1327
rect 3118 1193 3146 1194
rect 3118 1167 3119 1193
rect 3119 1167 3145 1193
rect 3145 1167 3146 1193
rect 3118 1166 3146 1167
rect 3118 1033 3146 1034
rect 3118 1007 3119 1033
rect 3119 1007 3145 1033
rect 3145 1007 3146 1033
rect 3118 1006 3146 1007
rect 3118 873 3146 874
rect 3118 847 3119 873
rect 3119 847 3145 873
rect 3145 847 3146 873
rect 3118 846 3146 847
rect 3118 713 3146 714
rect 3118 687 3119 713
rect 3119 687 3145 713
rect 3145 687 3146 713
rect 3118 686 3146 687
rect 3118 553 3146 554
rect 3118 527 3119 553
rect 3119 527 3145 553
rect 3145 527 3146 553
rect 3118 526 3146 527
rect 3118 393 3146 394
rect 3118 367 3119 393
rect 3119 367 3145 393
rect 3145 367 3146 393
rect 3118 366 3146 367
rect 3118 233 3146 234
rect 3118 207 3119 233
rect 3119 207 3145 233
rect 3145 207 3146 233
rect 3118 206 3146 207
rect 3118 73 3146 74
rect 3118 47 3119 73
rect 3119 47 3145 73
rect 3145 47 3146 73
rect 3118 46 3146 47
rect 3118 -87 3146 -86
rect 3118 -113 3119 -87
rect 3119 -113 3145 -87
rect 3145 -113 3146 -87
rect 3118 -114 3146 -113
rect 6851 3113 6879 3114
rect 6851 3087 6852 3113
rect 6852 3087 6878 3113
rect 6878 3087 6879 3113
rect 6851 3086 6879 3087
rect 6851 2953 6879 2954
rect 6851 2927 6852 2953
rect 6852 2927 6878 2953
rect 6878 2927 6879 2953
rect 6851 2926 6879 2927
rect 6851 2793 6879 2794
rect 6851 2767 6852 2793
rect 6852 2767 6878 2793
rect 6878 2767 6879 2793
rect 6851 2766 6879 2767
rect 6851 2633 6879 2634
rect 6851 2607 6852 2633
rect 6852 2607 6878 2633
rect 6878 2607 6879 2633
rect 6851 2606 6879 2607
rect 6851 2473 6879 2474
rect 6851 2447 6852 2473
rect 6852 2447 6878 2473
rect 6878 2447 6879 2473
rect 6851 2446 6879 2447
rect 6851 2313 6879 2314
rect 6851 2287 6852 2313
rect 6852 2287 6878 2313
rect 6878 2287 6879 2313
rect 6851 2286 6879 2287
rect 6851 2153 6879 2154
rect 6851 2127 6852 2153
rect 6852 2127 6878 2153
rect 6878 2127 6879 2153
rect 6851 2126 6879 2127
rect 6851 1993 6879 1994
rect 6851 1967 6852 1993
rect 6852 1967 6878 1993
rect 6878 1967 6879 1993
rect 6851 1966 6879 1967
rect 6851 1833 6879 1834
rect 6851 1807 6852 1833
rect 6852 1807 6878 1833
rect 6878 1807 6879 1833
rect 6851 1806 6879 1807
rect 6851 1673 6879 1674
rect 6851 1647 6852 1673
rect 6852 1647 6878 1673
rect 6878 1647 6879 1673
rect 6851 1646 6879 1647
rect 6851 1513 6879 1514
rect 6851 1487 6852 1513
rect 6852 1487 6878 1513
rect 6878 1487 6879 1513
rect 6851 1486 6879 1487
rect 6851 1353 6879 1354
rect 6851 1327 6852 1353
rect 6852 1327 6878 1353
rect 6878 1327 6879 1353
rect 6851 1326 6879 1327
rect 6851 1193 6879 1194
rect 6851 1167 6852 1193
rect 6852 1167 6878 1193
rect 6878 1167 6879 1193
rect 6851 1166 6879 1167
rect 6851 1033 6879 1034
rect 6851 1007 6852 1033
rect 6852 1007 6878 1033
rect 6878 1007 6879 1033
rect 6851 1006 6879 1007
rect 6851 873 6879 874
rect 6851 847 6852 873
rect 6852 847 6878 873
rect 6878 847 6879 873
rect 6851 846 6879 847
rect 6851 713 6879 714
rect 6851 687 6852 713
rect 6852 687 6878 713
rect 6878 687 6879 713
rect 6851 686 6879 687
rect 6851 553 6879 554
rect 6851 527 6852 553
rect 6852 527 6878 553
rect 6878 527 6879 553
rect 6851 526 6879 527
rect 6851 393 6879 394
rect 6851 367 6852 393
rect 6852 367 6878 393
rect 6878 367 6879 393
rect 6851 366 6879 367
rect 6851 233 6879 234
rect 6851 207 6852 233
rect 6852 207 6878 233
rect 6878 207 6879 233
rect 6851 206 6879 207
rect 6851 73 6879 74
rect 6851 47 6852 73
rect 6852 47 6878 73
rect 6878 47 6879 73
rect 6851 46 6879 47
rect 6851 -87 6879 -86
rect 6851 -113 6852 -87
rect 6852 -113 6878 -87
rect 6878 -113 6879 -87
rect 6851 -114 6879 -113
rect 3118 -247 3146 -246
rect 3118 -273 3119 -247
rect 3119 -273 3145 -247
rect 3145 -273 3146 -247
rect 3118 -274 3146 -273
rect 6851 -247 6879 -246
rect 6851 -273 6852 -247
rect 6852 -273 6878 -247
rect 6878 -273 6879 -247
rect 6851 -274 6879 -273
rect 3306 -350 3334 -349
rect 3306 -376 3307 -350
rect 3307 -376 3333 -350
rect 3333 -376 3334 -350
rect 3306 -377 3334 -376
rect 3466 -350 3494 -349
rect 3466 -376 3467 -350
rect 3467 -376 3493 -350
rect 3493 -376 3494 -350
rect 3466 -377 3494 -376
rect 3626 -350 3654 -349
rect 3626 -376 3627 -350
rect 3627 -376 3653 -350
rect 3653 -376 3654 -350
rect 3626 -377 3654 -376
rect 3786 -350 3814 -349
rect 3786 -376 3787 -350
rect 3787 -376 3813 -350
rect 3813 -376 3814 -350
rect 3786 -377 3814 -376
rect 3946 -350 3974 -349
rect 3946 -376 3947 -350
rect 3947 -376 3973 -350
rect 3973 -376 3974 -350
rect 3946 -377 3974 -376
rect 4106 -350 4134 -349
rect 4106 -376 4107 -350
rect 4107 -376 4133 -350
rect 4133 -376 4134 -350
rect 4106 -377 4134 -376
rect 4266 -350 4294 -349
rect 4266 -376 4267 -350
rect 4267 -376 4293 -350
rect 4293 -376 4294 -350
rect 4266 -377 4294 -376
rect 4426 -350 4454 -349
rect 4426 -376 4427 -350
rect 4427 -376 4453 -350
rect 4453 -376 4454 -350
rect 4426 -377 4454 -376
rect 4586 -350 4614 -349
rect 4586 -376 4587 -350
rect 4587 -376 4613 -350
rect 4613 -376 4614 -350
rect 4586 -377 4614 -376
rect 4746 -350 4774 -349
rect 4746 -376 4747 -350
rect 4747 -376 4773 -350
rect 4773 -376 4774 -350
rect 4746 -377 4774 -376
rect 4906 -350 4934 -349
rect 4906 -376 4907 -350
rect 4907 -376 4933 -350
rect 4933 -376 4934 -350
rect 4906 -377 4934 -376
rect 5066 -350 5094 -349
rect 5066 -376 5067 -350
rect 5067 -376 5093 -350
rect 5093 -376 5094 -350
rect 5066 -377 5094 -376
rect 5226 -350 5254 -349
rect 5226 -376 5227 -350
rect 5227 -376 5253 -350
rect 5253 -376 5254 -350
rect 5226 -377 5254 -376
rect 5386 -350 5414 -349
rect 5386 -376 5387 -350
rect 5387 -376 5413 -350
rect 5413 -376 5414 -350
rect 5386 -377 5414 -376
rect 5546 -350 5574 -349
rect 5546 -376 5547 -350
rect 5547 -376 5573 -350
rect 5573 -376 5574 -350
rect 5546 -377 5574 -376
rect 5706 -350 5734 -349
rect 5706 -376 5707 -350
rect 5707 -376 5733 -350
rect 5733 -376 5734 -350
rect 5706 -377 5734 -376
rect 5866 -350 5894 -349
rect 5866 -376 5867 -350
rect 5867 -376 5893 -350
rect 5893 -376 5894 -350
rect 5866 -377 5894 -376
rect 6026 -350 6054 -349
rect 6026 -376 6027 -350
rect 6027 -376 6053 -350
rect 6053 -376 6054 -350
rect 6026 -377 6054 -376
rect 6186 -350 6214 -349
rect 6186 -376 6187 -350
rect 6187 -376 6213 -350
rect 6213 -376 6214 -350
rect 6186 -377 6214 -376
rect 6346 -350 6374 -349
rect 6346 -376 6347 -350
rect 6347 -376 6373 -350
rect 6373 -376 6374 -350
rect 6346 -377 6374 -376
rect 6506 -350 6534 -349
rect 6506 -376 6507 -350
rect 6507 -376 6533 -350
rect 6533 -376 6534 -350
rect 6506 -377 6534 -376
rect 6666 -350 6694 -349
rect 6666 -376 6667 -350
rect 6667 -376 6693 -350
rect 6693 -376 6694 -350
rect 6666 -377 6694 -376
rect 9306 3378 9334 3379
rect 9306 3352 9307 3378
rect 9307 3352 9333 3378
rect 9333 3352 9334 3378
rect 9306 3351 9334 3352
rect 9466 3378 9494 3379
rect 9466 3352 9467 3378
rect 9467 3352 9493 3378
rect 9493 3352 9494 3378
rect 9466 3351 9494 3352
rect 9626 3378 9654 3379
rect 9626 3352 9627 3378
rect 9627 3352 9653 3378
rect 9653 3352 9654 3378
rect 9626 3351 9654 3352
rect 9786 3378 9814 3379
rect 9786 3352 9787 3378
rect 9787 3352 9813 3378
rect 9813 3352 9814 3378
rect 9786 3351 9814 3352
rect 9946 3378 9974 3379
rect 9946 3352 9947 3378
rect 9947 3352 9973 3378
rect 9973 3352 9974 3378
rect 9946 3351 9974 3352
rect 10106 3378 10134 3379
rect 10106 3352 10107 3378
rect 10107 3352 10133 3378
rect 10133 3352 10134 3378
rect 10106 3351 10134 3352
rect 10266 3378 10294 3379
rect 10266 3352 10267 3378
rect 10267 3352 10293 3378
rect 10293 3352 10294 3378
rect 10266 3351 10294 3352
rect 10426 3378 10454 3379
rect 10426 3352 10427 3378
rect 10427 3352 10453 3378
rect 10453 3352 10454 3378
rect 10426 3351 10454 3352
rect 10586 3378 10614 3379
rect 10586 3352 10587 3378
rect 10587 3352 10613 3378
rect 10613 3352 10614 3378
rect 10586 3351 10614 3352
rect 10746 3378 10774 3379
rect 10746 3352 10747 3378
rect 10747 3352 10773 3378
rect 10773 3352 10774 3378
rect 10746 3351 10774 3352
rect 10906 3378 10934 3379
rect 10906 3352 10907 3378
rect 10907 3352 10933 3378
rect 10933 3352 10934 3378
rect 10906 3351 10934 3352
rect 11066 3378 11094 3379
rect 11066 3352 11067 3378
rect 11067 3352 11093 3378
rect 11093 3352 11094 3378
rect 11066 3351 11094 3352
rect 11226 3378 11254 3379
rect 11226 3352 11227 3378
rect 11227 3352 11253 3378
rect 11253 3352 11254 3378
rect 11226 3351 11254 3352
rect 11386 3378 11414 3379
rect 11386 3352 11387 3378
rect 11387 3352 11413 3378
rect 11413 3352 11414 3378
rect 11386 3351 11414 3352
rect 11546 3378 11574 3379
rect 11546 3352 11547 3378
rect 11547 3352 11573 3378
rect 11573 3352 11574 3378
rect 11546 3351 11574 3352
rect 11706 3378 11734 3379
rect 11706 3352 11707 3378
rect 11707 3352 11733 3378
rect 11733 3352 11734 3378
rect 11706 3351 11734 3352
rect 11866 3378 11894 3379
rect 11866 3352 11867 3378
rect 11867 3352 11893 3378
rect 11893 3352 11894 3378
rect 11866 3351 11894 3352
rect 12026 3378 12054 3379
rect 12026 3352 12027 3378
rect 12027 3352 12053 3378
rect 12053 3352 12054 3378
rect 12026 3351 12054 3352
rect 12186 3378 12214 3379
rect 12186 3352 12187 3378
rect 12187 3352 12213 3378
rect 12213 3352 12214 3378
rect 12186 3351 12214 3352
rect 12346 3378 12374 3379
rect 12346 3352 12347 3378
rect 12347 3352 12373 3378
rect 12373 3352 12374 3378
rect 12346 3351 12374 3352
rect 12506 3378 12534 3379
rect 12506 3352 12507 3378
rect 12507 3352 12533 3378
rect 12533 3352 12534 3378
rect 12506 3351 12534 3352
rect 12666 3378 12694 3379
rect 12666 3352 12667 3378
rect 12667 3352 12693 3378
rect 12693 3352 12694 3378
rect 12666 3351 12694 3352
rect 9118 3273 9146 3274
rect 9118 3247 9119 3273
rect 9119 3247 9145 3273
rect 9145 3247 9146 3273
rect 9118 3246 9146 3247
rect 12851 3273 12879 3274
rect 12851 3247 12852 3273
rect 12852 3247 12878 3273
rect 12878 3247 12879 3273
rect 12851 3246 12879 3247
rect 9118 3113 9146 3114
rect 9118 3087 9119 3113
rect 9119 3087 9145 3113
rect 9145 3087 9146 3113
rect 9118 3086 9146 3087
rect 9118 2953 9146 2954
rect 9118 2927 9119 2953
rect 9119 2927 9145 2953
rect 9145 2927 9146 2953
rect 9118 2926 9146 2927
rect 9118 2793 9146 2794
rect 9118 2767 9119 2793
rect 9119 2767 9145 2793
rect 9145 2767 9146 2793
rect 9118 2766 9146 2767
rect 9118 2633 9146 2634
rect 9118 2607 9119 2633
rect 9119 2607 9145 2633
rect 9145 2607 9146 2633
rect 9118 2606 9146 2607
rect 9118 2473 9146 2474
rect 9118 2447 9119 2473
rect 9119 2447 9145 2473
rect 9145 2447 9146 2473
rect 9118 2446 9146 2447
rect 9118 2313 9146 2314
rect 9118 2287 9119 2313
rect 9119 2287 9145 2313
rect 9145 2287 9146 2313
rect 9118 2286 9146 2287
rect 9118 2153 9146 2154
rect 9118 2127 9119 2153
rect 9119 2127 9145 2153
rect 9145 2127 9146 2153
rect 9118 2126 9146 2127
rect 9118 1993 9146 1994
rect 9118 1967 9119 1993
rect 9119 1967 9145 1993
rect 9145 1967 9146 1993
rect 9118 1966 9146 1967
rect 9118 1833 9146 1834
rect 9118 1807 9119 1833
rect 9119 1807 9145 1833
rect 9145 1807 9146 1833
rect 9118 1806 9146 1807
rect 9118 1673 9146 1674
rect 9118 1647 9119 1673
rect 9119 1647 9145 1673
rect 9145 1647 9146 1673
rect 9118 1646 9146 1647
rect 9118 1513 9146 1514
rect 9118 1487 9119 1513
rect 9119 1487 9145 1513
rect 9145 1487 9146 1513
rect 9118 1486 9146 1487
rect 9118 1353 9146 1354
rect 9118 1327 9119 1353
rect 9119 1327 9145 1353
rect 9145 1327 9146 1353
rect 9118 1326 9146 1327
rect 9118 1193 9146 1194
rect 9118 1167 9119 1193
rect 9119 1167 9145 1193
rect 9145 1167 9146 1193
rect 9118 1166 9146 1167
rect 9118 1033 9146 1034
rect 9118 1007 9119 1033
rect 9119 1007 9145 1033
rect 9145 1007 9146 1033
rect 9118 1006 9146 1007
rect 9118 873 9146 874
rect 9118 847 9119 873
rect 9119 847 9145 873
rect 9145 847 9146 873
rect 9118 846 9146 847
rect 9118 713 9146 714
rect 9118 687 9119 713
rect 9119 687 9145 713
rect 9145 687 9146 713
rect 9118 686 9146 687
rect 9118 553 9146 554
rect 9118 527 9119 553
rect 9119 527 9145 553
rect 9145 527 9146 553
rect 9118 526 9146 527
rect 9118 393 9146 394
rect 9118 367 9119 393
rect 9119 367 9145 393
rect 9145 367 9146 393
rect 9118 366 9146 367
rect 9118 233 9146 234
rect 9118 207 9119 233
rect 9119 207 9145 233
rect 9145 207 9146 233
rect 9118 206 9146 207
rect 9118 73 9146 74
rect 9118 47 9119 73
rect 9119 47 9145 73
rect 9145 47 9146 73
rect 9118 46 9146 47
rect 9118 -87 9146 -86
rect 9118 -113 9119 -87
rect 9119 -113 9145 -87
rect 9145 -113 9146 -87
rect 9118 -114 9146 -113
rect 12851 3113 12879 3114
rect 12851 3087 12852 3113
rect 12852 3087 12878 3113
rect 12878 3087 12879 3113
rect 12851 3086 12879 3087
rect 12851 2953 12879 2954
rect 12851 2927 12852 2953
rect 12852 2927 12878 2953
rect 12878 2927 12879 2953
rect 12851 2926 12879 2927
rect 12851 2793 12879 2794
rect 12851 2767 12852 2793
rect 12852 2767 12878 2793
rect 12878 2767 12879 2793
rect 12851 2766 12879 2767
rect 12851 2633 12879 2634
rect 12851 2607 12852 2633
rect 12852 2607 12878 2633
rect 12878 2607 12879 2633
rect 12851 2606 12879 2607
rect 12851 2473 12879 2474
rect 12851 2447 12852 2473
rect 12852 2447 12878 2473
rect 12878 2447 12879 2473
rect 12851 2446 12879 2447
rect 12851 2313 12879 2314
rect 12851 2287 12852 2313
rect 12852 2287 12878 2313
rect 12878 2287 12879 2313
rect 12851 2286 12879 2287
rect 12851 2153 12879 2154
rect 12851 2127 12852 2153
rect 12852 2127 12878 2153
rect 12878 2127 12879 2153
rect 12851 2126 12879 2127
rect 12851 1993 12879 1994
rect 12851 1967 12852 1993
rect 12852 1967 12878 1993
rect 12878 1967 12879 1993
rect 12851 1966 12879 1967
rect 12851 1833 12879 1834
rect 12851 1807 12852 1833
rect 12852 1807 12878 1833
rect 12878 1807 12879 1833
rect 12851 1806 12879 1807
rect 12851 1673 12879 1674
rect 12851 1647 12852 1673
rect 12852 1647 12878 1673
rect 12878 1647 12879 1673
rect 12851 1646 12879 1647
rect 12851 1513 12879 1514
rect 12851 1487 12852 1513
rect 12852 1487 12878 1513
rect 12878 1487 12879 1513
rect 12851 1486 12879 1487
rect 12851 1353 12879 1354
rect 12851 1327 12852 1353
rect 12852 1327 12878 1353
rect 12878 1327 12879 1353
rect 12851 1326 12879 1327
rect 12851 1193 12879 1194
rect 12851 1167 12852 1193
rect 12852 1167 12878 1193
rect 12878 1167 12879 1193
rect 12851 1166 12879 1167
rect 12851 1033 12879 1034
rect 12851 1007 12852 1033
rect 12852 1007 12878 1033
rect 12878 1007 12879 1033
rect 12851 1006 12879 1007
rect 12851 873 12879 874
rect 12851 847 12852 873
rect 12852 847 12878 873
rect 12878 847 12879 873
rect 12851 846 12879 847
rect 12851 713 12879 714
rect 12851 687 12852 713
rect 12852 687 12878 713
rect 12878 687 12879 713
rect 12851 686 12879 687
rect 12851 553 12879 554
rect 12851 527 12852 553
rect 12852 527 12878 553
rect 12878 527 12879 553
rect 12851 526 12879 527
rect 12851 393 12879 394
rect 12851 367 12852 393
rect 12852 367 12878 393
rect 12878 367 12879 393
rect 12851 366 12879 367
rect 12851 233 12879 234
rect 12851 207 12852 233
rect 12852 207 12878 233
rect 12878 207 12879 233
rect 12851 206 12879 207
rect 12851 73 12879 74
rect 12851 47 12852 73
rect 12852 47 12878 73
rect 12878 47 12879 73
rect 12851 46 12879 47
rect 12851 -87 12879 -86
rect 12851 -113 12852 -87
rect 12852 -113 12878 -87
rect 12878 -113 12879 -87
rect 12851 -114 12879 -113
rect 9118 -247 9146 -246
rect 9118 -273 9119 -247
rect 9119 -273 9145 -247
rect 9145 -273 9146 -247
rect 9118 -274 9146 -273
rect 12851 -247 12879 -246
rect 12851 -273 12852 -247
rect 12852 -273 12878 -247
rect 12878 -273 12879 -247
rect 12851 -274 12879 -273
rect 9306 -350 9334 -349
rect 9306 -376 9307 -350
rect 9307 -376 9333 -350
rect 9333 -376 9334 -350
rect 9306 -377 9334 -376
rect 9466 -350 9494 -349
rect 9466 -376 9467 -350
rect 9467 -376 9493 -350
rect 9493 -376 9494 -350
rect 9466 -377 9494 -376
rect 9626 -350 9654 -349
rect 9626 -376 9627 -350
rect 9627 -376 9653 -350
rect 9653 -376 9654 -350
rect 9626 -377 9654 -376
rect 9786 -350 9814 -349
rect 9786 -376 9787 -350
rect 9787 -376 9813 -350
rect 9813 -376 9814 -350
rect 9786 -377 9814 -376
rect 9946 -350 9974 -349
rect 9946 -376 9947 -350
rect 9947 -376 9973 -350
rect 9973 -376 9974 -350
rect 9946 -377 9974 -376
rect 10106 -350 10134 -349
rect 10106 -376 10107 -350
rect 10107 -376 10133 -350
rect 10133 -376 10134 -350
rect 10106 -377 10134 -376
rect 10266 -350 10294 -349
rect 10266 -376 10267 -350
rect 10267 -376 10293 -350
rect 10293 -376 10294 -350
rect 10266 -377 10294 -376
rect 10426 -350 10454 -349
rect 10426 -376 10427 -350
rect 10427 -376 10453 -350
rect 10453 -376 10454 -350
rect 10426 -377 10454 -376
rect 10586 -350 10614 -349
rect 10586 -376 10587 -350
rect 10587 -376 10613 -350
rect 10613 -376 10614 -350
rect 10586 -377 10614 -376
rect 10746 -350 10774 -349
rect 10746 -376 10747 -350
rect 10747 -376 10773 -350
rect 10773 -376 10774 -350
rect 10746 -377 10774 -376
rect 10906 -350 10934 -349
rect 10906 -376 10907 -350
rect 10907 -376 10933 -350
rect 10933 -376 10934 -350
rect 10906 -377 10934 -376
rect 11066 -350 11094 -349
rect 11066 -376 11067 -350
rect 11067 -376 11093 -350
rect 11093 -376 11094 -350
rect 11066 -377 11094 -376
rect 11226 -350 11254 -349
rect 11226 -376 11227 -350
rect 11227 -376 11253 -350
rect 11253 -376 11254 -350
rect 11226 -377 11254 -376
rect 11386 -350 11414 -349
rect 11386 -376 11387 -350
rect 11387 -376 11413 -350
rect 11413 -376 11414 -350
rect 11386 -377 11414 -376
rect 11546 -350 11574 -349
rect 11546 -376 11547 -350
rect 11547 -376 11573 -350
rect 11573 -376 11574 -350
rect 11546 -377 11574 -376
rect 11706 -350 11734 -349
rect 11706 -376 11707 -350
rect 11707 -376 11733 -350
rect 11733 -376 11734 -350
rect 11706 -377 11734 -376
rect 11866 -350 11894 -349
rect 11866 -376 11867 -350
rect 11867 -376 11893 -350
rect 11893 -376 11894 -350
rect 11866 -377 11894 -376
rect 12026 -350 12054 -349
rect 12026 -376 12027 -350
rect 12027 -376 12053 -350
rect 12053 -376 12054 -350
rect 12026 -377 12054 -376
rect 12186 -350 12214 -349
rect 12186 -376 12187 -350
rect 12187 -376 12213 -350
rect 12213 -376 12214 -350
rect 12186 -377 12214 -376
rect 12346 -350 12374 -349
rect 12346 -376 12347 -350
rect 12347 -376 12373 -350
rect 12373 -376 12374 -350
rect 12346 -377 12374 -376
rect 12506 -350 12534 -349
rect 12506 -376 12507 -350
rect 12507 -376 12533 -350
rect 12533 -376 12534 -350
rect 12506 -377 12534 -376
rect 12666 -350 12694 -349
rect 12666 -376 12667 -350
rect 12667 -376 12693 -350
rect 12693 -376 12694 -350
rect 12666 -377 12694 -376
rect 15306 3378 15334 3379
rect 15306 3352 15307 3378
rect 15307 3352 15333 3378
rect 15333 3352 15334 3378
rect 15306 3351 15334 3352
rect 15466 3378 15494 3379
rect 15466 3352 15467 3378
rect 15467 3352 15493 3378
rect 15493 3352 15494 3378
rect 15466 3351 15494 3352
rect 15626 3378 15654 3379
rect 15626 3352 15627 3378
rect 15627 3352 15653 3378
rect 15653 3352 15654 3378
rect 15626 3351 15654 3352
rect 15786 3378 15814 3379
rect 15786 3352 15787 3378
rect 15787 3352 15813 3378
rect 15813 3352 15814 3378
rect 15786 3351 15814 3352
rect 15946 3378 15974 3379
rect 15946 3352 15947 3378
rect 15947 3352 15973 3378
rect 15973 3352 15974 3378
rect 15946 3351 15974 3352
rect 16106 3378 16134 3379
rect 16106 3352 16107 3378
rect 16107 3352 16133 3378
rect 16133 3352 16134 3378
rect 16106 3351 16134 3352
rect 16266 3378 16294 3379
rect 16266 3352 16267 3378
rect 16267 3352 16293 3378
rect 16293 3352 16294 3378
rect 16266 3351 16294 3352
rect 16426 3378 16454 3379
rect 16426 3352 16427 3378
rect 16427 3352 16453 3378
rect 16453 3352 16454 3378
rect 16426 3351 16454 3352
rect 16586 3378 16614 3379
rect 16586 3352 16587 3378
rect 16587 3352 16613 3378
rect 16613 3352 16614 3378
rect 16586 3351 16614 3352
rect 16746 3378 16774 3379
rect 16746 3352 16747 3378
rect 16747 3352 16773 3378
rect 16773 3352 16774 3378
rect 16746 3351 16774 3352
rect 16906 3378 16934 3379
rect 16906 3352 16907 3378
rect 16907 3352 16933 3378
rect 16933 3352 16934 3378
rect 16906 3351 16934 3352
rect 17066 3378 17094 3379
rect 17066 3352 17067 3378
rect 17067 3352 17093 3378
rect 17093 3352 17094 3378
rect 17066 3351 17094 3352
rect 17226 3378 17254 3379
rect 17226 3352 17227 3378
rect 17227 3352 17253 3378
rect 17253 3352 17254 3378
rect 17226 3351 17254 3352
rect 17386 3378 17414 3379
rect 17386 3352 17387 3378
rect 17387 3352 17413 3378
rect 17413 3352 17414 3378
rect 17386 3351 17414 3352
rect 17546 3378 17574 3379
rect 17546 3352 17547 3378
rect 17547 3352 17573 3378
rect 17573 3352 17574 3378
rect 17546 3351 17574 3352
rect 17706 3378 17734 3379
rect 17706 3352 17707 3378
rect 17707 3352 17733 3378
rect 17733 3352 17734 3378
rect 17706 3351 17734 3352
rect 17866 3378 17894 3379
rect 17866 3352 17867 3378
rect 17867 3352 17893 3378
rect 17893 3352 17894 3378
rect 17866 3351 17894 3352
rect 18026 3378 18054 3379
rect 18026 3352 18027 3378
rect 18027 3352 18053 3378
rect 18053 3352 18054 3378
rect 18026 3351 18054 3352
rect 18186 3378 18214 3379
rect 18186 3352 18187 3378
rect 18187 3352 18213 3378
rect 18213 3352 18214 3378
rect 18186 3351 18214 3352
rect 18346 3378 18374 3379
rect 18346 3352 18347 3378
rect 18347 3352 18373 3378
rect 18373 3352 18374 3378
rect 18346 3351 18374 3352
rect 18506 3378 18534 3379
rect 18506 3352 18507 3378
rect 18507 3352 18533 3378
rect 18533 3352 18534 3378
rect 18506 3351 18534 3352
rect 18666 3378 18694 3379
rect 18666 3352 18667 3378
rect 18667 3352 18693 3378
rect 18693 3352 18694 3378
rect 18666 3351 18694 3352
rect 15118 3273 15146 3274
rect 15118 3247 15119 3273
rect 15119 3247 15145 3273
rect 15145 3247 15146 3273
rect 15118 3246 15146 3247
rect 18851 3273 18879 3274
rect 18851 3247 18852 3273
rect 18852 3247 18878 3273
rect 18878 3247 18879 3273
rect 18851 3246 18879 3247
rect 15118 3113 15146 3114
rect 15118 3087 15119 3113
rect 15119 3087 15145 3113
rect 15145 3087 15146 3113
rect 15118 3086 15146 3087
rect 15118 2953 15146 2954
rect 15118 2927 15119 2953
rect 15119 2927 15145 2953
rect 15145 2927 15146 2953
rect 15118 2926 15146 2927
rect 15118 2793 15146 2794
rect 15118 2767 15119 2793
rect 15119 2767 15145 2793
rect 15145 2767 15146 2793
rect 15118 2766 15146 2767
rect 15118 2633 15146 2634
rect 15118 2607 15119 2633
rect 15119 2607 15145 2633
rect 15145 2607 15146 2633
rect 15118 2606 15146 2607
rect 15118 2473 15146 2474
rect 15118 2447 15119 2473
rect 15119 2447 15145 2473
rect 15145 2447 15146 2473
rect 15118 2446 15146 2447
rect 15118 2313 15146 2314
rect 15118 2287 15119 2313
rect 15119 2287 15145 2313
rect 15145 2287 15146 2313
rect 15118 2286 15146 2287
rect 15118 2153 15146 2154
rect 15118 2127 15119 2153
rect 15119 2127 15145 2153
rect 15145 2127 15146 2153
rect 15118 2126 15146 2127
rect 15118 1993 15146 1994
rect 15118 1967 15119 1993
rect 15119 1967 15145 1993
rect 15145 1967 15146 1993
rect 15118 1966 15146 1967
rect 15118 1833 15146 1834
rect 15118 1807 15119 1833
rect 15119 1807 15145 1833
rect 15145 1807 15146 1833
rect 15118 1806 15146 1807
rect 15118 1673 15146 1674
rect 15118 1647 15119 1673
rect 15119 1647 15145 1673
rect 15145 1647 15146 1673
rect 15118 1646 15146 1647
rect 15118 1513 15146 1514
rect 15118 1487 15119 1513
rect 15119 1487 15145 1513
rect 15145 1487 15146 1513
rect 15118 1486 15146 1487
rect 15118 1353 15146 1354
rect 15118 1327 15119 1353
rect 15119 1327 15145 1353
rect 15145 1327 15146 1353
rect 15118 1326 15146 1327
rect 15118 1193 15146 1194
rect 15118 1167 15119 1193
rect 15119 1167 15145 1193
rect 15145 1167 15146 1193
rect 15118 1166 15146 1167
rect 15118 1033 15146 1034
rect 15118 1007 15119 1033
rect 15119 1007 15145 1033
rect 15145 1007 15146 1033
rect 15118 1006 15146 1007
rect 15118 873 15146 874
rect 15118 847 15119 873
rect 15119 847 15145 873
rect 15145 847 15146 873
rect 15118 846 15146 847
rect 15118 713 15146 714
rect 15118 687 15119 713
rect 15119 687 15145 713
rect 15145 687 15146 713
rect 15118 686 15146 687
rect 15118 553 15146 554
rect 15118 527 15119 553
rect 15119 527 15145 553
rect 15145 527 15146 553
rect 15118 526 15146 527
rect 15118 393 15146 394
rect 15118 367 15119 393
rect 15119 367 15145 393
rect 15145 367 15146 393
rect 15118 366 15146 367
rect 15118 233 15146 234
rect 15118 207 15119 233
rect 15119 207 15145 233
rect 15145 207 15146 233
rect 15118 206 15146 207
rect 15118 73 15146 74
rect 15118 47 15119 73
rect 15119 47 15145 73
rect 15145 47 15146 73
rect 15118 46 15146 47
rect 15118 -87 15146 -86
rect 15118 -113 15119 -87
rect 15119 -113 15145 -87
rect 15145 -113 15146 -87
rect 15118 -114 15146 -113
rect 18851 3113 18879 3114
rect 18851 3087 18852 3113
rect 18852 3087 18878 3113
rect 18878 3087 18879 3113
rect 18851 3086 18879 3087
rect 18851 2953 18879 2954
rect 18851 2927 18852 2953
rect 18852 2927 18878 2953
rect 18878 2927 18879 2953
rect 18851 2926 18879 2927
rect 18851 2793 18879 2794
rect 18851 2767 18852 2793
rect 18852 2767 18878 2793
rect 18878 2767 18879 2793
rect 18851 2766 18879 2767
rect 18851 2633 18879 2634
rect 18851 2607 18852 2633
rect 18852 2607 18878 2633
rect 18878 2607 18879 2633
rect 18851 2606 18879 2607
rect 18851 2473 18879 2474
rect 18851 2447 18852 2473
rect 18852 2447 18878 2473
rect 18878 2447 18879 2473
rect 18851 2446 18879 2447
rect 18851 2313 18879 2314
rect 18851 2287 18852 2313
rect 18852 2287 18878 2313
rect 18878 2287 18879 2313
rect 18851 2286 18879 2287
rect 18851 2153 18879 2154
rect 18851 2127 18852 2153
rect 18852 2127 18878 2153
rect 18878 2127 18879 2153
rect 18851 2126 18879 2127
rect 18851 1993 18879 1994
rect 18851 1967 18852 1993
rect 18852 1967 18878 1993
rect 18878 1967 18879 1993
rect 18851 1966 18879 1967
rect 18851 1833 18879 1834
rect 18851 1807 18852 1833
rect 18852 1807 18878 1833
rect 18878 1807 18879 1833
rect 18851 1806 18879 1807
rect 18851 1673 18879 1674
rect 18851 1647 18852 1673
rect 18852 1647 18878 1673
rect 18878 1647 18879 1673
rect 18851 1646 18879 1647
rect 18851 1513 18879 1514
rect 18851 1487 18852 1513
rect 18852 1487 18878 1513
rect 18878 1487 18879 1513
rect 18851 1486 18879 1487
rect 18851 1353 18879 1354
rect 18851 1327 18852 1353
rect 18852 1327 18878 1353
rect 18878 1327 18879 1353
rect 18851 1326 18879 1327
rect 18851 1193 18879 1194
rect 18851 1167 18852 1193
rect 18852 1167 18878 1193
rect 18878 1167 18879 1193
rect 18851 1166 18879 1167
rect 18851 1033 18879 1034
rect 18851 1007 18852 1033
rect 18852 1007 18878 1033
rect 18878 1007 18879 1033
rect 18851 1006 18879 1007
rect 18851 873 18879 874
rect 18851 847 18852 873
rect 18852 847 18878 873
rect 18878 847 18879 873
rect 18851 846 18879 847
rect 18851 713 18879 714
rect 18851 687 18852 713
rect 18852 687 18878 713
rect 18878 687 18879 713
rect 18851 686 18879 687
rect 18851 553 18879 554
rect 18851 527 18852 553
rect 18852 527 18878 553
rect 18878 527 18879 553
rect 18851 526 18879 527
rect 18851 393 18879 394
rect 18851 367 18852 393
rect 18852 367 18878 393
rect 18878 367 18879 393
rect 18851 366 18879 367
rect 18851 233 18879 234
rect 18851 207 18852 233
rect 18852 207 18878 233
rect 18878 207 18879 233
rect 18851 206 18879 207
rect 18851 73 18879 74
rect 18851 47 18852 73
rect 18852 47 18878 73
rect 18878 47 18879 73
rect 18851 46 18879 47
rect 18851 -87 18879 -86
rect 18851 -113 18852 -87
rect 18852 -113 18878 -87
rect 18878 -113 18879 -87
rect 18851 -114 18879 -113
rect 15118 -247 15146 -246
rect 15118 -273 15119 -247
rect 15119 -273 15145 -247
rect 15145 -273 15146 -247
rect 15118 -274 15146 -273
rect 18851 -247 18879 -246
rect 18851 -273 18852 -247
rect 18852 -273 18878 -247
rect 18878 -273 18879 -247
rect 18851 -274 18879 -273
rect 21306 3378 21334 3379
rect 21306 3352 21307 3378
rect 21307 3352 21333 3378
rect 21333 3352 21334 3378
rect 21306 3351 21334 3352
rect 21466 3378 21494 3379
rect 21466 3352 21467 3378
rect 21467 3352 21493 3378
rect 21493 3352 21494 3378
rect 21466 3351 21494 3352
rect 21626 3378 21654 3379
rect 21626 3352 21627 3378
rect 21627 3352 21653 3378
rect 21653 3352 21654 3378
rect 21626 3351 21654 3352
rect 21786 3378 21814 3379
rect 21786 3352 21787 3378
rect 21787 3352 21813 3378
rect 21813 3352 21814 3378
rect 21786 3351 21814 3352
rect 21946 3378 21974 3379
rect 21946 3352 21947 3378
rect 21947 3352 21973 3378
rect 21973 3352 21974 3378
rect 21946 3351 21974 3352
rect 22106 3378 22134 3379
rect 22106 3352 22107 3378
rect 22107 3352 22133 3378
rect 22133 3352 22134 3378
rect 22106 3351 22134 3352
rect 22266 3378 22294 3379
rect 22266 3352 22267 3378
rect 22267 3352 22293 3378
rect 22293 3352 22294 3378
rect 22266 3351 22294 3352
rect 22426 3378 22454 3379
rect 22426 3352 22427 3378
rect 22427 3352 22453 3378
rect 22453 3352 22454 3378
rect 22426 3351 22454 3352
rect 22586 3378 22614 3379
rect 22586 3352 22587 3378
rect 22587 3352 22613 3378
rect 22613 3352 22614 3378
rect 22586 3351 22614 3352
rect 22746 3378 22774 3379
rect 22746 3352 22747 3378
rect 22747 3352 22773 3378
rect 22773 3352 22774 3378
rect 22746 3351 22774 3352
rect 22906 3378 22934 3379
rect 22906 3352 22907 3378
rect 22907 3352 22933 3378
rect 22933 3352 22934 3378
rect 22906 3351 22934 3352
rect 23066 3378 23094 3379
rect 23066 3352 23067 3378
rect 23067 3352 23093 3378
rect 23093 3352 23094 3378
rect 23066 3351 23094 3352
rect 23226 3378 23254 3379
rect 23226 3352 23227 3378
rect 23227 3352 23253 3378
rect 23253 3352 23254 3378
rect 23226 3351 23254 3352
rect 23386 3378 23414 3379
rect 23386 3352 23387 3378
rect 23387 3352 23413 3378
rect 23413 3352 23414 3378
rect 23386 3351 23414 3352
rect 23546 3378 23574 3379
rect 23546 3352 23547 3378
rect 23547 3352 23573 3378
rect 23573 3352 23574 3378
rect 23546 3351 23574 3352
rect 23706 3378 23734 3379
rect 23706 3352 23707 3378
rect 23707 3352 23733 3378
rect 23733 3352 23734 3378
rect 23706 3351 23734 3352
rect 23866 3378 23894 3379
rect 23866 3352 23867 3378
rect 23867 3352 23893 3378
rect 23893 3352 23894 3378
rect 23866 3351 23894 3352
rect 24026 3378 24054 3379
rect 24026 3352 24027 3378
rect 24027 3352 24053 3378
rect 24053 3352 24054 3378
rect 24026 3351 24054 3352
rect 24186 3378 24214 3379
rect 24186 3352 24187 3378
rect 24187 3352 24213 3378
rect 24213 3352 24214 3378
rect 24186 3351 24214 3352
rect 24346 3378 24374 3379
rect 24346 3352 24347 3378
rect 24347 3352 24373 3378
rect 24373 3352 24374 3378
rect 24346 3351 24374 3352
rect 24506 3378 24534 3379
rect 24506 3352 24507 3378
rect 24507 3352 24533 3378
rect 24533 3352 24534 3378
rect 24506 3351 24534 3352
rect 24666 3378 24694 3379
rect 24666 3352 24667 3378
rect 24667 3352 24693 3378
rect 24693 3352 24694 3378
rect 24666 3351 24694 3352
rect 21118 3273 21146 3274
rect 21118 3247 21119 3273
rect 21119 3247 21145 3273
rect 21145 3247 21146 3273
rect 21118 3246 21146 3247
rect 24851 3273 24879 3274
rect 24851 3247 24852 3273
rect 24852 3247 24878 3273
rect 24878 3247 24879 3273
rect 24851 3246 24879 3247
rect 21118 3113 21146 3114
rect 21118 3087 21119 3113
rect 21119 3087 21145 3113
rect 21145 3087 21146 3113
rect 21118 3086 21146 3087
rect 21118 2953 21146 2954
rect 21118 2927 21119 2953
rect 21119 2927 21145 2953
rect 21145 2927 21146 2953
rect 21118 2926 21146 2927
rect 21118 2793 21146 2794
rect 21118 2767 21119 2793
rect 21119 2767 21145 2793
rect 21145 2767 21146 2793
rect 21118 2766 21146 2767
rect 21118 2633 21146 2634
rect 21118 2607 21119 2633
rect 21119 2607 21145 2633
rect 21145 2607 21146 2633
rect 21118 2606 21146 2607
rect 21118 2473 21146 2474
rect 21118 2447 21119 2473
rect 21119 2447 21145 2473
rect 21145 2447 21146 2473
rect 21118 2446 21146 2447
rect 21118 2313 21146 2314
rect 21118 2287 21119 2313
rect 21119 2287 21145 2313
rect 21145 2287 21146 2313
rect 21118 2286 21146 2287
rect 21118 2153 21146 2154
rect 21118 2127 21119 2153
rect 21119 2127 21145 2153
rect 21145 2127 21146 2153
rect 21118 2126 21146 2127
rect 21118 1993 21146 1994
rect 21118 1967 21119 1993
rect 21119 1967 21145 1993
rect 21145 1967 21146 1993
rect 21118 1966 21146 1967
rect 21118 1833 21146 1834
rect 21118 1807 21119 1833
rect 21119 1807 21145 1833
rect 21145 1807 21146 1833
rect 21118 1806 21146 1807
rect 21118 1673 21146 1674
rect 21118 1647 21119 1673
rect 21119 1647 21145 1673
rect 21145 1647 21146 1673
rect 21118 1646 21146 1647
rect 21118 1513 21146 1514
rect 21118 1487 21119 1513
rect 21119 1487 21145 1513
rect 21145 1487 21146 1513
rect 21118 1486 21146 1487
rect 21118 1353 21146 1354
rect 21118 1327 21119 1353
rect 21119 1327 21145 1353
rect 21145 1327 21146 1353
rect 21118 1326 21146 1327
rect 21118 1193 21146 1194
rect 21118 1167 21119 1193
rect 21119 1167 21145 1193
rect 21145 1167 21146 1193
rect 21118 1166 21146 1167
rect 21118 1033 21146 1034
rect 21118 1007 21119 1033
rect 21119 1007 21145 1033
rect 21145 1007 21146 1033
rect 21118 1006 21146 1007
rect 21118 873 21146 874
rect 21118 847 21119 873
rect 21119 847 21145 873
rect 21145 847 21146 873
rect 21118 846 21146 847
rect 21118 713 21146 714
rect 21118 687 21119 713
rect 21119 687 21145 713
rect 21145 687 21146 713
rect 21118 686 21146 687
rect 21118 553 21146 554
rect 21118 527 21119 553
rect 21119 527 21145 553
rect 21145 527 21146 553
rect 21118 526 21146 527
rect 21118 393 21146 394
rect 21118 367 21119 393
rect 21119 367 21145 393
rect 21145 367 21146 393
rect 21118 366 21146 367
rect 21118 233 21146 234
rect 21118 207 21119 233
rect 21119 207 21145 233
rect 21145 207 21146 233
rect 21118 206 21146 207
rect 21118 73 21146 74
rect 21118 47 21119 73
rect 21119 47 21145 73
rect 21145 47 21146 73
rect 21118 46 21146 47
rect 21118 -87 21146 -86
rect 21118 -113 21119 -87
rect 21119 -113 21145 -87
rect 21145 -113 21146 -87
rect 21118 -114 21146 -113
rect 24851 3113 24879 3114
rect 24851 3087 24852 3113
rect 24852 3087 24878 3113
rect 24878 3087 24879 3113
rect 24851 3086 24879 3087
rect 24851 2953 24879 2954
rect 24851 2927 24852 2953
rect 24852 2927 24878 2953
rect 24878 2927 24879 2953
rect 24851 2926 24879 2927
rect 24851 2793 24879 2794
rect 24851 2767 24852 2793
rect 24852 2767 24878 2793
rect 24878 2767 24879 2793
rect 24851 2766 24879 2767
rect 24851 2633 24879 2634
rect 24851 2607 24852 2633
rect 24852 2607 24878 2633
rect 24878 2607 24879 2633
rect 24851 2606 24879 2607
rect 24851 2473 24879 2474
rect 24851 2447 24852 2473
rect 24852 2447 24878 2473
rect 24878 2447 24879 2473
rect 24851 2446 24879 2447
rect 24851 2313 24879 2314
rect 24851 2287 24852 2313
rect 24852 2287 24878 2313
rect 24878 2287 24879 2313
rect 24851 2286 24879 2287
rect 24851 2153 24879 2154
rect 24851 2127 24852 2153
rect 24852 2127 24878 2153
rect 24878 2127 24879 2153
rect 24851 2126 24879 2127
rect 24851 1993 24879 1994
rect 24851 1967 24852 1993
rect 24852 1967 24878 1993
rect 24878 1967 24879 1993
rect 24851 1966 24879 1967
rect 24851 1833 24879 1834
rect 24851 1807 24852 1833
rect 24852 1807 24878 1833
rect 24878 1807 24879 1833
rect 24851 1806 24879 1807
rect 24851 1673 24879 1674
rect 24851 1647 24852 1673
rect 24852 1647 24878 1673
rect 24878 1647 24879 1673
rect 24851 1646 24879 1647
rect 24851 1513 24879 1514
rect 24851 1487 24852 1513
rect 24852 1487 24878 1513
rect 24878 1487 24879 1513
rect 24851 1486 24879 1487
rect 24851 1353 24879 1354
rect 24851 1327 24852 1353
rect 24852 1327 24878 1353
rect 24878 1327 24879 1353
rect 24851 1326 24879 1327
rect 24851 1193 24879 1194
rect 24851 1167 24852 1193
rect 24852 1167 24878 1193
rect 24878 1167 24879 1193
rect 24851 1166 24879 1167
rect 24851 1033 24879 1034
rect 24851 1007 24852 1033
rect 24852 1007 24878 1033
rect 24878 1007 24879 1033
rect 24851 1006 24879 1007
rect 24851 873 24879 874
rect 24851 847 24852 873
rect 24852 847 24878 873
rect 24878 847 24879 873
rect 24851 846 24879 847
rect 24851 713 24879 714
rect 24851 687 24852 713
rect 24852 687 24878 713
rect 24878 687 24879 713
rect 24851 686 24879 687
rect 24851 553 24879 554
rect 24851 527 24852 553
rect 24852 527 24878 553
rect 24878 527 24879 553
rect 24851 526 24879 527
rect 24851 393 24879 394
rect 24851 367 24852 393
rect 24852 367 24878 393
rect 24878 367 24879 393
rect 24851 366 24879 367
rect 24851 233 24879 234
rect 24851 207 24852 233
rect 24852 207 24878 233
rect 24878 207 24879 233
rect 24851 206 24879 207
rect 24851 73 24879 74
rect 24851 47 24852 73
rect 24852 47 24878 73
rect 24878 47 24879 73
rect 24851 46 24879 47
rect 24851 -87 24879 -86
rect 24851 -113 24852 -87
rect 24852 -113 24878 -87
rect 24878 -113 24879 -87
rect 24851 -114 24879 -113
rect 21118 -247 21146 -246
rect 21118 -273 21119 -247
rect 21119 -273 21145 -247
rect 21145 -273 21146 -247
rect 21118 -274 21146 -273
rect 24851 -247 24879 -246
rect 24851 -273 24852 -247
rect 24852 -273 24878 -247
rect 24878 -273 24879 -247
rect 24851 -274 24879 -273
rect 15306 -350 15334 -349
rect 15306 -376 15307 -350
rect 15307 -376 15333 -350
rect 15333 -376 15334 -350
rect 15306 -377 15334 -376
rect 15466 -350 15494 -349
rect 15466 -376 15467 -350
rect 15467 -376 15493 -350
rect 15493 -376 15494 -350
rect 15466 -377 15494 -376
rect 15626 -350 15654 -349
rect 15626 -376 15627 -350
rect 15627 -376 15653 -350
rect 15653 -376 15654 -350
rect 15626 -377 15654 -376
rect 15786 -350 15814 -349
rect 15786 -376 15787 -350
rect 15787 -376 15813 -350
rect 15813 -376 15814 -350
rect 15786 -377 15814 -376
rect 15946 -350 15974 -349
rect 15946 -376 15947 -350
rect 15947 -376 15973 -350
rect 15973 -376 15974 -350
rect 15946 -377 15974 -376
rect 16106 -350 16134 -349
rect 16106 -376 16107 -350
rect 16107 -376 16133 -350
rect 16133 -376 16134 -350
rect 16106 -377 16134 -376
rect 16266 -350 16294 -349
rect 16266 -376 16267 -350
rect 16267 -376 16293 -350
rect 16293 -376 16294 -350
rect 16266 -377 16294 -376
rect 16426 -350 16454 -349
rect 16426 -376 16427 -350
rect 16427 -376 16453 -350
rect 16453 -376 16454 -350
rect 16426 -377 16454 -376
rect 16586 -350 16614 -349
rect 16586 -376 16587 -350
rect 16587 -376 16613 -350
rect 16613 -376 16614 -350
rect 16586 -377 16614 -376
rect 16746 -350 16774 -349
rect 16746 -376 16747 -350
rect 16747 -376 16773 -350
rect 16773 -376 16774 -350
rect 16746 -377 16774 -376
rect 16906 -350 16934 -349
rect 16906 -376 16907 -350
rect 16907 -376 16933 -350
rect 16933 -376 16934 -350
rect 16906 -377 16934 -376
rect 17066 -350 17094 -349
rect 17066 -376 17067 -350
rect 17067 -376 17093 -350
rect 17093 -376 17094 -350
rect 17066 -377 17094 -376
rect 17226 -350 17254 -349
rect 17226 -376 17227 -350
rect 17227 -376 17253 -350
rect 17253 -376 17254 -350
rect 17226 -377 17254 -376
rect 17386 -350 17414 -349
rect 17386 -376 17387 -350
rect 17387 -376 17413 -350
rect 17413 -376 17414 -350
rect 17386 -377 17414 -376
rect 17546 -350 17574 -349
rect 17546 -376 17547 -350
rect 17547 -376 17573 -350
rect 17573 -376 17574 -350
rect 17546 -377 17574 -376
rect 17706 -350 17734 -349
rect 17706 -376 17707 -350
rect 17707 -376 17733 -350
rect 17733 -376 17734 -350
rect 17706 -377 17734 -376
rect 17866 -350 17894 -349
rect 17866 -376 17867 -350
rect 17867 -376 17893 -350
rect 17893 -376 17894 -350
rect 17866 -377 17894 -376
rect 18026 -350 18054 -349
rect 18026 -376 18027 -350
rect 18027 -376 18053 -350
rect 18053 -376 18054 -350
rect 18026 -377 18054 -376
rect 18186 -350 18214 -349
rect 18186 -376 18187 -350
rect 18187 -376 18213 -350
rect 18213 -376 18214 -350
rect 18186 -377 18214 -376
rect 18346 -350 18374 -349
rect 18346 -376 18347 -350
rect 18347 -376 18373 -350
rect 18373 -376 18374 -350
rect 18346 -377 18374 -376
rect 18506 -350 18534 -349
rect 18506 -376 18507 -350
rect 18507 -376 18533 -350
rect 18533 -376 18534 -350
rect 18506 -377 18534 -376
rect 18666 -350 18694 -349
rect 18666 -376 18667 -350
rect 18667 -376 18693 -350
rect 18693 -376 18694 -350
rect 18666 -377 18694 -376
rect 21306 -350 21334 -349
rect 21306 -376 21307 -350
rect 21307 -376 21333 -350
rect 21333 -376 21334 -350
rect 21306 -377 21334 -376
rect 21466 -350 21494 -349
rect 21466 -376 21467 -350
rect 21467 -376 21493 -350
rect 21493 -376 21494 -350
rect 21466 -377 21494 -376
rect 21626 -350 21654 -349
rect 21626 -376 21627 -350
rect 21627 -376 21653 -350
rect 21653 -376 21654 -350
rect 21626 -377 21654 -376
rect 21786 -350 21814 -349
rect 21786 -376 21787 -350
rect 21787 -376 21813 -350
rect 21813 -376 21814 -350
rect 21786 -377 21814 -376
rect 21946 -350 21974 -349
rect 21946 -376 21947 -350
rect 21947 -376 21973 -350
rect 21973 -376 21974 -350
rect 21946 -377 21974 -376
rect 22106 -350 22134 -349
rect 22106 -376 22107 -350
rect 22107 -376 22133 -350
rect 22133 -376 22134 -350
rect 22106 -377 22134 -376
rect 22266 -350 22294 -349
rect 22266 -376 22267 -350
rect 22267 -376 22293 -350
rect 22293 -376 22294 -350
rect 22266 -377 22294 -376
rect 22426 -350 22454 -349
rect 22426 -376 22427 -350
rect 22427 -376 22453 -350
rect 22453 -376 22454 -350
rect 22426 -377 22454 -376
rect 22586 -350 22614 -349
rect 22586 -376 22587 -350
rect 22587 -376 22613 -350
rect 22613 -376 22614 -350
rect 22586 -377 22614 -376
rect 22746 -350 22774 -349
rect 22746 -376 22747 -350
rect 22747 -376 22773 -350
rect 22773 -376 22774 -350
rect 22746 -377 22774 -376
rect 22906 -350 22934 -349
rect 22906 -376 22907 -350
rect 22907 -376 22933 -350
rect 22933 -376 22934 -350
rect 22906 -377 22934 -376
rect 23066 -350 23094 -349
rect 23066 -376 23067 -350
rect 23067 -376 23093 -350
rect 23093 -376 23094 -350
rect 23066 -377 23094 -376
rect 23226 -350 23254 -349
rect 23226 -376 23227 -350
rect 23227 -376 23253 -350
rect 23253 -376 23254 -350
rect 23226 -377 23254 -376
rect 23386 -350 23414 -349
rect 23386 -376 23387 -350
rect 23387 -376 23413 -350
rect 23413 -376 23414 -350
rect 23386 -377 23414 -376
rect 23546 -350 23574 -349
rect 23546 -376 23547 -350
rect 23547 -376 23573 -350
rect 23573 -376 23574 -350
rect 23546 -377 23574 -376
rect 23706 -350 23734 -349
rect 23706 -376 23707 -350
rect 23707 -376 23733 -350
rect 23733 -376 23734 -350
rect 23706 -377 23734 -376
rect 23866 -350 23894 -349
rect 23866 -376 23867 -350
rect 23867 -376 23893 -350
rect 23893 -376 23894 -350
rect 23866 -377 23894 -376
rect 24026 -350 24054 -349
rect 24026 -376 24027 -350
rect 24027 -376 24053 -350
rect 24053 -376 24054 -350
rect 24026 -377 24054 -376
rect 24186 -350 24214 -349
rect 24186 -376 24187 -350
rect 24187 -376 24213 -350
rect 24213 -376 24214 -350
rect 24186 -377 24214 -376
rect 24346 -350 24374 -349
rect 24346 -376 24347 -350
rect 24347 -376 24373 -350
rect 24373 -376 24374 -350
rect 24346 -377 24374 -376
rect 24506 -350 24534 -349
rect 24506 -376 24507 -350
rect 24507 -376 24533 -350
rect 24533 -376 24534 -350
rect 24506 -377 24534 -376
rect 24666 -350 24694 -349
rect 24666 -376 24667 -350
rect 24667 -376 24693 -350
rect 24693 -376 24694 -350
rect 24666 -377 24694 -376
rect 19440 -690 19480 -630
rect 20035 -1170 20065 -1140
rect 19965 -1245 19995 -1215
rect 20070 -1240 20100 -1210
rect 16155 -2100 16225 -2070
rect 16295 -2260 16365 -2230
rect 11635 -3770 11705 -3740
rect 11775 -3930 11845 -3900
rect 8200 -4790 8230 -4760
rect 8305 -4785 8335 -4755
rect 8235 -4860 8265 -4830
rect 8520 -5370 8560 -5310
rect 3306 -5624 3334 -5623
rect 3306 -5650 3307 -5624
rect 3307 -5650 3333 -5624
rect 3333 -5650 3334 -5624
rect 3306 -5651 3334 -5650
rect 3466 -5624 3494 -5623
rect 3466 -5650 3467 -5624
rect 3467 -5650 3493 -5624
rect 3493 -5650 3494 -5624
rect 3466 -5651 3494 -5650
rect 3626 -5624 3654 -5623
rect 3626 -5650 3627 -5624
rect 3627 -5650 3653 -5624
rect 3653 -5650 3654 -5624
rect 3626 -5651 3654 -5650
rect 3786 -5624 3814 -5623
rect 3786 -5650 3787 -5624
rect 3787 -5650 3813 -5624
rect 3813 -5650 3814 -5624
rect 3786 -5651 3814 -5650
rect 3946 -5624 3974 -5623
rect 3946 -5650 3947 -5624
rect 3947 -5650 3973 -5624
rect 3973 -5650 3974 -5624
rect 3946 -5651 3974 -5650
rect 4106 -5624 4134 -5623
rect 4106 -5650 4107 -5624
rect 4107 -5650 4133 -5624
rect 4133 -5650 4134 -5624
rect 4106 -5651 4134 -5650
rect 4266 -5624 4294 -5623
rect 4266 -5650 4267 -5624
rect 4267 -5650 4293 -5624
rect 4293 -5650 4294 -5624
rect 4266 -5651 4294 -5650
rect 4426 -5624 4454 -5623
rect 4426 -5650 4427 -5624
rect 4427 -5650 4453 -5624
rect 4453 -5650 4454 -5624
rect 4426 -5651 4454 -5650
rect 4586 -5624 4614 -5623
rect 4586 -5650 4587 -5624
rect 4587 -5650 4613 -5624
rect 4613 -5650 4614 -5624
rect 4586 -5651 4614 -5650
rect 4746 -5624 4774 -5623
rect 4746 -5650 4747 -5624
rect 4747 -5650 4773 -5624
rect 4773 -5650 4774 -5624
rect 4746 -5651 4774 -5650
rect 4906 -5624 4934 -5623
rect 4906 -5650 4907 -5624
rect 4907 -5650 4933 -5624
rect 4933 -5650 4934 -5624
rect 4906 -5651 4934 -5650
rect 5066 -5624 5094 -5623
rect 5066 -5650 5067 -5624
rect 5067 -5650 5093 -5624
rect 5093 -5650 5094 -5624
rect 5066 -5651 5094 -5650
rect 5226 -5624 5254 -5623
rect 5226 -5650 5227 -5624
rect 5227 -5650 5253 -5624
rect 5253 -5650 5254 -5624
rect 5226 -5651 5254 -5650
rect 5386 -5624 5414 -5623
rect 5386 -5650 5387 -5624
rect 5387 -5650 5413 -5624
rect 5413 -5650 5414 -5624
rect 5386 -5651 5414 -5650
rect 5546 -5624 5574 -5623
rect 5546 -5650 5547 -5624
rect 5547 -5650 5573 -5624
rect 5573 -5650 5574 -5624
rect 5546 -5651 5574 -5650
rect 5706 -5624 5734 -5623
rect 5706 -5650 5707 -5624
rect 5707 -5650 5733 -5624
rect 5733 -5650 5734 -5624
rect 5706 -5651 5734 -5650
rect 5866 -5624 5894 -5623
rect 5866 -5650 5867 -5624
rect 5867 -5650 5893 -5624
rect 5893 -5650 5894 -5624
rect 5866 -5651 5894 -5650
rect 6026 -5624 6054 -5623
rect 6026 -5650 6027 -5624
rect 6027 -5650 6053 -5624
rect 6053 -5650 6054 -5624
rect 6026 -5651 6054 -5650
rect 6186 -5624 6214 -5623
rect 6186 -5650 6187 -5624
rect 6187 -5650 6213 -5624
rect 6213 -5650 6214 -5624
rect 6186 -5651 6214 -5650
rect 6346 -5624 6374 -5623
rect 6346 -5650 6347 -5624
rect 6347 -5650 6373 -5624
rect 6373 -5650 6374 -5624
rect 6346 -5651 6374 -5650
rect 6506 -5624 6534 -5623
rect 6506 -5650 6507 -5624
rect 6507 -5650 6533 -5624
rect 6533 -5650 6534 -5624
rect 6506 -5651 6534 -5650
rect 6666 -5624 6694 -5623
rect 6666 -5650 6667 -5624
rect 6667 -5650 6693 -5624
rect 6693 -5650 6694 -5624
rect 6666 -5651 6694 -5650
rect 9306 -5624 9334 -5623
rect 9306 -5650 9307 -5624
rect 9307 -5650 9333 -5624
rect 9333 -5650 9334 -5624
rect 9306 -5651 9334 -5650
rect 9466 -5624 9494 -5623
rect 9466 -5650 9467 -5624
rect 9467 -5650 9493 -5624
rect 9493 -5650 9494 -5624
rect 9466 -5651 9494 -5650
rect 9626 -5624 9654 -5623
rect 9626 -5650 9627 -5624
rect 9627 -5650 9653 -5624
rect 9653 -5650 9654 -5624
rect 9626 -5651 9654 -5650
rect 9786 -5624 9814 -5623
rect 9786 -5650 9787 -5624
rect 9787 -5650 9813 -5624
rect 9813 -5650 9814 -5624
rect 9786 -5651 9814 -5650
rect 9946 -5624 9974 -5623
rect 9946 -5650 9947 -5624
rect 9947 -5650 9973 -5624
rect 9973 -5650 9974 -5624
rect 9946 -5651 9974 -5650
rect 10106 -5624 10134 -5623
rect 10106 -5650 10107 -5624
rect 10107 -5650 10133 -5624
rect 10133 -5650 10134 -5624
rect 10106 -5651 10134 -5650
rect 10266 -5624 10294 -5623
rect 10266 -5650 10267 -5624
rect 10267 -5650 10293 -5624
rect 10293 -5650 10294 -5624
rect 10266 -5651 10294 -5650
rect 10426 -5624 10454 -5623
rect 10426 -5650 10427 -5624
rect 10427 -5650 10453 -5624
rect 10453 -5650 10454 -5624
rect 10426 -5651 10454 -5650
rect 10586 -5624 10614 -5623
rect 10586 -5650 10587 -5624
rect 10587 -5650 10613 -5624
rect 10613 -5650 10614 -5624
rect 10586 -5651 10614 -5650
rect 10746 -5624 10774 -5623
rect 10746 -5650 10747 -5624
rect 10747 -5650 10773 -5624
rect 10773 -5650 10774 -5624
rect 10746 -5651 10774 -5650
rect 10906 -5624 10934 -5623
rect 10906 -5650 10907 -5624
rect 10907 -5650 10933 -5624
rect 10933 -5650 10934 -5624
rect 10906 -5651 10934 -5650
rect 11066 -5624 11094 -5623
rect 11066 -5650 11067 -5624
rect 11067 -5650 11093 -5624
rect 11093 -5650 11094 -5624
rect 11066 -5651 11094 -5650
rect 11226 -5624 11254 -5623
rect 11226 -5650 11227 -5624
rect 11227 -5650 11253 -5624
rect 11253 -5650 11254 -5624
rect 11226 -5651 11254 -5650
rect 11386 -5624 11414 -5623
rect 11386 -5650 11387 -5624
rect 11387 -5650 11413 -5624
rect 11413 -5650 11414 -5624
rect 11386 -5651 11414 -5650
rect 11546 -5624 11574 -5623
rect 11546 -5650 11547 -5624
rect 11547 -5650 11573 -5624
rect 11573 -5650 11574 -5624
rect 11546 -5651 11574 -5650
rect 11706 -5624 11734 -5623
rect 11706 -5650 11707 -5624
rect 11707 -5650 11733 -5624
rect 11733 -5650 11734 -5624
rect 11706 -5651 11734 -5650
rect 11866 -5624 11894 -5623
rect 11866 -5650 11867 -5624
rect 11867 -5650 11893 -5624
rect 11893 -5650 11894 -5624
rect 11866 -5651 11894 -5650
rect 12026 -5624 12054 -5623
rect 12026 -5650 12027 -5624
rect 12027 -5650 12053 -5624
rect 12053 -5650 12054 -5624
rect 12026 -5651 12054 -5650
rect 12186 -5624 12214 -5623
rect 12186 -5650 12187 -5624
rect 12187 -5650 12213 -5624
rect 12213 -5650 12214 -5624
rect 12186 -5651 12214 -5650
rect 12346 -5624 12374 -5623
rect 12346 -5650 12347 -5624
rect 12347 -5650 12373 -5624
rect 12373 -5650 12374 -5624
rect 12346 -5651 12374 -5650
rect 12506 -5624 12534 -5623
rect 12506 -5650 12507 -5624
rect 12507 -5650 12533 -5624
rect 12533 -5650 12534 -5624
rect 12506 -5651 12534 -5650
rect 12666 -5624 12694 -5623
rect 12666 -5650 12667 -5624
rect 12667 -5650 12693 -5624
rect 12693 -5650 12694 -5624
rect 12666 -5651 12694 -5650
rect 3121 -5727 3149 -5726
rect 3121 -5753 3122 -5727
rect 3122 -5753 3148 -5727
rect 3148 -5753 3149 -5727
rect 3121 -5754 3149 -5753
rect 6854 -5727 6882 -5726
rect 6854 -5753 6855 -5727
rect 6855 -5753 6881 -5727
rect 6881 -5753 6882 -5727
rect 6854 -5754 6882 -5753
rect 3121 -5887 3149 -5886
rect 3121 -5913 3122 -5887
rect 3122 -5913 3148 -5887
rect 3148 -5913 3149 -5887
rect 3121 -5914 3149 -5913
rect 3121 -6047 3149 -6046
rect 3121 -6073 3122 -6047
rect 3122 -6073 3148 -6047
rect 3148 -6073 3149 -6047
rect 3121 -6074 3149 -6073
rect 3121 -6207 3149 -6206
rect 3121 -6233 3122 -6207
rect 3122 -6233 3148 -6207
rect 3148 -6233 3149 -6207
rect 3121 -6234 3149 -6233
rect 3121 -6367 3149 -6366
rect 3121 -6393 3122 -6367
rect 3122 -6393 3148 -6367
rect 3148 -6393 3149 -6367
rect 3121 -6394 3149 -6393
rect 3121 -6527 3149 -6526
rect 3121 -6553 3122 -6527
rect 3122 -6553 3148 -6527
rect 3148 -6553 3149 -6527
rect 3121 -6554 3149 -6553
rect 3121 -6687 3149 -6686
rect 3121 -6713 3122 -6687
rect 3122 -6713 3148 -6687
rect 3148 -6713 3149 -6687
rect 3121 -6714 3149 -6713
rect 3121 -6847 3149 -6846
rect 3121 -6873 3122 -6847
rect 3122 -6873 3148 -6847
rect 3148 -6873 3149 -6847
rect 3121 -6874 3149 -6873
rect 3121 -7007 3149 -7006
rect 3121 -7033 3122 -7007
rect 3122 -7033 3148 -7007
rect 3148 -7033 3149 -7007
rect 3121 -7034 3149 -7033
rect 3121 -7167 3149 -7166
rect 3121 -7193 3122 -7167
rect 3122 -7193 3148 -7167
rect 3148 -7193 3149 -7167
rect 3121 -7194 3149 -7193
rect 3121 -7327 3149 -7326
rect 3121 -7353 3122 -7327
rect 3122 -7353 3148 -7327
rect 3148 -7353 3149 -7327
rect 3121 -7354 3149 -7353
rect 3121 -7487 3149 -7486
rect 3121 -7513 3122 -7487
rect 3122 -7513 3148 -7487
rect 3148 -7513 3149 -7487
rect 3121 -7514 3149 -7513
rect 3121 -7647 3149 -7646
rect 3121 -7673 3122 -7647
rect 3122 -7673 3148 -7647
rect 3148 -7673 3149 -7647
rect 3121 -7674 3149 -7673
rect 3121 -7807 3149 -7806
rect 3121 -7833 3122 -7807
rect 3122 -7833 3148 -7807
rect 3148 -7833 3149 -7807
rect 3121 -7834 3149 -7833
rect 3121 -7967 3149 -7966
rect 3121 -7993 3122 -7967
rect 3122 -7993 3148 -7967
rect 3148 -7993 3149 -7967
rect 3121 -7994 3149 -7993
rect 3121 -8127 3149 -8126
rect 3121 -8153 3122 -8127
rect 3122 -8153 3148 -8127
rect 3148 -8153 3149 -8127
rect 3121 -8154 3149 -8153
rect 3121 -8287 3149 -8286
rect 3121 -8313 3122 -8287
rect 3122 -8313 3148 -8287
rect 3148 -8313 3149 -8287
rect 3121 -8314 3149 -8313
rect 3121 -8447 3149 -8446
rect 3121 -8473 3122 -8447
rect 3122 -8473 3148 -8447
rect 3148 -8473 3149 -8447
rect 3121 -8474 3149 -8473
rect 3121 -8607 3149 -8606
rect 3121 -8633 3122 -8607
rect 3122 -8633 3148 -8607
rect 3148 -8633 3149 -8607
rect 3121 -8634 3149 -8633
rect 3121 -8767 3149 -8766
rect 3121 -8793 3122 -8767
rect 3122 -8793 3148 -8767
rect 3148 -8793 3149 -8767
rect 3121 -8794 3149 -8793
rect 3121 -8927 3149 -8926
rect 3121 -8953 3122 -8927
rect 3122 -8953 3148 -8927
rect 3148 -8953 3149 -8927
rect 3121 -8954 3149 -8953
rect 3121 -9087 3149 -9086
rect 3121 -9113 3122 -9087
rect 3122 -9113 3148 -9087
rect 3148 -9113 3149 -9087
rect 3121 -9114 3149 -9113
rect 6854 -5887 6882 -5886
rect 6854 -5913 6855 -5887
rect 6855 -5913 6881 -5887
rect 6881 -5913 6882 -5887
rect 6854 -5914 6882 -5913
rect 6854 -6047 6882 -6046
rect 6854 -6073 6855 -6047
rect 6855 -6073 6881 -6047
rect 6881 -6073 6882 -6047
rect 6854 -6074 6882 -6073
rect 6854 -6207 6882 -6206
rect 6854 -6233 6855 -6207
rect 6855 -6233 6881 -6207
rect 6881 -6233 6882 -6207
rect 6854 -6234 6882 -6233
rect 6854 -6367 6882 -6366
rect 6854 -6393 6855 -6367
rect 6855 -6393 6881 -6367
rect 6881 -6393 6882 -6367
rect 6854 -6394 6882 -6393
rect 6854 -6527 6882 -6526
rect 6854 -6553 6855 -6527
rect 6855 -6553 6881 -6527
rect 6881 -6553 6882 -6527
rect 6854 -6554 6882 -6553
rect 6854 -6687 6882 -6686
rect 6854 -6713 6855 -6687
rect 6855 -6713 6881 -6687
rect 6881 -6713 6882 -6687
rect 6854 -6714 6882 -6713
rect 6854 -6847 6882 -6846
rect 6854 -6873 6855 -6847
rect 6855 -6873 6881 -6847
rect 6881 -6873 6882 -6847
rect 6854 -6874 6882 -6873
rect 6854 -7007 6882 -7006
rect 6854 -7033 6855 -7007
rect 6855 -7033 6881 -7007
rect 6881 -7033 6882 -7007
rect 6854 -7034 6882 -7033
rect 6854 -7167 6882 -7166
rect 6854 -7193 6855 -7167
rect 6855 -7193 6881 -7167
rect 6881 -7193 6882 -7167
rect 6854 -7194 6882 -7193
rect 6854 -7327 6882 -7326
rect 6854 -7353 6855 -7327
rect 6855 -7353 6881 -7327
rect 6881 -7353 6882 -7327
rect 6854 -7354 6882 -7353
rect 6854 -7487 6882 -7486
rect 6854 -7513 6855 -7487
rect 6855 -7513 6881 -7487
rect 6881 -7513 6882 -7487
rect 6854 -7514 6882 -7513
rect 6854 -7647 6882 -7646
rect 6854 -7673 6855 -7647
rect 6855 -7673 6881 -7647
rect 6881 -7673 6882 -7647
rect 6854 -7674 6882 -7673
rect 6854 -7807 6882 -7806
rect 6854 -7833 6855 -7807
rect 6855 -7833 6881 -7807
rect 6881 -7833 6882 -7807
rect 6854 -7834 6882 -7833
rect 6854 -7967 6882 -7966
rect 6854 -7993 6855 -7967
rect 6855 -7993 6881 -7967
rect 6881 -7993 6882 -7967
rect 6854 -7994 6882 -7993
rect 6854 -8127 6882 -8126
rect 6854 -8153 6855 -8127
rect 6855 -8153 6881 -8127
rect 6881 -8153 6882 -8127
rect 6854 -8154 6882 -8153
rect 6854 -8287 6882 -8286
rect 6854 -8313 6855 -8287
rect 6855 -8313 6881 -8287
rect 6881 -8313 6882 -8287
rect 6854 -8314 6882 -8313
rect 6854 -8447 6882 -8446
rect 6854 -8473 6855 -8447
rect 6855 -8473 6881 -8447
rect 6881 -8473 6882 -8447
rect 6854 -8474 6882 -8473
rect 6854 -8607 6882 -8606
rect 6854 -8633 6855 -8607
rect 6855 -8633 6881 -8607
rect 6881 -8633 6882 -8607
rect 6854 -8634 6882 -8633
rect 6854 -8767 6882 -8766
rect 6854 -8793 6855 -8767
rect 6855 -8793 6881 -8767
rect 6881 -8793 6882 -8767
rect 6854 -8794 6882 -8793
rect 6854 -8927 6882 -8926
rect 6854 -8953 6855 -8927
rect 6855 -8953 6881 -8927
rect 6881 -8953 6882 -8927
rect 6854 -8954 6882 -8953
rect 6854 -9087 6882 -9086
rect 6854 -9113 6855 -9087
rect 6855 -9113 6881 -9087
rect 6881 -9113 6882 -9087
rect 6854 -9114 6882 -9113
rect 3121 -9247 3149 -9246
rect 3121 -9273 3122 -9247
rect 3122 -9273 3148 -9247
rect 3148 -9273 3149 -9247
rect 3121 -9274 3149 -9273
rect 6854 -9247 6882 -9246
rect 6854 -9273 6855 -9247
rect 6855 -9273 6881 -9247
rect 6881 -9273 6882 -9247
rect 6854 -9274 6882 -9273
rect 3306 -9352 3334 -9351
rect 3306 -9378 3307 -9352
rect 3307 -9378 3333 -9352
rect 3333 -9378 3334 -9352
rect 3306 -9379 3334 -9378
rect 3466 -9352 3494 -9351
rect 3466 -9378 3467 -9352
rect 3467 -9378 3493 -9352
rect 3493 -9378 3494 -9352
rect 3466 -9379 3494 -9378
rect 3626 -9352 3654 -9351
rect 3626 -9378 3627 -9352
rect 3627 -9378 3653 -9352
rect 3653 -9378 3654 -9352
rect 3626 -9379 3654 -9378
rect 3786 -9352 3814 -9351
rect 3786 -9378 3787 -9352
rect 3787 -9378 3813 -9352
rect 3813 -9378 3814 -9352
rect 3786 -9379 3814 -9378
rect 3946 -9352 3974 -9351
rect 3946 -9378 3947 -9352
rect 3947 -9378 3973 -9352
rect 3973 -9378 3974 -9352
rect 3946 -9379 3974 -9378
rect 4106 -9352 4134 -9351
rect 4106 -9378 4107 -9352
rect 4107 -9378 4133 -9352
rect 4133 -9378 4134 -9352
rect 4106 -9379 4134 -9378
rect 4266 -9352 4294 -9351
rect 4266 -9378 4267 -9352
rect 4267 -9378 4293 -9352
rect 4293 -9378 4294 -9352
rect 4266 -9379 4294 -9378
rect 4426 -9352 4454 -9351
rect 4426 -9378 4427 -9352
rect 4427 -9378 4453 -9352
rect 4453 -9378 4454 -9352
rect 4426 -9379 4454 -9378
rect 4586 -9352 4614 -9351
rect 4586 -9378 4587 -9352
rect 4587 -9378 4613 -9352
rect 4613 -9378 4614 -9352
rect 4586 -9379 4614 -9378
rect 4746 -9352 4774 -9351
rect 4746 -9378 4747 -9352
rect 4747 -9378 4773 -9352
rect 4773 -9378 4774 -9352
rect 4746 -9379 4774 -9378
rect 4906 -9352 4934 -9351
rect 4906 -9378 4907 -9352
rect 4907 -9378 4933 -9352
rect 4933 -9378 4934 -9352
rect 4906 -9379 4934 -9378
rect 5066 -9352 5094 -9351
rect 5066 -9378 5067 -9352
rect 5067 -9378 5093 -9352
rect 5093 -9378 5094 -9352
rect 5066 -9379 5094 -9378
rect 5226 -9352 5254 -9351
rect 5226 -9378 5227 -9352
rect 5227 -9378 5253 -9352
rect 5253 -9378 5254 -9352
rect 5226 -9379 5254 -9378
rect 5386 -9352 5414 -9351
rect 5386 -9378 5387 -9352
rect 5387 -9378 5413 -9352
rect 5413 -9378 5414 -9352
rect 5386 -9379 5414 -9378
rect 5546 -9352 5574 -9351
rect 5546 -9378 5547 -9352
rect 5547 -9378 5573 -9352
rect 5573 -9378 5574 -9352
rect 5546 -9379 5574 -9378
rect 5706 -9352 5734 -9351
rect 5706 -9378 5707 -9352
rect 5707 -9378 5733 -9352
rect 5733 -9378 5734 -9352
rect 5706 -9379 5734 -9378
rect 5866 -9352 5894 -9351
rect 5866 -9378 5867 -9352
rect 5867 -9378 5893 -9352
rect 5893 -9378 5894 -9352
rect 5866 -9379 5894 -9378
rect 6026 -9352 6054 -9351
rect 6026 -9378 6027 -9352
rect 6027 -9378 6053 -9352
rect 6053 -9378 6054 -9352
rect 6026 -9379 6054 -9378
rect 6186 -9352 6214 -9351
rect 6186 -9378 6187 -9352
rect 6187 -9378 6213 -9352
rect 6213 -9378 6214 -9352
rect 6186 -9379 6214 -9378
rect 6346 -9352 6374 -9351
rect 6346 -9378 6347 -9352
rect 6347 -9378 6373 -9352
rect 6373 -9378 6374 -9352
rect 6346 -9379 6374 -9378
rect 6506 -9352 6534 -9351
rect 6506 -9378 6507 -9352
rect 6507 -9378 6533 -9352
rect 6533 -9378 6534 -9352
rect 6506 -9379 6534 -9378
rect 6666 -9352 6694 -9351
rect 6666 -9378 6667 -9352
rect 6667 -9378 6693 -9352
rect 6693 -9378 6694 -9352
rect 6666 -9379 6694 -9378
rect 9121 -5727 9149 -5726
rect 9121 -5753 9122 -5727
rect 9122 -5753 9148 -5727
rect 9148 -5753 9149 -5727
rect 9121 -5754 9149 -5753
rect 12854 -5727 12882 -5726
rect 12854 -5753 12855 -5727
rect 12855 -5753 12881 -5727
rect 12881 -5753 12882 -5727
rect 12854 -5754 12882 -5753
rect 9121 -5887 9149 -5886
rect 9121 -5913 9122 -5887
rect 9122 -5913 9148 -5887
rect 9148 -5913 9149 -5887
rect 9121 -5914 9149 -5913
rect 9121 -6047 9149 -6046
rect 9121 -6073 9122 -6047
rect 9122 -6073 9148 -6047
rect 9148 -6073 9149 -6047
rect 9121 -6074 9149 -6073
rect 9121 -6207 9149 -6206
rect 9121 -6233 9122 -6207
rect 9122 -6233 9148 -6207
rect 9148 -6233 9149 -6207
rect 9121 -6234 9149 -6233
rect 9121 -6367 9149 -6366
rect 9121 -6393 9122 -6367
rect 9122 -6393 9148 -6367
rect 9148 -6393 9149 -6367
rect 9121 -6394 9149 -6393
rect 9121 -6527 9149 -6526
rect 9121 -6553 9122 -6527
rect 9122 -6553 9148 -6527
rect 9148 -6553 9149 -6527
rect 9121 -6554 9149 -6553
rect 9121 -6687 9149 -6686
rect 9121 -6713 9122 -6687
rect 9122 -6713 9148 -6687
rect 9148 -6713 9149 -6687
rect 9121 -6714 9149 -6713
rect 9121 -6847 9149 -6846
rect 9121 -6873 9122 -6847
rect 9122 -6873 9148 -6847
rect 9148 -6873 9149 -6847
rect 9121 -6874 9149 -6873
rect 9121 -7007 9149 -7006
rect 9121 -7033 9122 -7007
rect 9122 -7033 9148 -7007
rect 9148 -7033 9149 -7007
rect 9121 -7034 9149 -7033
rect 9121 -7167 9149 -7166
rect 9121 -7193 9122 -7167
rect 9122 -7193 9148 -7167
rect 9148 -7193 9149 -7167
rect 9121 -7194 9149 -7193
rect 9121 -7327 9149 -7326
rect 9121 -7353 9122 -7327
rect 9122 -7353 9148 -7327
rect 9148 -7353 9149 -7327
rect 9121 -7354 9149 -7353
rect 9121 -7487 9149 -7486
rect 9121 -7513 9122 -7487
rect 9122 -7513 9148 -7487
rect 9148 -7513 9149 -7487
rect 9121 -7514 9149 -7513
rect 9121 -7647 9149 -7646
rect 9121 -7673 9122 -7647
rect 9122 -7673 9148 -7647
rect 9148 -7673 9149 -7647
rect 9121 -7674 9149 -7673
rect 9121 -7807 9149 -7806
rect 9121 -7833 9122 -7807
rect 9122 -7833 9148 -7807
rect 9148 -7833 9149 -7807
rect 9121 -7834 9149 -7833
rect 9121 -7967 9149 -7966
rect 9121 -7993 9122 -7967
rect 9122 -7993 9148 -7967
rect 9148 -7993 9149 -7967
rect 9121 -7994 9149 -7993
rect 9121 -8127 9149 -8126
rect 9121 -8153 9122 -8127
rect 9122 -8153 9148 -8127
rect 9148 -8153 9149 -8127
rect 9121 -8154 9149 -8153
rect 9121 -8287 9149 -8286
rect 9121 -8313 9122 -8287
rect 9122 -8313 9148 -8287
rect 9148 -8313 9149 -8287
rect 9121 -8314 9149 -8313
rect 9121 -8447 9149 -8446
rect 9121 -8473 9122 -8447
rect 9122 -8473 9148 -8447
rect 9148 -8473 9149 -8447
rect 9121 -8474 9149 -8473
rect 9121 -8607 9149 -8606
rect 9121 -8633 9122 -8607
rect 9122 -8633 9148 -8607
rect 9148 -8633 9149 -8607
rect 9121 -8634 9149 -8633
rect 9121 -8767 9149 -8766
rect 9121 -8793 9122 -8767
rect 9122 -8793 9148 -8767
rect 9148 -8793 9149 -8767
rect 9121 -8794 9149 -8793
rect 9121 -8927 9149 -8926
rect 9121 -8953 9122 -8927
rect 9122 -8953 9148 -8927
rect 9148 -8953 9149 -8927
rect 9121 -8954 9149 -8953
rect 9121 -9087 9149 -9086
rect 9121 -9113 9122 -9087
rect 9122 -9113 9148 -9087
rect 9148 -9113 9149 -9087
rect 9121 -9114 9149 -9113
rect 12854 -5887 12882 -5886
rect 12854 -5913 12855 -5887
rect 12855 -5913 12881 -5887
rect 12881 -5913 12882 -5887
rect 12854 -5914 12882 -5913
rect 12854 -6047 12882 -6046
rect 12854 -6073 12855 -6047
rect 12855 -6073 12881 -6047
rect 12881 -6073 12882 -6047
rect 12854 -6074 12882 -6073
rect 12854 -6207 12882 -6206
rect 12854 -6233 12855 -6207
rect 12855 -6233 12881 -6207
rect 12881 -6233 12882 -6207
rect 12854 -6234 12882 -6233
rect 12854 -6367 12882 -6366
rect 12854 -6393 12855 -6367
rect 12855 -6393 12881 -6367
rect 12881 -6393 12882 -6367
rect 12854 -6394 12882 -6393
rect 12854 -6527 12882 -6526
rect 12854 -6553 12855 -6527
rect 12855 -6553 12881 -6527
rect 12881 -6553 12882 -6527
rect 12854 -6554 12882 -6553
rect 12854 -6687 12882 -6686
rect 12854 -6713 12855 -6687
rect 12855 -6713 12881 -6687
rect 12881 -6713 12882 -6687
rect 12854 -6714 12882 -6713
rect 12854 -6847 12882 -6846
rect 12854 -6873 12855 -6847
rect 12855 -6873 12881 -6847
rect 12881 -6873 12882 -6847
rect 12854 -6874 12882 -6873
rect 12854 -7007 12882 -7006
rect 12854 -7033 12855 -7007
rect 12855 -7033 12881 -7007
rect 12881 -7033 12882 -7007
rect 12854 -7034 12882 -7033
rect 12854 -7167 12882 -7166
rect 12854 -7193 12855 -7167
rect 12855 -7193 12881 -7167
rect 12881 -7193 12882 -7167
rect 12854 -7194 12882 -7193
rect 12854 -7327 12882 -7326
rect 12854 -7353 12855 -7327
rect 12855 -7353 12881 -7327
rect 12881 -7353 12882 -7327
rect 12854 -7354 12882 -7353
rect 12854 -7487 12882 -7486
rect 12854 -7513 12855 -7487
rect 12855 -7513 12881 -7487
rect 12881 -7513 12882 -7487
rect 12854 -7514 12882 -7513
rect 12854 -7647 12882 -7646
rect 12854 -7673 12855 -7647
rect 12855 -7673 12881 -7647
rect 12881 -7673 12882 -7647
rect 12854 -7674 12882 -7673
rect 12854 -7807 12882 -7806
rect 12854 -7833 12855 -7807
rect 12855 -7833 12881 -7807
rect 12881 -7833 12882 -7807
rect 12854 -7834 12882 -7833
rect 12854 -7967 12882 -7966
rect 12854 -7993 12855 -7967
rect 12855 -7993 12881 -7967
rect 12881 -7993 12882 -7967
rect 12854 -7994 12882 -7993
rect 12854 -8127 12882 -8126
rect 12854 -8153 12855 -8127
rect 12855 -8153 12881 -8127
rect 12881 -8153 12882 -8127
rect 12854 -8154 12882 -8153
rect 12854 -8287 12882 -8286
rect 12854 -8313 12855 -8287
rect 12855 -8313 12881 -8287
rect 12881 -8313 12882 -8287
rect 12854 -8314 12882 -8313
rect 12854 -8447 12882 -8446
rect 12854 -8473 12855 -8447
rect 12855 -8473 12881 -8447
rect 12881 -8473 12882 -8447
rect 12854 -8474 12882 -8473
rect 12854 -8607 12882 -8606
rect 12854 -8633 12855 -8607
rect 12855 -8633 12881 -8607
rect 12881 -8633 12882 -8607
rect 12854 -8634 12882 -8633
rect 12854 -8767 12882 -8766
rect 12854 -8793 12855 -8767
rect 12855 -8793 12881 -8767
rect 12881 -8793 12882 -8767
rect 12854 -8794 12882 -8793
rect 12854 -8927 12882 -8926
rect 12854 -8953 12855 -8927
rect 12855 -8953 12881 -8927
rect 12881 -8953 12882 -8927
rect 12854 -8954 12882 -8953
rect 12854 -9087 12882 -9086
rect 12854 -9113 12855 -9087
rect 12855 -9113 12881 -9087
rect 12881 -9113 12882 -9087
rect 12854 -9114 12882 -9113
rect 9121 -9247 9149 -9246
rect 9121 -9273 9122 -9247
rect 9122 -9273 9148 -9247
rect 9148 -9273 9149 -9247
rect 9121 -9274 9149 -9273
rect 12854 -9247 12882 -9246
rect 12854 -9273 12855 -9247
rect 12855 -9273 12881 -9247
rect 12881 -9273 12882 -9247
rect 12854 -9274 12882 -9273
rect 9306 -9352 9334 -9351
rect 9306 -9378 9307 -9352
rect 9307 -9378 9333 -9352
rect 9333 -9378 9334 -9352
rect 9306 -9379 9334 -9378
rect 9466 -9352 9494 -9351
rect 9466 -9378 9467 -9352
rect 9467 -9378 9493 -9352
rect 9493 -9378 9494 -9352
rect 9466 -9379 9494 -9378
rect 9626 -9352 9654 -9351
rect 9626 -9378 9627 -9352
rect 9627 -9378 9653 -9352
rect 9653 -9378 9654 -9352
rect 9626 -9379 9654 -9378
rect 9786 -9352 9814 -9351
rect 9786 -9378 9787 -9352
rect 9787 -9378 9813 -9352
rect 9813 -9378 9814 -9352
rect 9786 -9379 9814 -9378
rect 9946 -9352 9974 -9351
rect 9946 -9378 9947 -9352
rect 9947 -9378 9973 -9352
rect 9973 -9378 9974 -9352
rect 9946 -9379 9974 -9378
rect 10106 -9352 10134 -9351
rect 10106 -9378 10107 -9352
rect 10107 -9378 10133 -9352
rect 10133 -9378 10134 -9352
rect 10106 -9379 10134 -9378
rect 10266 -9352 10294 -9351
rect 10266 -9378 10267 -9352
rect 10267 -9378 10293 -9352
rect 10293 -9378 10294 -9352
rect 10266 -9379 10294 -9378
rect 10426 -9352 10454 -9351
rect 10426 -9378 10427 -9352
rect 10427 -9378 10453 -9352
rect 10453 -9378 10454 -9352
rect 10426 -9379 10454 -9378
rect 10586 -9352 10614 -9351
rect 10586 -9378 10587 -9352
rect 10587 -9378 10613 -9352
rect 10613 -9378 10614 -9352
rect 10586 -9379 10614 -9378
rect 10746 -9352 10774 -9351
rect 10746 -9378 10747 -9352
rect 10747 -9378 10773 -9352
rect 10773 -9378 10774 -9352
rect 10746 -9379 10774 -9378
rect 10906 -9352 10934 -9351
rect 10906 -9378 10907 -9352
rect 10907 -9378 10933 -9352
rect 10933 -9378 10934 -9352
rect 10906 -9379 10934 -9378
rect 11066 -9352 11094 -9351
rect 11066 -9378 11067 -9352
rect 11067 -9378 11093 -9352
rect 11093 -9378 11094 -9352
rect 11066 -9379 11094 -9378
rect 11226 -9352 11254 -9351
rect 11226 -9378 11227 -9352
rect 11227 -9378 11253 -9352
rect 11253 -9378 11254 -9352
rect 11226 -9379 11254 -9378
rect 11386 -9352 11414 -9351
rect 11386 -9378 11387 -9352
rect 11387 -9378 11413 -9352
rect 11413 -9378 11414 -9352
rect 11386 -9379 11414 -9378
rect 11546 -9352 11574 -9351
rect 11546 -9378 11547 -9352
rect 11547 -9378 11573 -9352
rect 11573 -9378 11574 -9352
rect 11546 -9379 11574 -9378
rect 11706 -9352 11734 -9351
rect 11706 -9378 11707 -9352
rect 11707 -9378 11733 -9352
rect 11733 -9378 11734 -9352
rect 11706 -9379 11734 -9378
rect 11866 -9352 11894 -9351
rect 11866 -9378 11867 -9352
rect 11867 -9378 11893 -9352
rect 11893 -9378 11894 -9352
rect 11866 -9379 11894 -9378
rect 12026 -9352 12054 -9351
rect 12026 -9378 12027 -9352
rect 12027 -9378 12053 -9352
rect 12053 -9378 12054 -9352
rect 12026 -9379 12054 -9378
rect 12186 -9352 12214 -9351
rect 12186 -9378 12187 -9352
rect 12187 -9378 12213 -9352
rect 12213 -9378 12214 -9352
rect 12186 -9379 12214 -9378
rect 12346 -9352 12374 -9351
rect 12346 -9378 12347 -9352
rect 12347 -9378 12373 -9352
rect 12373 -9378 12374 -9352
rect 12346 -9379 12374 -9378
rect 12506 -9352 12534 -9351
rect 12506 -9378 12507 -9352
rect 12507 -9378 12533 -9352
rect 12533 -9378 12534 -9352
rect 12506 -9379 12534 -9378
rect 12666 -9352 12694 -9351
rect 12666 -9378 12667 -9352
rect 12667 -9378 12693 -9352
rect 12693 -9378 12694 -9352
rect 12666 -9379 12694 -9378
rect 15306 -5624 15334 -5623
rect 15306 -5650 15307 -5624
rect 15307 -5650 15333 -5624
rect 15333 -5650 15334 -5624
rect 15306 -5651 15334 -5650
rect 15466 -5624 15494 -5623
rect 15466 -5650 15467 -5624
rect 15467 -5650 15493 -5624
rect 15493 -5650 15494 -5624
rect 15466 -5651 15494 -5650
rect 15626 -5624 15654 -5623
rect 15626 -5650 15627 -5624
rect 15627 -5650 15653 -5624
rect 15653 -5650 15654 -5624
rect 15626 -5651 15654 -5650
rect 15786 -5624 15814 -5623
rect 15786 -5650 15787 -5624
rect 15787 -5650 15813 -5624
rect 15813 -5650 15814 -5624
rect 15786 -5651 15814 -5650
rect 15946 -5624 15974 -5623
rect 15946 -5650 15947 -5624
rect 15947 -5650 15973 -5624
rect 15973 -5650 15974 -5624
rect 15946 -5651 15974 -5650
rect 16106 -5624 16134 -5623
rect 16106 -5650 16107 -5624
rect 16107 -5650 16133 -5624
rect 16133 -5650 16134 -5624
rect 16106 -5651 16134 -5650
rect 16266 -5624 16294 -5623
rect 16266 -5650 16267 -5624
rect 16267 -5650 16293 -5624
rect 16293 -5650 16294 -5624
rect 16266 -5651 16294 -5650
rect 16426 -5624 16454 -5623
rect 16426 -5650 16427 -5624
rect 16427 -5650 16453 -5624
rect 16453 -5650 16454 -5624
rect 16426 -5651 16454 -5650
rect 16586 -5624 16614 -5623
rect 16586 -5650 16587 -5624
rect 16587 -5650 16613 -5624
rect 16613 -5650 16614 -5624
rect 16586 -5651 16614 -5650
rect 16746 -5624 16774 -5623
rect 16746 -5650 16747 -5624
rect 16747 -5650 16773 -5624
rect 16773 -5650 16774 -5624
rect 16746 -5651 16774 -5650
rect 16906 -5624 16934 -5623
rect 16906 -5650 16907 -5624
rect 16907 -5650 16933 -5624
rect 16933 -5650 16934 -5624
rect 16906 -5651 16934 -5650
rect 17066 -5624 17094 -5623
rect 17066 -5650 17067 -5624
rect 17067 -5650 17093 -5624
rect 17093 -5650 17094 -5624
rect 17066 -5651 17094 -5650
rect 17226 -5624 17254 -5623
rect 17226 -5650 17227 -5624
rect 17227 -5650 17253 -5624
rect 17253 -5650 17254 -5624
rect 17226 -5651 17254 -5650
rect 17386 -5624 17414 -5623
rect 17386 -5650 17387 -5624
rect 17387 -5650 17413 -5624
rect 17413 -5650 17414 -5624
rect 17386 -5651 17414 -5650
rect 17546 -5624 17574 -5623
rect 17546 -5650 17547 -5624
rect 17547 -5650 17573 -5624
rect 17573 -5650 17574 -5624
rect 17546 -5651 17574 -5650
rect 17706 -5624 17734 -5623
rect 17706 -5650 17707 -5624
rect 17707 -5650 17733 -5624
rect 17733 -5650 17734 -5624
rect 17706 -5651 17734 -5650
rect 17866 -5624 17894 -5623
rect 17866 -5650 17867 -5624
rect 17867 -5650 17893 -5624
rect 17893 -5650 17894 -5624
rect 17866 -5651 17894 -5650
rect 18026 -5624 18054 -5623
rect 18026 -5650 18027 -5624
rect 18027 -5650 18053 -5624
rect 18053 -5650 18054 -5624
rect 18026 -5651 18054 -5650
rect 18186 -5624 18214 -5623
rect 18186 -5650 18187 -5624
rect 18187 -5650 18213 -5624
rect 18213 -5650 18214 -5624
rect 18186 -5651 18214 -5650
rect 18346 -5624 18374 -5623
rect 18346 -5650 18347 -5624
rect 18347 -5650 18373 -5624
rect 18373 -5650 18374 -5624
rect 18346 -5651 18374 -5650
rect 18506 -5624 18534 -5623
rect 18506 -5650 18507 -5624
rect 18507 -5650 18533 -5624
rect 18533 -5650 18534 -5624
rect 18506 -5651 18534 -5650
rect 18666 -5624 18694 -5623
rect 18666 -5650 18667 -5624
rect 18667 -5650 18693 -5624
rect 18693 -5650 18694 -5624
rect 18666 -5651 18694 -5650
rect 15121 -5727 15149 -5726
rect 15121 -5753 15122 -5727
rect 15122 -5753 15148 -5727
rect 15148 -5753 15149 -5727
rect 15121 -5754 15149 -5753
rect 18854 -5727 18882 -5726
rect 18854 -5753 18855 -5727
rect 18855 -5753 18881 -5727
rect 18881 -5753 18882 -5727
rect 18854 -5754 18882 -5753
rect 15121 -5887 15149 -5886
rect 15121 -5913 15122 -5887
rect 15122 -5913 15148 -5887
rect 15148 -5913 15149 -5887
rect 15121 -5914 15149 -5913
rect 15121 -6047 15149 -6046
rect 15121 -6073 15122 -6047
rect 15122 -6073 15148 -6047
rect 15148 -6073 15149 -6047
rect 15121 -6074 15149 -6073
rect 15121 -6207 15149 -6206
rect 15121 -6233 15122 -6207
rect 15122 -6233 15148 -6207
rect 15148 -6233 15149 -6207
rect 15121 -6234 15149 -6233
rect 15121 -6367 15149 -6366
rect 15121 -6393 15122 -6367
rect 15122 -6393 15148 -6367
rect 15148 -6393 15149 -6367
rect 15121 -6394 15149 -6393
rect 15121 -6527 15149 -6526
rect 15121 -6553 15122 -6527
rect 15122 -6553 15148 -6527
rect 15148 -6553 15149 -6527
rect 15121 -6554 15149 -6553
rect 15121 -6687 15149 -6686
rect 15121 -6713 15122 -6687
rect 15122 -6713 15148 -6687
rect 15148 -6713 15149 -6687
rect 15121 -6714 15149 -6713
rect 15121 -6847 15149 -6846
rect 15121 -6873 15122 -6847
rect 15122 -6873 15148 -6847
rect 15148 -6873 15149 -6847
rect 15121 -6874 15149 -6873
rect 15121 -7007 15149 -7006
rect 15121 -7033 15122 -7007
rect 15122 -7033 15148 -7007
rect 15148 -7033 15149 -7007
rect 15121 -7034 15149 -7033
rect 15121 -7167 15149 -7166
rect 15121 -7193 15122 -7167
rect 15122 -7193 15148 -7167
rect 15148 -7193 15149 -7167
rect 15121 -7194 15149 -7193
rect 15121 -7327 15149 -7326
rect 15121 -7353 15122 -7327
rect 15122 -7353 15148 -7327
rect 15148 -7353 15149 -7327
rect 15121 -7354 15149 -7353
rect 15121 -7487 15149 -7486
rect 15121 -7513 15122 -7487
rect 15122 -7513 15148 -7487
rect 15148 -7513 15149 -7487
rect 15121 -7514 15149 -7513
rect 15121 -7647 15149 -7646
rect 15121 -7673 15122 -7647
rect 15122 -7673 15148 -7647
rect 15148 -7673 15149 -7647
rect 15121 -7674 15149 -7673
rect 15121 -7807 15149 -7806
rect 15121 -7833 15122 -7807
rect 15122 -7833 15148 -7807
rect 15148 -7833 15149 -7807
rect 15121 -7834 15149 -7833
rect 15121 -7967 15149 -7966
rect 15121 -7993 15122 -7967
rect 15122 -7993 15148 -7967
rect 15148 -7993 15149 -7967
rect 15121 -7994 15149 -7993
rect 15121 -8127 15149 -8126
rect 15121 -8153 15122 -8127
rect 15122 -8153 15148 -8127
rect 15148 -8153 15149 -8127
rect 15121 -8154 15149 -8153
rect 15121 -8287 15149 -8286
rect 15121 -8313 15122 -8287
rect 15122 -8313 15148 -8287
rect 15148 -8313 15149 -8287
rect 15121 -8314 15149 -8313
rect 15121 -8447 15149 -8446
rect 15121 -8473 15122 -8447
rect 15122 -8473 15148 -8447
rect 15148 -8473 15149 -8447
rect 15121 -8474 15149 -8473
rect 15121 -8607 15149 -8606
rect 15121 -8633 15122 -8607
rect 15122 -8633 15148 -8607
rect 15148 -8633 15149 -8607
rect 15121 -8634 15149 -8633
rect 15121 -8767 15149 -8766
rect 15121 -8793 15122 -8767
rect 15122 -8793 15148 -8767
rect 15148 -8793 15149 -8767
rect 15121 -8794 15149 -8793
rect 15121 -8927 15149 -8926
rect 15121 -8953 15122 -8927
rect 15122 -8953 15148 -8927
rect 15148 -8953 15149 -8927
rect 15121 -8954 15149 -8953
rect 15121 -9087 15149 -9086
rect 15121 -9113 15122 -9087
rect 15122 -9113 15148 -9087
rect 15148 -9113 15149 -9087
rect 15121 -9114 15149 -9113
rect 18854 -5887 18882 -5886
rect 18854 -5913 18855 -5887
rect 18855 -5913 18881 -5887
rect 18881 -5913 18882 -5887
rect 18854 -5914 18882 -5913
rect 18854 -6047 18882 -6046
rect 18854 -6073 18855 -6047
rect 18855 -6073 18881 -6047
rect 18881 -6073 18882 -6047
rect 18854 -6074 18882 -6073
rect 18854 -6207 18882 -6206
rect 18854 -6233 18855 -6207
rect 18855 -6233 18881 -6207
rect 18881 -6233 18882 -6207
rect 18854 -6234 18882 -6233
rect 18854 -6367 18882 -6366
rect 18854 -6393 18855 -6367
rect 18855 -6393 18881 -6367
rect 18881 -6393 18882 -6367
rect 18854 -6394 18882 -6393
rect 18854 -6527 18882 -6526
rect 18854 -6553 18855 -6527
rect 18855 -6553 18881 -6527
rect 18881 -6553 18882 -6527
rect 18854 -6554 18882 -6553
rect 18854 -6687 18882 -6686
rect 18854 -6713 18855 -6687
rect 18855 -6713 18881 -6687
rect 18881 -6713 18882 -6687
rect 18854 -6714 18882 -6713
rect 18854 -6847 18882 -6846
rect 18854 -6873 18855 -6847
rect 18855 -6873 18881 -6847
rect 18881 -6873 18882 -6847
rect 18854 -6874 18882 -6873
rect 18854 -7007 18882 -7006
rect 18854 -7033 18855 -7007
rect 18855 -7033 18881 -7007
rect 18881 -7033 18882 -7007
rect 18854 -7034 18882 -7033
rect 18854 -7167 18882 -7166
rect 18854 -7193 18855 -7167
rect 18855 -7193 18881 -7167
rect 18881 -7193 18882 -7167
rect 18854 -7194 18882 -7193
rect 18854 -7327 18882 -7326
rect 18854 -7353 18855 -7327
rect 18855 -7353 18881 -7327
rect 18881 -7353 18882 -7327
rect 18854 -7354 18882 -7353
rect 18854 -7487 18882 -7486
rect 18854 -7513 18855 -7487
rect 18855 -7513 18881 -7487
rect 18881 -7513 18882 -7487
rect 18854 -7514 18882 -7513
rect 18854 -7647 18882 -7646
rect 18854 -7673 18855 -7647
rect 18855 -7673 18881 -7647
rect 18881 -7673 18882 -7647
rect 18854 -7674 18882 -7673
rect 18854 -7807 18882 -7806
rect 18854 -7833 18855 -7807
rect 18855 -7833 18881 -7807
rect 18881 -7833 18882 -7807
rect 18854 -7834 18882 -7833
rect 18854 -7967 18882 -7966
rect 18854 -7993 18855 -7967
rect 18855 -7993 18881 -7967
rect 18881 -7993 18882 -7967
rect 18854 -7994 18882 -7993
rect 18854 -8127 18882 -8126
rect 18854 -8153 18855 -8127
rect 18855 -8153 18881 -8127
rect 18881 -8153 18882 -8127
rect 18854 -8154 18882 -8153
rect 18854 -8287 18882 -8286
rect 18854 -8313 18855 -8287
rect 18855 -8313 18881 -8287
rect 18881 -8313 18882 -8287
rect 18854 -8314 18882 -8313
rect 18854 -8447 18882 -8446
rect 18854 -8473 18855 -8447
rect 18855 -8473 18881 -8447
rect 18881 -8473 18882 -8447
rect 18854 -8474 18882 -8473
rect 18854 -8607 18882 -8606
rect 18854 -8633 18855 -8607
rect 18855 -8633 18881 -8607
rect 18881 -8633 18882 -8607
rect 18854 -8634 18882 -8633
rect 18854 -8767 18882 -8766
rect 18854 -8793 18855 -8767
rect 18855 -8793 18881 -8767
rect 18881 -8793 18882 -8767
rect 18854 -8794 18882 -8793
rect 18854 -8927 18882 -8926
rect 18854 -8953 18855 -8927
rect 18855 -8953 18881 -8927
rect 18881 -8953 18882 -8927
rect 18854 -8954 18882 -8953
rect 18854 -9087 18882 -9086
rect 18854 -9113 18855 -9087
rect 18855 -9113 18881 -9087
rect 18881 -9113 18882 -9087
rect 18854 -9114 18882 -9113
rect 15121 -9247 15149 -9246
rect 15121 -9273 15122 -9247
rect 15122 -9273 15148 -9247
rect 15148 -9273 15149 -9247
rect 15121 -9274 15149 -9273
rect 18854 -9247 18882 -9246
rect 18854 -9273 18855 -9247
rect 18855 -9273 18881 -9247
rect 18881 -9273 18882 -9247
rect 18854 -9274 18882 -9273
rect 15306 -9352 15334 -9351
rect 15306 -9378 15307 -9352
rect 15307 -9378 15333 -9352
rect 15333 -9378 15334 -9352
rect 15306 -9379 15334 -9378
rect 15466 -9352 15494 -9351
rect 15466 -9378 15467 -9352
rect 15467 -9378 15493 -9352
rect 15493 -9378 15494 -9352
rect 15466 -9379 15494 -9378
rect 15626 -9352 15654 -9351
rect 15626 -9378 15627 -9352
rect 15627 -9378 15653 -9352
rect 15653 -9378 15654 -9352
rect 15626 -9379 15654 -9378
rect 15786 -9352 15814 -9351
rect 15786 -9378 15787 -9352
rect 15787 -9378 15813 -9352
rect 15813 -9378 15814 -9352
rect 15786 -9379 15814 -9378
rect 15946 -9352 15974 -9351
rect 15946 -9378 15947 -9352
rect 15947 -9378 15973 -9352
rect 15973 -9378 15974 -9352
rect 15946 -9379 15974 -9378
rect 16106 -9352 16134 -9351
rect 16106 -9378 16107 -9352
rect 16107 -9378 16133 -9352
rect 16133 -9378 16134 -9352
rect 16106 -9379 16134 -9378
rect 16266 -9352 16294 -9351
rect 16266 -9378 16267 -9352
rect 16267 -9378 16293 -9352
rect 16293 -9378 16294 -9352
rect 16266 -9379 16294 -9378
rect 16426 -9352 16454 -9351
rect 16426 -9378 16427 -9352
rect 16427 -9378 16453 -9352
rect 16453 -9378 16454 -9352
rect 16426 -9379 16454 -9378
rect 16586 -9352 16614 -9351
rect 16586 -9378 16587 -9352
rect 16587 -9378 16613 -9352
rect 16613 -9378 16614 -9352
rect 16586 -9379 16614 -9378
rect 16746 -9352 16774 -9351
rect 16746 -9378 16747 -9352
rect 16747 -9378 16773 -9352
rect 16773 -9378 16774 -9352
rect 16746 -9379 16774 -9378
rect 16906 -9352 16934 -9351
rect 16906 -9378 16907 -9352
rect 16907 -9378 16933 -9352
rect 16933 -9378 16934 -9352
rect 16906 -9379 16934 -9378
rect 17066 -9352 17094 -9351
rect 17066 -9378 17067 -9352
rect 17067 -9378 17093 -9352
rect 17093 -9378 17094 -9352
rect 17066 -9379 17094 -9378
rect 17226 -9352 17254 -9351
rect 17226 -9378 17227 -9352
rect 17227 -9378 17253 -9352
rect 17253 -9378 17254 -9352
rect 17226 -9379 17254 -9378
rect 17386 -9352 17414 -9351
rect 17386 -9378 17387 -9352
rect 17387 -9378 17413 -9352
rect 17413 -9378 17414 -9352
rect 17386 -9379 17414 -9378
rect 17546 -9352 17574 -9351
rect 17546 -9378 17547 -9352
rect 17547 -9378 17573 -9352
rect 17573 -9378 17574 -9352
rect 17546 -9379 17574 -9378
rect 17706 -9352 17734 -9351
rect 17706 -9378 17707 -9352
rect 17707 -9378 17733 -9352
rect 17733 -9378 17734 -9352
rect 17706 -9379 17734 -9378
rect 17866 -9352 17894 -9351
rect 17866 -9378 17867 -9352
rect 17867 -9378 17893 -9352
rect 17893 -9378 17894 -9352
rect 17866 -9379 17894 -9378
rect 18026 -9352 18054 -9351
rect 18026 -9378 18027 -9352
rect 18027 -9378 18053 -9352
rect 18053 -9378 18054 -9352
rect 18026 -9379 18054 -9378
rect 18186 -9352 18214 -9351
rect 18186 -9378 18187 -9352
rect 18187 -9378 18213 -9352
rect 18213 -9378 18214 -9352
rect 18186 -9379 18214 -9378
rect 18346 -9352 18374 -9351
rect 18346 -9378 18347 -9352
rect 18347 -9378 18373 -9352
rect 18373 -9378 18374 -9352
rect 18346 -9379 18374 -9378
rect 18506 -9352 18534 -9351
rect 18506 -9378 18507 -9352
rect 18507 -9378 18533 -9352
rect 18533 -9378 18534 -9352
rect 18506 -9379 18534 -9378
rect 18666 -9352 18694 -9351
rect 18666 -9378 18667 -9352
rect 18667 -9378 18693 -9352
rect 18693 -9378 18694 -9352
rect 18666 -9379 18694 -9378
rect 21306 -5624 21334 -5623
rect 21306 -5650 21307 -5624
rect 21307 -5650 21333 -5624
rect 21333 -5650 21334 -5624
rect 21306 -5651 21334 -5650
rect 21466 -5624 21494 -5623
rect 21466 -5650 21467 -5624
rect 21467 -5650 21493 -5624
rect 21493 -5650 21494 -5624
rect 21466 -5651 21494 -5650
rect 21626 -5624 21654 -5623
rect 21626 -5650 21627 -5624
rect 21627 -5650 21653 -5624
rect 21653 -5650 21654 -5624
rect 21626 -5651 21654 -5650
rect 21786 -5624 21814 -5623
rect 21786 -5650 21787 -5624
rect 21787 -5650 21813 -5624
rect 21813 -5650 21814 -5624
rect 21786 -5651 21814 -5650
rect 21946 -5624 21974 -5623
rect 21946 -5650 21947 -5624
rect 21947 -5650 21973 -5624
rect 21973 -5650 21974 -5624
rect 21946 -5651 21974 -5650
rect 22106 -5624 22134 -5623
rect 22106 -5650 22107 -5624
rect 22107 -5650 22133 -5624
rect 22133 -5650 22134 -5624
rect 22106 -5651 22134 -5650
rect 22266 -5624 22294 -5623
rect 22266 -5650 22267 -5624
rect 22267 -5650 22293 -5624
rect 22293 -5650 22294 -5624
rect 22266 -5651 22294 -5650
rect 22426 -5624 22454 -5623
rect 22426 -5650 22427 -5624
rect 22427 -5650 22453 -5624
rect 22453 -5650 22454 -5624
rect 22426 -5651 22454 -5650
rect 22586 -5624 22614 -5623
rect 22586 -5650 22587 -5624
rect 22587 -5650 22613 -5624
rect 22613 -5650 22614 -5624
rect 22586 -5651 22614 -5650
rect 22746 -5624 22774 -5623
rect 22746 -5650 22747 -5624
rect 22747 -5650 22773 -5624
rect 22773 -5650 22774 -5624
rect 22746 -5651 22774 -5650
rect 22906 -5624 22934 -5623
rect 22906 -5650 22907 -5624
rect 22907 -5650 22933 -5624
rect 22933 -5650 22934 -5624
rect 22906 -5651 22934 -5650
rect 23066 -5624 23094 -5623
rect 23066 -5650 23067 -5624
rect 23067 -5650 23093 -5624
rect 23093 -5650 23094 -5624
rect 23066 -5651 23094 -5650
rect 23226 -5624 23254 -5623
rect 23226 -5650 23227 -5624
rect 23227 -5650 23253 -5624
rect 23253 -5650 23254 -5624
rect 23226 -5651 23254 -5650
rect 23386 -5624 23414 -5623
rect 23386 -5650 23387 -5624
rect 23387 -5650 23413 -5624
rect 23413 -5650 23414 -5624
rect 23386 -5651 23414 -5650
rect 23546 -5624 23574 -5623
rect 23546 -5650 23547 -5624
rect 23547 -5650 23573 -5624
rect 23573 -5650 23574 -5624
rect 23546 -5651 23574 -5650
rect 23706 -5624 23734 -5623
rect 23706 -5650 23707 -5624
rect 23707 -5650 23733 -5624
rect 23733 -5650 23734 -5624
rect 23706 -5651 23734 -5650
rect 23866 -5624 23894 -5623
rect 23866 -5650 23867 -5624
rect 23867 -5650 23893 -5624
rect 23893 -5650 23894 -5624
rect 23866 -5651 23894 -5650
rect 24026 -5624 24054 -5623
rect 24026 -5650 24027 -5624
rect 24027 -5650 24053 -5624
rect 24053 -5650 24054 -5624
rect 24026 -5651 24054 -5650
rect 24186 -5624 24214 -5623
rect 24186 -5650 24187 -5624
rect 24187 -5650 24213 -5624
rect 24213 -5650 24214 -5624
rect 24186 -5651 24214 -5650
rect 24346 -5624 24374 -5623
rect 24346 -5650 24347 -5624
rect 24347 -5650 24373 -5624
rect 24373 -5650 24374 -5624
rect 24346 -5651 24374 -5650
rect 24506 -5624 24534 -5623
rect 24506 -5650 24507 -5624
rect 24507 -5650 24533 -5624
rect 24533 -5650 24534 -5624
rect 24506 -5651 24534 -5650
rect 24666 -5624 24694 -5623
rect 24666 -5650 24667 -5624
rect 24667 -5650 24693 -5624
rect 24693 -5650 24694 -5624
rect 24666 -5651 24694 -5650
rect 21121 -5727 21149 -5726
rect 21121 -5753 21122 -5727
rect 21122 -5753 21148 -5727
rect 21148 -5753 21149 -5727
rect 21121 -5754 21149 -5753
rect 24854 -5727 24882 -5726
rect 24854 -5753 24855 -5727
rect 24855 -5753 24881 -5727
rect 24881 -5753 24882 -5727
rect 24854 -5754 24882 -5753
rect 21121 -5887 21149 -5886
rect 21121 -5913 21122 -5887
rect 21122 -5913 21148 -5887
rect 21148 -5913 21149 -5887
rect 21121 -5914 21149 -5913
rect 21121 -6047 21149 -6046
rect 21121 -6073 21122 -6047
rect 21122 -6073 21148 -6047
rect 21148 -6073 21149 -6047
rect 21121 -6074 21149 -6073
rect 21121 -6207 21149 -6206
rect 21121 -6233 21122 -6207
rect 21122 -6233 21148 -6207
rect 21148 -6233 21149 -6207
rect 21121 -6234 21149 -6233
rect 21121 -6367 21149 -6366
rect 21121 -6393 21122 -6367
rect 21122 -6393 21148 -6367
rect 21148 -6393 21149 -6367
rect 21121 -6394 21149 -6393
rect 21121 -6527 21149 -6526
rect 21121 -6553 21122 -6527
rect 21122 -6553 21148 -6527
rect 21148 -6553 21149 -6527
rect 21121 -6554 21149 -6553
rect 21121 -6687 21149 -6686
rect 21121 -6713 21122 -6687
rect 21122 -6713 21148 -6687
rect 21148 -6713 21149 -6687
rect 21121 -6714 21149 -6713
rect 21121 -6847 21149 -6846
rect 21121 -6873 21122 -6847
rect 21122 -6873 21148 -6847
rect 21148 -6873 21149 -6847
rect 21121 -6874 21149 -6873
rect 21121 -7007 21149 -7006
rect 21121 -7033 21122 -7007
rect 21122 -7033 21148 -7007
rect 21148 -7033 21149 -7007
rect 21121 -7034 21149 -7033
rect 21121 -7167 21149 -7166
rect 21121 -7193 21122 -7167
rect 21122 -7193 21148 -7167
rect 21148 -7193 21149 -7167
rect 21121 -7194 21149 -7193
rect 21121 -7327 21149 -7326
rect 21121 -7353 21122 -7327
rect 21122 -7353 21148 -7327
rect 21148 -7353 21149 -7327
rect 21121 -7354 21149 -7353
rect 21121 -7487 21149 -7486
rect 21121 -7513 21122 -7487
rect 21122 -7513 21148 -7487
rect 21148 -7513 21149 -7487
rect 21121 -7514 21149 -7513
rect 21121 -7647 21149 -7646
rect 21121 -7673 21122 -7647
rect 21122 -7673 21148 -7647
rect 21148 -7673 21149 -7647
rect 21121 -7674 21149 -7673
rect 21121 -7807 21149 -7806
rect 21121 -7833 21122 -7807
rect 21122 -7833 21148 -7807
rect 21148 -7833 21149 -7807
rect 21121 -7834 21149 -7833
rect 21121 -7967 21149 -7966
rect 21121 -7993 21122 -7967
rect 21122 -7993 21148 -7967
rect 21148 -7993 21149 -7967
rect 21121 -7994 21149 -7993
rect 21121 -8127 21149 -8126
rect 21121 -8153 21122 -8127
rect 21122 -8153 21148 -8127
rect 21148 -8153 21149 -8127
rect 21121 -8154 21149 -8153
rect 21121 -8287 21149 -8286
rect 21121 -8313 21122 -8287
rect 21122 -8313 21148 -8287
rect 21148 -8313 21149 -8287
rect 21121 -8314 21149 -8313
rect 21121 -8447 21149 -8446
rect 21121 -8473 21122 -8447
rect 21122 -8473 21148 -8447
rect 21148 -8473 21149 -8447
rect 21121 -8474 21149 -8473
rect 21121 -8607 21149 -8606
rect 21121 -8633 21122 -8607
rect 21122 -8633 21148 -8607
rect 21148 -8633 21149 -8607
rect 21121 -8634 21149 -8633
rect 21121 -8767 21149 -8766
rect 21121 -8793 21122 -8767
rect 21122 -8793 21148 -8767
rect 21148 -8793 21149 -8767
rect 21121 -8794 21149 -8793
rect 21121 -8927 21149 -8926
rect 21121 -8953 21122 -8927
rect 21122 -8953 21148 -8927
rect 21148 -8953 21149 -8927
rect 21121 -8954 21149 -8953
rect 21121 -9087 21149 -9086
rect 21121 -9113 21122 -9087
rect 21122 -9113 21148 -9087
rect 21148 -9113 21149 -9087
rect 21121 -9114 21149 -9113
rect 24854 -5887 24882 -5886
rect 24854 -5913 24855 -5887
rect 24855 -5913 24881 -5887
rect 24881 -5913 24882 -5887
rect 24854 -5914 24882 -5913
rect 24854 -6047 24882 -6046
rect 24854 -6073 24855 -6047
rect 24855 -6073 24881 -6047
rect 24881 -6073 24882 -6047
rect 24854 -6074 24882 -6073
rect 24854 -6207 24882 -6206
rect 24854 -6233 24855 -6207
rect 24855 -6233 24881 -6207
rect 24881 -6233 24882 -6207
rect 24854 -6234 24882 -6233
rect 24854 -6367 24882 -6366
rect 24854 -6393 24855 -6367
rect 24855 -6393 24881 -6367
rect 24881 -6393 24882 -6367
rect 24854 -6394 24882 -6393
rect 24854 -6527 24882 -6526
rect 24854 -6553 24855 -6527
rect 24855 -6553 24881 -6527
rect 24881 -6553 24882 -6527
rect 24854 -6554 24882 -6553
rect 24854 -6687 24882 -6686
rect 24854 -6713 24855 -6687
rect 24855 -6713 24881 -6687
rect 24881 -6713 24882 -6687
rect 24854 -6714 24882 -6713
rect 24854 -6847 24882 -6846
rect 24854 -6873 24855 -6847
rect 24855 -6873 24881 -6847
rect 24881 -6873 24882 -6847
rect 24854 -6874 24882 -6873
rect 24854 -7007 24882 -7006
rect 24854 -7033 24855 -7007
rect 24855 -7033 24881 -7007
rect 24881 -7033 24882 -7007
rect 24854 -7034 24882 -7033
rect 24854 -7167 24882 -7166
rect 24854 -7193 24855 -7167
rect 24855 -7193 24881 -7167
rect 24881 -7193 24882 -7167
rect 24854 -7194 24882 -7193
rect 24854 -7327 24882 -7326
rect 24854 -7353 24855 -7327
rect 24855 -7353 24881 -7327
rect 24881 -7353 24882 -7327
rect 24854 -7354 24882 -7353
rect 24854 -7487 24882 -7486
rect 24854 -7513 24855 -7487
rect 24855 -7513 24881 -7487
rect 24881 -7513 24882 -7487
rect 24854 -7514 24882 -7513
rect 24854 -7647 24882 -7646
rect 24854 -7673 24855 -7647
rect 24855 -7673 24881 -7647
rect 24881 -7673 24882 -7647
rect 24854 -7674 24882 -7673
rect 24854 -7807 24882 -7806
rect 24854 -7833 24855 -7807
rect 24855 -7833 24881 -7807
rect 24881 -7833 24882 -7807
rect 24854 -7834 24882 -7833
rect 24854 -7967 24882 -7966
rect 24854 -7993 24855 -7967
rect 24855 -7993 24881 -7967
rect 24881 -7993 24882 -7967
rect 24854 -7994 24882 -7993
rect 24854 -8127 24882 -8126
rect 24854 -8153 24855 -8127
rect 24855 -8153 24881 -8127
rect 24881 -8153 24882 -8127
rect 24854 -8154 24882 -8153
rect 24854 -8287 24882 -8286
rect 24854 -8313 24855 -8287
rect 24855 -8313 24881 -8287
rect 24881 -8313 24882 -8287
rect 24854 -8314 24882 -8313
rect 24854 -8447 24882 -8446
rect 24854 -8473 24855 -8447
rect 24855 -8473 24881 -8447
rect 24881 -8473 24882 -8447
rect 24854 -8474 24882 -8473
rect 24854 -8607 24882 -8606
rect 24854 -8633 24855 -8607
rect 24855 -8633 24881 -8607
rect 24881 -8633 24882 -8607
rect 24854 -8634 24882 -8633
rect 24854 -8767 24882 -8766
rect 24854 -8793 24855 -8767
rect 24855 -8793 24881 -8767
rect 24881 -8793 24882 -8767
rect 24854 -8794 24882 -8793
rect 24854 -8927 24882 -8926
rect 24854 -8953 24855 -8927
rect 24855 -8953 24881 -8927
rect 24881 -8953 24882 -8927
rect 24854 -8954 24882 -8953
rect 24854 -9087 24882 -9086
rect 24854 -9113 24855 -9087
rect 24855 -9113 24881 -9087
rect 24881 -9113 24882 -9087
rect 24854 -9114 24882 -9113
rect 21121 -9247 21149 -9246
rect 21121 -9273 21122 -9247
rect 21122 -9273 21148 -9247
rect 21148 -9273 21149 -9247
rect 21121 -9274 21149 -9273
rect 24854 -9247 24882 -9246
rect 24854 -9273 24855 -9247
rect 24855 -9273 24881 -9247
rect 24881 -9273 24882 -9247
rect 24854 -9274 24882 -9273
rect 21306 -9352 21334 -9351
rect 21306 -9378 21307 -9352
rect 21307 -9378 21333 -9352
rect 21333 -9378 21334 -9352
rect 21306 -9379 21334 -9378
rect 21466 -9352 21494 -9351
rect 21466 -9378 21467 -9352
rect 21467 -9378 21493 -9352
rect 21493 -9378 21494 -9352
rect 21466 -9379 21494 -9378
rect 21626 -9352 21654 -9351
rect 21626 -9378 21627 -9352
rect 21627 -9378 21653 -9352
rect 21653 -9378 21654 -9352
rect 21626 -9379 21654 -9378
rect 21786 -9352 21814 -9351
rect 21786 -9378 21787 -9352
rect 21787 -9378 21813 -9352
rect 21813 -9378 21814 -9352
rect 21786 -9379 21814 -9378
rect 21946 -9352 21974 -9351
rect 21946 -9378 21947 -9352
rect 21947 -9378 21973 -9352
rect 21973 -9378 21974 -9352
rect 21946 -9379 21974 -9378
rect 22106 -9352 22134 -9351
rect 22106 -9378 22107 -9352
rect 22107 -9378 22133 -9352
rect 22133 -9378 22134 -9352
rect 22106 -9379 22134 -9378
rect 22266 -9352 22294 -9351
rect 22266 -9378 22267 -9352
rect 22267 -9378 22293 -9352
rect 22293 -9378 22294 -9352
rect 22266 -9379 22294 -9378
rect 22426 -9352 22454 -9351
rect 22426 -9378 22427 -9352
rect 22427 -9378 22453 -9352
rect 22453 -9378 22454 -9352
rect 22426 -9379 22454 -9378
rect 22586 -9352 22614 -9351
rect 22586 -9378 22587 -9352
rect 22587 -9378 22613 -9352
rect 22613 -9378 22614 -9352
rect 22586 -9379 22614 -9378
rect 22746 -9352 22774 -9351
rect 22746 -9378 22747 -9352
rect 22747 -9378 22773 -9352
rect 22773 -9378 22774 -9352
rect 22746 -9379 22774 -9378
rect 22906 -9352 22934 -9351
rect 22906 -9378 22907 -9352
rect 22907 -9378 22933 -9352
rect 22933 -9378 22934 -9352
rect 22906 -9379 22934 -9378
rect 23066 -9352 23094 -9351
rect 23066 -9378 23067 -9352
rect 23067 -9378 23093 -9352
rect 23093 -9378 23094 -9352
rect 23066 -9379 23094 -9378
rect 23226 -9352 23254 -9351
rect 23226 -9378 23227 -9352
rect 23227 -9378 23253 -9352
rect 23253 -9378 23254 -9352
rect 23226 -9379 23254 -9378
rect 23386 -9352 23414 -9351
rect 23386 -9378 23387 -9352
rect 23387 -9378 23413 -9352
rect 23413 -9378 23414 -9352
rect 23386 -9379 23414 -9378
rect 23546 -9352 23574 -9351
rect 23546 -9378 23547 -9352
rect 23547 -9378 23573 -9352
rect 23573 -9378 23574 -9352
rect 23546 -9379 23574 -9378
rect 23706 -9352 23734 -9351
rect 23706 -9378 23707 -9352
rect 23707 -9378 23733 -9352
rect 23733 -9378 23734 -9352
rect 23706 -9379 23734 -9378
rect 23866 -9352 23894 -9351
rect 23866 -9378 23867 -9352
rect 23867 -9378 23893 -9352
rect 23893 -9378 23894 -9352
rect 23866 -9379 23894 -9378
rect 24026 -9352 24054 -9351
rect 24026 -9378 24027 -9352
rect 24027 -9378 24053 -9352
rect 24053 -9378 24054 -9352
rect 24026 -9379 24054 -9378
rect 24186 -9352 24214 -9351
rect 24186 -9378 24187 -9352
rect 24187 -9378 24213 -9352
rect 24213 -9378 24214 -9352
rect 24186 -9379 24214 -9378
rect 24346 -9352 24374 -9351
rect 24346 -9378 24347 -9352
rect 24347 -9378 24373 -9352
rect 24373 -9378 24374 -9352
rect 24346 -9379 24374 -9378
rect 24506 -9352 24534 -9351
rect 24506 -9378 24507 -9352
rect 24507 -9378 24533 -9352
rect 24533 -9378 24534 -9352
rect 24506 -9379 24534 -9378
rect 24666 -9352 24694 -9351
rect 24666 -9378 24667 -9352
rect 24667 -9378 24693 -9352
rect 24693 -9378 24694 -9352
rect 24666 -9379 24694 -9378
rect 3306 -11624 3334 -11623
rect 3306 -11650 3307 -11624
rect 3307 -11650 3333 -11624
rect 3333 -11650 3334 -11624
rect 3306 -11651 3334 -11650
rect 3466 -11624 3494 -11623
rect 3466 -11650 3467 -11624
rect 3467 -11650 3493 -11624
rect 3493 -11650 3494 -11624
rect 3466 -11651 3494 -11650
rect 3626 -11624 3654 -11623
rect 3626 -11650 3627 -11624
rect 3627 -11650 3653 -11624
rect 3653 -11650 3654 -11624
rect 3626 -11651 3654 -11650
rect 3786 -11624 3814 -11623
rect 3786 -11650 3787 -11624
rect 3787 -11650 3813 -11624
rect 3813 -11650 3814 -11624
rect 3786 -11651 3814 -11650
rect 3946 -11624 3974 -11623
rect 3946 -11650 3947 -11624
rect 3947 -11650 3973 -11624
rect 3973 -11650 3974 -11624
rect 3946 -11651 3974 -11650
rect 4106 -11624 4134 -11623
rect 4106 -11650 4107 -11624
rect 4107 -11650 4133 -11624
rect 4133 -11650 4134 -11624
rect 4106 -11651 4134 -11650
rect 4266 -11624 4294 -11623
rect 4266 -11650 4267 -11624
rect 4267 -11650 4293 -11624
rect 4293 -11650 4294 -11624
rect 4266 -11651 4294 -11650
rect 4426 -11624 4454 -11623
rect 4426 -11650 4427 -11624
rect 4427 -11650 4453 -11624
rect 4453 -11650 4454 -11624
rect 4426 -11651 4454 -11650
rect 4586 -11624 4614 -11623
rect 4586 -11650 4587 -11624
rect 4587 -11650 4613 -11624
rect 4613 -11650 4614 -11624
rect 4586 -11651 4614 -11650
rect 4746 -11624 4774 -11623
rect 4746 -11650 4747 -11624
rect 4747 -11650 4773 -11624
rect 4773 -11650 4774 -11624
rect 4746 -11651 4774 -11650
rect 4906 -11624 4934 -11623
rect 4906 -11650 4907 -11624
rect 4907 -11650 4933 -11624
rect 4933 -11650 4934 -11624
rect 4906 -11651 4934 -11650
rect 5066 -11624 5094 -11623
rect 5066 -11650 5067 -11624
rect 5067 -11650 5093 -11624
rect 5093 -11650 5094 -11624
rect 5066 -11651 5094 -11650
rect 5226 -11624 5254 -11623
rect 5226 -11650 5227 -11624
rect 5227 -11650 5253 -11624
rect 5253 -11650 5254 -11624
rect 5226 -11651 5254 -11650
rect 5386 -11624 5414 -11623
rect 5386 -11650 5387 -11624
rect 5387 -11650 5413 -11624
rect 5413 -11650 5414 -11624
rect 5386 -11651 5414 -11650
rect 5546 -11624 5574 -11623
rect 5546 -11650 5547 -11624
rect 5547 -11650 5573 -11624
rect 5573 -11650 5574 -11624
rect 5546 -11651 5574 -11650
rect 5706 -11624 5734 -11623
rect 5706 -11650 5707 -11624
rect 5707 -11650 5733 -11624
rect 5733 -11650 5734 -11624
rect 5706 -11651 5734 -11650
rect 5866 -11624 5894 -11623
rect 5866 -11650 5867 -11624
rect 5867 -11650 5893 -11624
rect 5893 -11650 5894 -11624
rect 5866 -11651 5894 -11650
rect 6026 -11624 6054 -11623
rect 6026 -11650 6027 -11624
rect 6027 -11650 6053 -11624
rect 6053 -11650 6054 -11624
rect 6026 -11651 6054 -11650
rect 6186 -11624 6214 -11623
rect 6186 -11650 6187 -11624
rect 6187 -11650 6213 -11624
rect 6213 -11650 6214 -11624
rect 6186 -11651 6214 -11650
rect 6346 -11624 6374 -11623
rect 6346 -11650 6347 -11624
rect 6347 -11650 6373 -11624
rect 6373 -11650 6374 -11624
rect 6346 -11651 6374 -11650
rect 6506 -11624 6534 -11623
rect 6506 -11650 6507 -11624
rect 6507 -11650 6533 -11624
rect 6533 -11650 6534 -11624
rect 6506 -11651 6534 -11650
rect 6666 -11624 6694 -11623
rect 6666 -11650 6667 -11624
rect 6667 -11650 6693 -11624
rect 6693 -11650 6694 -11624
rect 6666 -11651 6694 -11650
rect 3121 -11727 3149 -11726
rect 3121 -11753 3122 -11727
rect 3122 -11753 3148 -11727
rect 3148 -11753 3149 -11727
rect 3121 -11754 3149 -11753
rect 6854 -11727 6882 -11726
rect 6854 -11753 6855 -11727
rect 6855 -11753 6881 -11727
rect 6881 -11753 6882 -11727
rect 6854 -11754 6882 -11753
rect 3121 -11887 3149 -11886
rect 3121 -11913 3122 -11887
rect 3122 -11913 3148 -11887
rect 3148 -11913 3149 -11887
rect 3121 -11914 3149 -11913
rect 3121 -12047 3149 -12046
rect 3121 -12073 3122 -12047
rect 3122 -12073 3148 -12047
rect 3148 -12073 3149 -12047
rect 3121 -12074 3149 -12073
rect 3121 -12207 3149 -12206
rect 3121 -12233 3122 -12207
rect 3122 -12233 3148 -12207
rect 3148 -12233 3149 -12207
rect 3121 -12234 3149 -12233
rect 3121 -12367 3149 -12366
rect 3121 -12393 3122 -12367
rect 3122 -12393 3148 -12367
rect 3148 -12393 3149 -12367
rect 3121 -12394 3149 -12393
rect 3121 -12527 3149 -12526
rect 3121 -12553 3122 -12527
rect 3122 -12553 3148 -12527
rect 3148 -12553 3149 -12527
rect 3121 -12554 3149 -12553
rect 3121 -12687 3149 -12686
rect 3121 -12713 3122 -12687
rect 3122 -12713 3148 -12687
rect 3148 -12713 3149 -12687
rect 3121 -12714 3149 -12713
rect 3121 -12847 3149 -12846
rect 3121 -12873 3122 -12847
rect 3122 -12873 3148 -12847
rect 3148 -12873 3149 -12847
rect 3121 -12874 3149 -12873
rect 3121 -13007 3149 -13006
rect 3121 -13033 3122 -13007
rect 3122 -13033 3148 -13007
rect 3148 -13033 3149 -13007
rect 3121 -13034 3149 -13033
rect 3121 -13167 3149 -13166
rect 3121 -13193 3122 -13167
rect 3122 -13193 3148 -13167
rect 3148 -13193 3149 -13167
rect 3121 -13194 3149 -13193
rect 3121 -13327 3149 -13326
rect 3121 -13353 3122 -13327
rect 3122 -13353 3148 -13327
rect 3148 -13353 3149 -13327
rect 3121 -13354 3149 -13353
rect 3121 -13487 3149 -13486
rect 3121 -13513 3122 -13487
rect 3122 -13513 3148 -13487
rect 3148 -13513 3149 -13487
rect 3121 -13514 3149 -13513
rect 3121 -13647 3149 -13646
rect 3121 -13673 3122 -13647
rect 3122 -13673 3148 -13647
rect 3148 -13673 3149 -13647
rect 3121 -13674 3149 -13673
rect 3121 -13807 3149 -13806
rect 3121 -13833 3122 -13807
rect 3122 -13833 3148 -13807
rect 3148 -13833 3149 -13807
rect 3121 -13834 3149 -13833
rect 3121 -13967 3149 -13966
rect 3121 -13993 3122 -13967
rect 3122 -13993 3148 -13967
rect 3148 -13993 3149 -13967
rect 3121 -13994 3149 -13993
rect 3121 -14127 3149 -14126
rect 3121 -14153 3122 -14127
rect 3122 -14153 3148 -14127
rect 3148 -14153 3149 -14127
rect 3121 -14154 3149 -14153
rect 3121 -14287 3149 -14286
rect 3121 -14313 3122 -14287
rect 3122 -14313 3148 -14287
rect 3148 -14313 3149 -14287
rect 3121 -14314 3149 -14313
rect 3121 -14447 3149 -14446
rect 3121 -14473 3122 -14447
rect 3122 -14473 3148 -14447
rect 3148 -14473 3149 -14447
rect 3121 -14474 3149 -14473
rect 3121 -14607 3149 -14606
rect 3121 -14633 3122 -14607
rect 3122 -14633 3148 -14607
rect 3148 -14633 3149 -14607
rect 3121 -14634 3149 -14633
rect 3121 -14767 3149 -14766
rect 3121 -14793 3122 -14767
rect 3122 -14793 3148 -14767
rect 3148 -14793 3149 -14767
rect 3121 -14794 3149 -14793
rect 3121 -14927 3149 -14926
rect 3121 -14953 3122 -14927
rect 3122 -14953 3148 -14927
rect 3148 -14953 3149 -14927
rect 3121 -14954 3149 -14953
rect 3121 -15087 3149 -15086
rect 3121 -15113 3122 -15087
rect 3122 -15113 3148 -15087
rect 3148 -15113 3149 -15087
rect 3121 -15114 3149 -15113
rect 6854 -11887 6882 -11886
rect 6854 -11913 6855 -11887
rect 6855 -11913 6881 -11887
rect 6881 -11913 6882 -11887
rect 6854 -11914 6882 -11913
rect 6854 -12047 6882 -12046
rect 6854 -12073 6855 -12047
rect 6855 -12073 6881 -12047
rect 6881 -12073 6882 -12047
rect 6854 -12074 6882 -12073
rect 6854 -12207 6882 -12206
rect 6854 -12233 6855 -12207
rect 6855 -12233 6881 -12207
rect 6881 -12233 6882 -12207
rect 6854 -12234 6882 -12233
rect 6854 -12367 6882 -12366
rect 6854 -12393 6855 -12367
rect 6855 -12393 6881 -12367
rect 6881 -12393 6882 -12367
rect 6854 -12394 6882 -12393
rect 6854 -12527 6882 -12526
rect 6854 -12553 6855 -12527
rect 6855 -12553 6881 -12527
rect 6881 -12553 6882 -12527
rect 6854 -12554 6882 -12553
rect 6854 -12687 6882 -12686
rect 6854 -12713 6855 -12687
rect 6855 -12713 6881 -12687
rect 6881 -12713 6882 -12687
rect 6854 -12714 6882 -12713
rect 6854 -12847 6882 -12846
rect 6854 -12873 6855 -12847
rect 6855 -12873 6881 -12847
rect 6881 -12873 6882 -12847
rect 6854 -12874 6882 -12873
rect 6854 -13007 6882 -13006
rect 6854 -13033 6855 -13007
rect 6855 -13033 6881 -13007
rect 6881 -13033 6882 -13007
rect 6854 -13034 6882 -13033
rect 6854 -13167 6882 -13166
rect 6854 -13193 6855 -13167
rect 6855 -13193 6881 -13167
rect 6881 -13193 6882 -13167
rect 6854 -13194 6882 -13193
rect 6854 -13327 6882 -13326
rect 6854 -13353 6855 -13327
rect 6855 -13353 6881 -13327
rect 6881 -13353 6882 -13327
rect 6854 -13354 6882 -13353
rect 6854 -13487 6882 -13486
rect 6854 -13513 6855 -13487
rect 6855 -13513 6881 -13487
rect 6881 -13513 6882 -13487
rect 6854 -13514 6882 -13513
rect 6854 -13647 6882 -13646
rect 6854 -13673 6855 -13647
rect 6855 -13673 6881 -13647
rect 6881 -13673 6882 -13647
rect 6854 -13674 6882 -13673
rect 6854 -13807 6882 -13806
rect 6854 -13833 6855 -13807
rect 6855 -13833 6881 -13807
rect 6881 -13833 6882 -13807
rect 6854 -13834 6882 -13833
rect 6854 -13967 6882 -13966
rect 6854 -13993 6855 -13967
rect 6855 -13993 6881 -13967
rect 6881 -13993 6882 -13967
rect 6854 -13994 6882 -13993
rect 6854 -14127 6882 -14126
rect 6854 -14153 6855 -14127
rect 6855 -14153 6881 -14127
rect 6881 -14153 6882 -14127
rect 6854 -14154 6882 -14153
rect 6854 -14287 6882 -14286
rect 6854 -14313 6855 -14287
rect 6855 -14313 6881 -14287
rect 6881 -14313 6882 -14287
rect 6854 -14314 6882 -14313
rect 6854 -14447 6882 -14446
rect 6854 -14473 6855 -14447
rect 6855 -14473 6881 -14447
rect 6881 -14473 6882 -14447
rect 6854 -14474 6882 -14473
rect 6854 -14607 6882 -14606
rect 6854 -14633 6855 -14607
rect 6855 -14633 6881 -14607
rect 6881 -14633 6882 -14607
rect 6854 -14634 6882 -14633
rect 6854 -14767 6882 -14766
rect 6854 -14793 6855 -14767
rect 6855 -14793 6881 -14767
rect 6881 -14793 6882 -14767
rect 6854 -14794 6882 -14793
rect 6854 -14927 6882 -14926
rect 6854 -14953 6855 -14927
rect 6855 -14953 6881 -14927
rect 6881 -14953 6882 -14927
rect 6854 -14954 6882 -14953
rect 6854 -15087 6882 -15086
rect 6854 -15113 6855 -15087
rect 6855 -15113 6881 -15087
rect 6881 -15113 6882 -15087
rect 6854 -15114 6882 -15113
rect 3121 -15247 3149 -15246
rect 3121 -15273 3122 -15247
rect 3122 -15273 3148 -15247
rect 3148 -15273 3149 -15247
rect 3121 -15274 3149 -15273
rect 6854 -15247 6882 -15246
rect 6854 -15273 6855 -15247
rect 6855 -15273 6881 -15247
rect 6881 -15273 6882 -15247
rect 6854 -15274 6882 -15273
rect 3306 -15352 3334 -15351
rect 3306 -15378 3307 -15352
rect 3307 -15378 3333 -15352
rect 3333 -15378 3334 -15352
rect 3306 -15379 3334 -15378
rect 3466 -15352 3494 -15351
rect 3466 -15378 3467 -15352
rect 3467 -15378 3493 -15352
rect 3493 -15378 3494 -15352
rect 3466 -15379 3494 -15378
rect 3626 -15352 3654 -15351
rect 3626 -15378 3627 -15352
rect 3627 -15378 3653 -15352
rect 3653 -15378 3654 -15352
rect 3626 -15379 3654 -15378
rect 3786 -15352 3814 -15351
rect 3786 -15378 3787 -15352
rect 3787 -15378 3813 -15352
rect 3813 -15378 3814 -15352
rect 3786 -15379 3814 -15378
rect 3946 -15352 3974 -15351
rect 3946 -15378 3947 -15352
rect 3947 -15378 3973 -15352
rect 3973 -15378 3974 -15352
rect 3946 -15379 3974 -15378
rect 4106 -15352 4134 -15351
rect 4106 -15378 4107 -15352
rect 4107 -15378 4133 -15352
rect 4133 -15378 4134 -15352
rect 4106 -15379 4134 -15378
rect 4266 -15352 4294 -15351
rect 4266 -15378 4267 -15352
rect 4267 -15378 4293 -15352
rect 4293 -15378 4294 -15352
rect 4266 -15379 4294 -15378
rect 4426 -15352 4454 -15351
rect 4426 -15378 4427 -15352
rect 4427 -15378 4453 -15352
rect 4453 -15378 4454 -15352
rect 4426 -15379 4454 -15378
rect 4586 -15352 4614 -15351
rect 4586 -15378 4587 -15352
rect 4587 -15378 4613 -15352
rect 4613 -15378 4614 -15352
rect 4586 -15379 4614 -15378
rect 4746 -15352 4774 -15351
rect 4746 -15378 4747 -15352
rect 4747 -15378 4773 -15352
rect 4773 -15378 4774 -15352
rect 4746 -15379 4774 -15378
rect 4906 -15352 4934 -15351
rect 4906 -15378 4907 -15352
rect 4907 -15378 4933 -15352
rect 4933 -15378 4934 -15352
rect 4906 -15379 4934 -15378
rect 5066 -15352 5094 -15351
rect 5066 -15378 5067 -15352
rect 5067 -15378 5093 -15352
rect 5093 -15378 5094 -15352
rect 5066 -15379 5094 -15378
rect 5226 -15352 5254 -15351
rect 5226 -15378 5227 -15352
rect 5227 -15378 5253 -15352
rect 5253 -15378 5254 -15352
rect 5226 -15379 5254 -15378
rect 5386 -15352 5414 -15351
rect 5386 -15378 5387 -15352
rect 5387 -15378 5413 -15352
rect 5413 -15378 5414 -15352
rect 5386 -15379 5414 -15378
rect 5546 -15352 5574 -15351
rect 5546 -15378 5547 -15352
rect 5547 -15378 5573 -15352
rect 5573 -15378 5574 -15352
rect 5546 -15379 5574 -15378
rect 5706 -15352 5734 -15351
rect 5706 -15378 5707 -15352
rect 5707 -15378 5733 -15352
rect 5733 -15378 5734 -15352
rect 5706 -15379 5734 -15378
rect 5866 -15352 5894 -15351
rect 5866 -15378 5867 -15352
rect 5867 -15378 5893 -15352
rect 5893 -15378 5894 -15352
rect 5866 -15379 5894 -15378
rect 6026 -15352 6054 -15351
rect 6026 -15378 6027 -15352
rect 6027 -15378 6053 -15352
rect 6053 -15378 6054 -15352
rect 6026 -15379 6054 -15378
rect 6186 -15352 6214 -15351
rect 6186 -15378 6187 -15352
rect 6187 -15378 6213 -15352
rect 6213 -15378 6214 -15352
rect 6186 -15379 6214 -15378
rect 6346 -15352 6374 -15351
rect 6346 -15378 6347 -15352
rect 6347 -15378 6373 -15352
rect 6373 -15378 6374 -15352
rect 6346 -15379 6374 -15378
rect 6506 -15352 6534 -15351
rect 6506 -15378 6507 -15352
rect 6507 -15378 6533 -15352
rect 6533 -15378 6534 -15352
rect 6506 -15379 6534 -15378
rect 6666 -15352 6694 -15351
rect 6666 -15378 6667 -15352
rect 6667 -15378 6693 -15352
rect 6693 -15378 6694 -15352
rect 6666 -15379 6694 -15378
rect 9306 -11624 9334 -11623
rect 9306 -11650 9307 -11624
rect 9307 -11650 9333 -11624
rect 9333 -11650 9334 -11624
rect 9306 -11651 9334 -11650
rect 9466 -11624 9494 -11623
rect 9466 -11650 9467 -11624
rect 9467 -11650 9493 -11624
rect 9493 -11650 9494 -11624
rect 9466 -11651 9494 -11650
rect 9626 -11624 9654 -11623
rect 9626 -11650 9627 -11624
rect 9627 -11650 9653 -11624
rect 9653 -11650 9654 -11624
rect 9626 -11651 9654 -11650
rect 9786 -11624 9814 -11623
rect 9786 -11650 9787 -11624
rect 9787 -11650 9813 -11624
rect 9813 -11650 9814 -11624
rect 9786 -11651 9814 -11650
rect 9946 -11624 9974 -11623
rect 9946 -11650 9947 -11624
rect 9947 -11650 9973 -11624
rect 9973 -11650 9974 -11624
rect 9946 -11651 9974 -11650
rect 10106 -11624 10134 -11623
rect 10106 -11650 10107 -11624
rect 10107 -11650 10133 -11624
rect 10133 -11650 10134 -11624
rect 10106 -11651 10134 -11650
rect 10266 -11624 10294 -11623
rect 10266 -11650 10267 -11624
rect 10267 -11650 10293 -11624
rect 10293 -11650 10294 -11624
rect 10266 -11651 10294 -11650
rect 10426 -11624 10454 -11623
rect 10426 -11650 10427 -11624
rect 10427 -11650 10453 -11624
rect 10453 -11650 10454 -11624
rect 10426 -11651 10454 -11650
rect 10586 -11624 10614 -11623
rect 10586 -11650 10587 -11624
rect 10587 -11650 10613 -11624
rect 10613 -11650 10614 -11624
rect 10586 -11651 10614 -11650
rect 10746 -11624 10774 -11623
rect 10746 -11650 10747 -11624
rect 10747 -11650 10773 -11624
rect 10773 -11650 10774 -11624
rect 10746 -11651 10774 -11650
rect 10906 -11624 10934 -11623
rect 10906 -11650 10907 -11624
rect 10907 -11650 10933 -11624
rect 10933 -11650 10934 -11624
rect 10906 -11651 10934 -11650
rect 11066 -11624 11094 -11623
rect 11066 -11650 11067 -11624
rect 11067 -11650 11093 -11624
rect 11093 -11650 11094 -11624
rect 11066 -11651 11094 -11650
rect 11226 -11624 11254 -11623
rect 11226 -11650 11227 -11624
rect 11227 -11650 11253 -11624
rect 11253 -11650 11254 -11624
rect 11226 -11651 11254 -11650
rect 11386 -11624 11414 -11623
rect 11386 -11650 11387 -11624
rect 11387 -11650 11413 -11624
rect 11413 -11650 11414 -11624
rect 11386 -11651 11414 -11650
rect 11546 -11624 11574 -11623
rect 11546 -11650 11547 -11624
rect 11547 -11650 11573 -11624
rect 11573 -11650 11574 -11624
rect 11546 -11651 11574 -11650
rect 11706 -11624 11734 -11623
rect 11706 -11650 11707 -11624
rect 11707 -11650 11733 -11624
rect 11733 -11650 11734 -11624
rect 11706 -11651 11734 -11650
rect 11866 -11624 11894 -11623
rect 11866 -11650 11867 -11624
rect 11867 -11650 11893 -11624
rect 11893 -11650 11894 -11624
rect 11866 -11651 11894 -11650
rect 12026 -11624 12054 -11623
rect 12026 -11650 12027 -11624
rect 12027 -11650 12053 -11624
rect 12053 -11650 12054 -11624
rect 12026 -11651 12054 -11650
rect 12186 -11624 12214 -11623
rect 12186 -11650 12187 -11624
rect 12187 -11650 12213 -11624
rect 12213 -11650 12214 -11624
rect 12186 -11651 12214 -11650
rect 12346 -11624 12374 -11623
rect 12346 -11650 12347 -11624
rect 12347 -11650 12373 -11624
rect 12373 -11650 12374 -11624
rect 12346 -11651 12374 -11650
rect 12506 -11624 12534 -11623
rect 12506 -11650 12507 -11624
rect 12507 -11650 12533 -11624
rect 12533 -11650 12534 -11624
rect 12506 -11651 12534 -11650
rect 12666 -11624 12694 -11623
rect 12666 -11650 12667 -11624
rect 12667 -11650 12693 -11624
rect 12693 -11650 12694 -11624
rect 12666 -11651 12694 -11650
rect 9121 -11727 9149 -11726
rect 9121 -11753 9122 -11727
rect 9122 -11753 9148 -11727
rect 9148 -11753 9149 -11727
rect 9121 -11754 9149 -11753
rect 12854 -11727 12882 -11726
rect 12854 -11753 12855 -11727
rect 12855 -11753 12881 -11727
rect 12881 -11753 12882 -11727
rect 12854 -11754 12882 -11753
rect 9121 -11887 9149 -11886
rect 9121 -11913 9122 -11887
rect 9122 -11913 9148 -11887
rect 9148 -11913 9149 -11887
rect 9121 -11914 9149 -11913
rect 9121 -12047 9149 -12046
rect 9121 -12073 9122 -12047
rect 9122 -12073 9148 -12047
rect 9148 -12073 9149 -12047
rect 9121 -12074 9149 -12073
rect 9121 -12207 9149 -12206
rect 9121 -12233 9122 -12207
rect 9122 -12233 9148 -12207
rect 9148 -12233 9149 -12207
rect 9121 -12234 9149 -12233
rect 9121 -12367 9149 -12366
rect 9121 -12393 9122 -12367
rect 9122 -12393 9148 -12367
rect 9148 -12393 9149 -12367
rect 9121 -12394 9149 -12393
rect 9121 -12527 9149 -12526
rect 9121 -12553 9122 -12527
rect 9122 -12553 9148 -12527
rect 9148 -12553 9149 -12527
rect 9121 -12554 9149 -12553
rect 9121 -12687 9149 -12686
rect 9121 -12713 9122 -12687
rect 9122 -12713 9148 -12687
rect 9148 -12713 9149 -12687
rect 9121 -12714 9149 -12713
rect 9121 -12847 9149 -12846
rect 9121 -12873 9122 -12847
rect 9122 -12873 9148 -12847
rect 9148 -12873 9149 -12847
rect 9121 -12874 9149 -12873
rect 9121 -13007 9149 -13006
rect 9121 -13033 9122 -13007
rect 9122 -13033 9148 -13007
rect 9148 -13033 9149 -13007
rect 9121 -13034 9149 -13033
rect 9121 -13167 9149 -13166
rect 9121 -13193 9122 -13167
rect 9122 -13193 9148 -13167
rect 9148 -13193 9149 -13167
rect 9121 -13194 9149 -13193
rect 9121 -13327 9149 -13326
rect 9121 -13353 9122 -13327
rect 9122 -13353 9148 -13327
rect 9148 -13353 9149 -13327
rect 9121 -13354 9149 -13353
rect 9121 -13487 9149 -13486
rect 9121 -13513 9122 -13487
rect 9122 -13513 9148 -13487
rect 9148 -13513 9149 -13487
rect 9121 -13514 9149 -13513
rect 9121 -13647 9149 -13646
rect 9121 -13673 9122 -13647
rect 9122 -13673 9148 -13647
rect 9148 -13673 9149 -13647
rect 9121 -13674 9149 -13673
rect 9121 -13807 9149 -13806
rect 9121 -13833 9122 -13807
rect 9122 -13833 9148 -13807
rect 9148 -13833 9149 -13807
rect 9121 -13834 9149 -13833
rect 9121 -13967 9149 -13966
rect 9121 -13993 9122 -13967
rect 9122 -13993 9148 -13967
rect 9148 -13993 9149 -13967
rect 9121 -13994 9149 -13993
rect 9121 -14127 9149 -14126
rect 9121 -14153 9122 -14127
rect 9122 -14153 9148 -14127
rect 9148 -14153 9149 -14127
rect 9121 -14154 9149 -14153
rect 9121 -14287 9149 -14286
rect 9121 -14313 9122 -14287
rect 9122 -14313 9148 -14287
rect 9148 -14313 9149 -14287
rect 9121 -14314 9149 -14313
rect 9121 -14447 9149 -14446
rect 9121 -14473 9122 -14447
rect 9122 -14473 9148 -14447
rect 9148 -14473 9149 -14447
rect 9121 -14474 9149 -14473
rect 9121 -14607 9149 -14606
rect 9121 -14633 9122 -14607
rect 9122 -14633 9148 -14607
rect 9148 -14633 9149 -14607
rect 9121 -14634 9149 -14633
rect 9121 -14767 9149 -14766
rect 9121 -14793 9122 -14767
rect 9122 -14793 9148 -14767
rect 9148 -14793 9149 -14767
rect 9121 -14794 9149 -14793
rect 9121 -14927 9149 -14926
rect 9121 -14953 9122 -14927
rect 9122 -14953 9148 -14927
rect 9148 -14953 9149 -14927
rect 9121 -14954 9149 -14953
rect 9121 -15087 9149 -15086
rect 9121 -15113 9122 -15087
rect 9122 -15113 9148 -15087
rect 9148 -15113 9149 -15087
rect 9121 -15114 9149 -15113
rect 12854 -11887 12882 -11886
rect 12854 -11913 12855 -11887
rect 12855 -11913 12881 -11887
rect 12881 -11913 12882 -11887
rect 12854 -11914 12882 -11913
rect 12854 -12047 12882 -12046
rect 12854 -12073 12855 -12047
rect 12855 -12073 12881 -12047
rect 12881 -12073 12882 -12047
rect 12854 -12074 12882 -12073
rect 12854 -12207 12882 -12206
rect 12854 -12233 12855 -12207
rect 12855 -12233 12881 -12207
rect 12881 -12233 12882 -12207
rect 12854 -12234 12882 -12233
rect 12854 -12367 12882 -12366
rect 12854 -12393 12855 -12367
rect 12855 -12393 12881 -12367
rect 12881 -12393 12882 -12367
rect 12854 -12394 12882 -12393
rect 12854 -12527 12882 -12526
rect 12854 -12553 12855 -12527
rect 12855 -12553 12881 -12527
rect 12881 -12553 12882 -12527
rect 12854 -12554 12882 -12553
rect 12854 -12687 12882 -12686
rect 12854 -12713 12855 -12687
rect 12855 -12713 12881 -12687
rect 12881 -12713 12882 -12687
rect 12854 -12714 12882 -12713
rect 12854 -12847 12882 -12846
rect 12854 -12873 12855 -12847
rect 12855 -12873 12881 -12847
rect 12881 -12873 12882 -12847
rect 12854 -12874 12882 -12873
rect 12854 -13007 12882 -13006
rect 12854 -13033 12855 -13007
rect 12855 -13033 12881 -13007
rect 12881 -13033 12882 -13007
rect 12854 -13034 12882 -13033
rect 12854 -13167 12882 -13166
rect 12854 -13193 12855 -13167
rect 12855 -13193 12881 -13167
rect 12881 -13193 12882 -13167
rect 12854 -13194 12882 -13193
rect 12854 -13327 12882 -13326
rect 12854 -13353 12855 -13327
rect 12855 -13353 12881 -13327
rect 12881 -13353 12882 -13327
rect 12854 -13354 12882 -13353
rect 12854 -13487 12882 -13486
rect 12854 -13513 12855 -13487
rect 12855 -13513 12881 -13487
rect 12881 -13513 12882 -13487
rect 12854 -13514 12882 -13513
rect 12854 -13647 12882 -13646
rect 12854 -13673 12855 -13647
rect 12855 -13673 12881 -13647
rect 12881 -13673 12882 -13647
rect 12854 -13674 12882 -13673
rect 12854 -13807 12882 -13806
rect 12854 -13833 12855 -13807
rect 12855 -13833 12881 -13807
rect 12881 -13833 12882 -13807
rect 12854 -13834 12882 -13833
rect 12854 -13967 12882 -13966
rect 12854 -13993 12855 -13967
rect 12855 -13993 12881 -13967
rect 12881 -13993 12882 -13967
rect 12854 -13994 12882 -13993
rect 12854 -14127 12882 -14126
rect 12854 -14153 12855 -14127
rect 12855 -14153 12881 -14127
rect 12881 -14153 12882 -14127
rect 12854 -14154 12882 -14153
rect 12854 -14287 12882 -14286
rect 12854 -14313 12855 -14287
rect 12855 -14313 12881 -14287
rect 12881 -14313 12882 -14287
rect 12854 -14314 12882 -14313
rect 12854 -14447 12882 -14446
rect 12854 -14473 12855 -14447
rect 12855 -14473 12881 -14447
rect 12881 -14473 12882 -14447
rect 12854 -14474 12882 -14473
rect 12854 -14607 12882 -14606
rect 12854 -14633 12855 -14607
rect 12855 -14633 12881 -14607
rect 12881 -14633 12882 -14607
rect 12854 -14634 12882 -14633
rect 12854 -14767 12882 -14766
rect 12854 -14793 12855 -14767
rect 12855 -14793 12881 -14767
rect 12881 -14793 12882 -14767
rect 12854 -14794 12882 -14793
rect 12854 -14927 12882 -14926
rect 12854 -14953 12855 -14927
rect 12855 -14953 12881 -14927
rect 12881 -14953 12882 -14927
rect 12854 -14954 12882 -14953
rect 12854 -15087 12882 -15086
rect 12854 -15113 12855 -15087
rect 12855 -15113 12881 -15087
rect 12881 -15113 12882 -15087
rect 12854 -15114 12882 -15113
rect 9121 -15247 9149 -15246
rect 9121 -15273 9122 -15247
rect 9122 -15273 9148 -15247
rect 9148 -15273 9149 -15247
rect 9121 -15274 9149 -15273
rect 12854 -15247 12882 -15246
rect 12854 -15273 12855 -15247
rect 12855 -15273 12881 -15247
rect 12881 -15273 12882 -15247
rect 12854 -15274 12882 -15273
rect 9306 -15352 9334 -15351
rect 9306 -15378 9307 -15352
rect 9307 -15378 9333 -15352
rect 9333 -15378 9334 -15352
rect 9306 -15379 9334 -15378
rect 9466 -15352 9494 -15351
rect 9466 -15378 9467 -15352
rect 9467 -15378 9493 -15352
rect 9493 -15378 9494 -15352
rect 9466 -15379 9494 -15378
rect 9626 -15352 9654 -15351
rect 9626 -15378 9627 -15352
rect 9627 -15378 9653 -15352
rect 9653 -15378 9654 -15352
rect 9626 -15379 9654 -15378
rect 9786 -15352 9814 -15351
rect 9786 -15378 9787 -15352
rect 9787 -15378 9813 -15352
rect 9813 -15378 9814 -15352
rect 9786 -15379 9814 -15378
rect 9946 -15352 9974 -15351
rect 9946 -15378 9947 -15352
rect 9947 -15378 9973 -15352
rect 9973 -15378 9974 -15352
rect 9946 -15379 9974 -15378
rect 10106 -15352 10134 -15351
rect 10106 -15378 10107 -15352
rect 10107 -15378 10133 -15352
rect 10133 -15378 10134 -15352
rect 10106 -15379 10134 -15378
rect 10266 -15352 10294 -15351
rect 10266 -15378 10267 -15352
rect 10267 -15378 10293 -15352
rect 10293 -15378 10294 -15352
rect 10266 -15379 10294 -15378
rect 10426 -15352 10454 -15351
rect 10426 -15378 10427 -15352
rect 10427 -15378 10453 -15352
rect 10453 -15378 10454 -15352
rect 10426 -15379 10454 -15378
rect 10586 -15352 10614 -15351
rect 10586 -15378 10587 -15352
rect 10587 -15378 10613 -15352
rect 10613 -15378 10614 -15352
rect 10586 -15379 10614 -15378
rect 10746 -15352 10774 -15351
rect 10746 -15378 10747 -15352
rect 10747 -15378 10773 -15352
rect 10773 -15378 10774 -15352
rect 10746 -15379 10774 -15378
rect 10906 -15352 10934 -15351
rect 10906 -15378 10907 -15352
rect 10907 -15378 10933 -15352
rect 10933 -15378 10934 -15352
rect 10906 -15379 10934 -15378
rect 11066 -15352 11094 -15351
rect 11066 -15378 11067 -15352
rect 11067 -15378 11093 -15352
rect 11093 -15378 11094 -15352
rect 11066 -15379 11094 -15378
rect 11226 -15352 11254 -15351
rect 11226 -15378 11227 -15352
rect 11227 -15378 11253 -15352
rect 11253 -15378 11254 -15352
rect 11226 -15379 11254 -15378
rect 11386 -15352 11414 -15351
rect 11386 -15378 11387 -15352
rect 11387 -15378 11413 -15352
rect 11413 -15378 11414 -15352
rect 11386 -15379 11414 -15378
rect 11546 -15352 11574 -15351
rect 11546 -15378 11547 -15352
rect 11547 -15378 11573 -15352
rect 11573 -15378 11574 -15352
rect 11546 -15379 11574 -15378
rect 11706 -15352 11734 -15351
rect 11706 -15378 11707 -15352
rect 11707 -15378 11733 -15352
rect 11733 -15378 11734 -15352
rect 11706 -15379 11734 -15378
rect 11866 -15352 11894 -15351
rect 11866 -15378 11867 -15352
rect 11867 -15378 11893 -15352
rect 11893 -15378 11894 -15352
rect 11866 -15379 11894 -15378
rect 12026 -15352 12054 -15351
rect 12026 -15378 12027 -15352
rect 12027 -15378 12053 -15352
rect 12053 -15378 12054 -15352
rect 12026 -15379 12054 -15378
rect 12186 -15352 12214 -15351
rect 12186 -15378 12187 -15352
rect 12187 -15378 12213 -15352
rect 12213 -15378 12214 -15352
rect 12186 -15379 12214 -15378
rect 12346 -15352 12374 -15351
rect 12346 -15378 12347 -15352
rect 12347 -15378 12373 -15352
rect 12373 -15378 12374 -15352
rect 12346 -15379 12374 -15378
rect 12506 -15352 12534 -15351
rect 12506 -15378 12507 -15352
rect 12507 -15378 12533 -15352
rect 12533 -15378 12534 -15352
rect 12506 -15379 12534 -15378
rect 12666 -15352 12694 -15351
rect 12666 -15378 12667 -15352
rect 12667 -15378 12693 -15352
rect 12693 -15378 12694 -15352
rect 12666 -15379 12694 -15378
rect 15306 -11624 15334 -11623
rect 15306 -11650 15307 -11624
rect 15307 -11650 15333 -11624
rect 15333 -11650 15334 -11624
rect 15306 -11651 15334 -11650
rect 15466 -11624 15494 -11623
rect 15466 -11650 15467 -11624
rect 15467 -11650 15493 -11624
rect 15493 -11650 15494 -11624
rect 15466 -11651 15494 -11650
rect 15626 -11624 15654 -11623
rect 15626 -11650 15627 -11624
rect 15627 -11650 15653 -11624
rect 15653 -11650 15654 -11624
rect 15626 -11651 15654 -11650
rect 15786 -11624 15814 -11623
rect 15786 -11650 15787 -11624
rect 15787 -11650 15813 -11624
rect 15813 -11650 15814 -11624
rect 15786 -11651 15814 -11650
rect 15946 -11624 15974 -11623
rect 15946 -11650 15947 -11624
rect 15947 -11650 15973 -11624
rect 15973 -11650 15974 -11624
rect 15946 -11651 15974 -11650
rect 16106 -11624 16134 -11623
rect 16106 -11650 16107 -11624
rect 16107 -11650 16133 -11624
rect 16133 -11650 16134 -11624
rect 16106 -11651 16134 -11650
rect 16266 -11624 16294 -11623
rect 16266 -11650 16267 -11624
rect 16267 -11650 16293 -11624
rect 16293 -11650 16294 -11624
rect 16266 -11651 16294 -11650
rect 16426 -11624 16454 -11623
rect 16426 -11650 16427 -11624
rect 16427 -11650 16453 -11624
rect 16453 -11650 16454 -11624
rect 16426 -11651 16454 -11650
rect 16586 -11624 16614 -11623
rect 16586 -11650 16587 -11624
rect 16587 -11650 16613 -11624
rect 16613 -11650 16614 -11624
rect 16586 -11651 16614 -11650
rect 16746 -11624 16774 -11623
rect 16746 -11650 16747 -11624
rect 16747 -11650 16773 -11624
rect 16773 -11650 16774 -11624
rect 16746 -11651 16774 -11650
rect 16906 -11624 16934 -11623
rect 16906 -11650 16907 -11624
rect 16907 -11650 16933 -11624
rect 16933 -11650 16934 -11624
rect 16906 -11651 16934 -11650
rect 17066 -11624 17094 -11623
rect 17066 -11650 17067 -11624
rect 17067 -11650 17093 -11624
rect 17093 -11650 17094 -11624
rect 17066 -11651 17094 -11650
rect 17226 -11624 17254 -11623
rect 17226 -11650 17227 -11624
rect 17227 -11650 17253 -11624
rect 17253 -11650 17254 -11624
rect 17226 -11651 17254 -11650
rect 17386 -11624 17414 -11623
rect 17386 -11650 17387 -11624
rect 17387 -11650 17413 -11624
rect 17413 -11650 17414 -11624
rect 17386 -11651 17414 -11650
rect 17546 -11624 17574 -11623
rect 17546 -11650 17547 -11624
rect 17547 -11650 17573 -11624
rect 17573 -11650 17574 -11624
rect 17546 -11651 17574 -11650
rect 17706 -11624 17734 -11623
rect 17706 -11650 17707 -11624
rect 17707 -11650 17733 -11624
rect 17733 -11650 17734 -11624
rect 17706 -11651 17734 -11650
rect 17866 -11624 17894 -11623
rect 17866 -11650 17867 -11624
rect 17867 -11650 17893 -11624
rect 17893 -11650 17894 -11624
rect 17866 -11651 17894 -11650
rect 18026 -11624 18054 -11623
rect 18026 -11650 18027 -11624
rect 18027 -11650 18053 -11624
rect 18053 -11650 18054 -11624
rect 18026 -11651 18054 -11650
rect 18186 -11624 18214 -11623
rect 18186 -11650 18187 -11624
rect 18187 -11650 18213 -11624
rect 18213 -11650 18214 -11624
rect 18186 -11651 18214 -11650
rect 18346 -11624 18374 -11623
rect 18346 -11650 18347 -11624
rect 18347 -11650 18373 -11624
rect 18373 -11650 18374 -11624
rect 18346 -11651 18374 -11650
rect 18506 -11624 18534 -11623
rect 18506 -11650 18507 -11624
rect 18507 -11650 18533 -11624
rect 18533 -11650 18534 -11624
rect 18506 -11651 18534 -11650
rect 18666 -11624 18694 -11623
rect 18666 -11650 18667 -11624
rect 18667 -11650 18693 -11624
rect 18693 -11650 18694 -11624
rect 18666 -11651 18694 -11650
rect 15121 -11727 15149 -11726
rect 15121 -11753 15122 -11727
rect 15122 -11753 15148 -11727
rect 15148 -11753 15149 -11727
rect 15121 -11754 15149 -11753
rect 18854 -11727 18882 -11726
rect 18854 -11753 18855 -11727
rect 18855 -11753 18881 -11727
rect 18881 -11753 18882 -11727
rect 18854 -11754 18882 -11753
rect 15121 -11887 15149 -11886
rect 15121 -11913 15122 -11887
rect 15122 -11913 15148 -11887
rect 15148 -11913 15149 -11887
rect 15121 -11914 15149 -11913
rect 15121 -12047 15149 -12046
rect 15121 -12073 15122 -12047
rect 15122 -12073 15148 -12047
rect 15148 -12073 15149 -12047
rect 15121 -12074 15149 -12073
rect 15121 -12207 15149 -12206
rect 15121 -12233 15122 -12207
rect 15122 -12233 15148 -12207
rect 15148 -12233 15149 -12207
rect 15121 -12234 15149 -12233
rect 15121 -12367 15149 -12366
rect 15121 -12393 15122 -12367
rect 15122 -12393 15148 -12367
rect 15148 -12393 15149 -12367
rect 15121 -12394 15149 -12393
rect 15121 -12527 15149 -12526
rect 15121 -12553 15122 -12527
rect 15122 -12553 15148 -12527
rect 15148 -12553 15149 -12527
rect 15121 -12554 15149 -12553
rect 15121 -12687 15149 -12686
rect 15121 -12713 15122 -12687
rect 15122 -12713 15148 -12687
rect 15148 -12713 15149 -12687
rect 15121 -12714 15149 -12713
rect 15121 -12847 15149 -12846
rect 15121 -12873 15122 -12847
rect 15122 -12873 15148 -12847
rect 15148 -12873 15149 -12847
rect 15121 -12874 15149 -12873
rect 15121 -13007 15149 -13006
rect 15121 -13033 15122 -13007
rect 15122 -13033 15148 -13007
rect 15148 -13033 15149 -13007
rect 15121 -13034 15149 -13033
rect 15121 -13167 15149 -13166
rect 15121 -13193 15122 -13167
rect 15122 -13193 15148 -13167
rect 15148 -13193 15149 -13167
rect 15121 -13194 15149 -13193
rect 15121 -13327 15149 -13326
rect 15121 -13353 15122 -13327
rect 15122 -13353 15148 -13327
rect 15148 -13353 15149 -13327
rect 15121 -13354 15149 -13353
rect 15121 -13487 15149 -13486
rect 15121 -13513 15122 -13487
rect 15122 -13513 15148 -13487
rect 15148 -13513 15149 -13487
rect 15121 -13514 15149 -13513
rect 15121 -13647 15149 -13646
rect 15121 -13673 15122 -13647
rect 15122 -13673 15148 -13647
rect 15148 -13673 15149 -13647
rect 15121 -13674 15149 -13673
rect 15121 -13807 15149 -13806
rect 15121 -13833 15122 -13807
rect 15122 -13833 15148 -13807
rect 15148 -13833 15149 -13807
rect 15121 -13834 15149 -13833
rect 15121 -13967 15149 -13966
rect 15121 -13993 15122 -13967
rect 15122 -13993 15148 -13967
rect 15148 -13993 15149 -13967
rect 15121 -13994 15149 -13993
rect 15121 -14127 15149 -14126
rect 15121 -14153 15122 -14127
rect 15122 -14153 15148 -14127
rect 15148 -14153 15149 -14127
rect 15121 -14154 15149 -14153
rect 15121 -14287 15149 -14286
rect 15121 -14313 15122 -14287
rect 15122 -14313 15148 -14287
rect 15148 -14313 15149 -14287
rect 15121 -14314 15149 -14313
rect 15121 -14447 15149 -14446
rect 15121 -14473 15122 -14447
rect 15122 -14473 15148 -14447
rect 15148 -14473 15149 -14447
rect 15121 -14474 15149 -14473
rect 15121 -14607 15149 -14606
rect 15121 -14633 15122 -14607
rect 15122 -14633 15148 -14607
rect 15148 -14633 15149 -14607
rect 15121 -14634 15149 -14633
rect 15121 -14767 15149 -14766
rect 15121 -14793 15122 -14767
rect 15122 -14793 15148 -14767
rect 15148 -14793 15149 -14767
rect 15121 -14794 15149 -14793
rect 15121 -14927 15149 -14926
rect 15121 -14953 15122 -14927
rect 15122 -14953 15148 -14927
rect 15148 -14953 15149 -14927
rect 15121 -14954 15149 -14953
rect 15121 -15087 15149 -15086
rect 15121 -15113 15122 -15087
rect 15122 -15113 15148 -15087
rect 15148 -15113 15149 -15087
rect 15121 -15114 15149 -15113
rect 18854 -11887 18882 -11886
rect 18854 -11913 18855 -11887
rect 18855 -11913 18881 -11887
rect 18881 -11913 18882 -11887
rect 18854 -11914 18882 -11913
rect 18854 -12047 18882 -12046
rect 18854 -12073 18855 -12047
rect 18855 -12073 18881 -12047
rect 18881 -12073 18882 -12047
rect 18854 -12074 18882 -12073
rect 18854 -12207 18882 -12206
rect 18854 -12233 18855 -12207
rect 18855 -12233 18881 -12207
rect 18881 -12233 18882 -12207
rect 18854 -12234 18882 -12233
rect 18854 -12367 18882 -12366
rect 18854 -12393 18855 -12367
rect 18855 -12393 18881 -12367
rect 18881 -12393 18882 -12367
rect 18854 -12394 18882 -12393
rect 18854 -12527 18882 -12526
rect 18854 -12553 18855 -12527
rect 18855 -12553 18881 -12527
rect 18881 -12553 18882 -12527
rect 18854 -12554 18882 -12553
rect 18854 -12687 18882 -12686
rect 18854 -12713 18855 -12687
rect 18855 -12713 18881 -12687
rect 18881 -12713 18882 -12687
rect 18854 -12714 18882 -12713
rect 18854 -12847 18882 -12846
rect 18854 -12873 18855 -12847
rect 18855 -12873 18881 -12847
rect 18881 -12873 18882 -12847
rect 18854 -12874 18882 -12873
rect 18854 -13007 18882 -13006
rect 18854 -13033 18855 -13007
rect 18855 -13033 18881 -13007
rect 18881 -13033 18882 -13007
rect 18854 -13034 18882 -13033
rect 18854 -13167 18882 -13166
rect 18854 -13193 18855 -13167
rect 18855 -13193 18881 -13167
rect 18881 -13193 18882 -13167
rect 18854 -13194 18882 -13193
rect 18854 -13327 18882 -13326
rect 18854 -13353 18855 -13327
rect 18855 -13353 18881 -13327
rect 18881 -13353 18882 -13327
rect 18854 -13354 18882 -13353
rect 18854 -13487 18882 -13486
rect 18854 -13513 18855 -13487
rect 18855 -13513 18881 -13487
rect 18881 -13513 18882 -13487
rect 18854 -13514 18882 -13513
rect 18854 -13647 18882 -13646
rect 18854 -13673 18855 -13647
rect 18855 -13673 18881 -13647
rect 18881 -13673 18882 -13647
rect 18854 -13674 18882 -13673
rect 18854 -13807 18882 -13806
rect 18854 -13833 18855 -13807
rect 18855 -13833 18881 -13807
rect 18881 -13833 18882 -13807
rect 18854 -13834 18882 -13833
rect 18854 -13967 18882 -13966
rect 18854 -13993 18855 -13967
rect 18855 -13993 18881 -13967
rect 18881 -13993 18882 -13967
rect 18854 -13994 18882 -13993
rect 18854 -14127 18882 -14126
rect 18854 -14153 18855 -14127
rect 18855 -14153 18881 -14127
rect 18881 -14153 18882 -14127
rect 18854 -14154 18882 -14153
rect 18854 -14287 18882 -14286
rect 18854 -14313 18855 -14287
rect 18855 -14313 18881 -14287
rect 18881 -14313 18882 -14287
rect 18854 -14314 18882 -14313
rect 18854 -14447 18882 -14446
rect 18854 -14473 18855 -14447
rect 18855 -14473 18881 -14447
rect 18881 -14473 18882 -14447
rect 18854 -14474 18882 -14473
rect 18854 -14607 18882 -14606
rect 18854 -14633 18855 -14607
rect 18855 -14633 18881 -14607
rect 18881 -14633 18882 -14607
rect 18854 -14634 18882 -14633
rect 18854 -14767 18882 -14766
rect 18854 -14793 18855 -14767
rect 18855 -14793 18881 -14767
rect 18881 -14793 18882 -14767
rect 18854 -14794 18882 -14793
rect 18854 -14927 18882 -14926
rect 18854 -14953 18855 -14927
rect 18855 -14953 18881 -14927
rect 18881 -14953 18882 -14927
rect 18854 -14954 18882 -14953
rect 18854 -15087 18882 -15086
rect 18854 -15113 18855 -15087
rect 18855 -15113 18881 -15087
rect 18881 -15113 18882 -15087
rect 18854 -15114 18882 -15113
rect 15121 -15247 15149 -15246
rect 15121 -15273 15122 -15247
rect 15122 -15273 15148 -15247
rect 15148 -15273 15149 -15247
rect 15121 -15274 15149 -15273
rect 18854 -15247 18882 -15246
rect 18854 -15273 18855 -15247
rect 18855 -15273 18881 -15247
rect 18881 -15273 18882 -15247
rect 18854 -15274 18882 -15273
rect 15306 -15352 15334 -15351
rect 15306 -15378 15307 -15352
rect 15307 -15378 15333 -15352
rect 15333 -15378 15334 -15352
rect 15306 -15379 15334 -15378
rect 15466 -15352 15494 -15351
rect 15466 -15378 15467 -15352
rect 15467 -15378 15493 -15352
rect 15493 -15378 15494 -15352
rect 15466 -15379 15494 -15378
rect 15626 -15352 15654 -15351
rect 15626 -15378 15627 -15352
rect 15627 -15378 15653 -15352
rect 15653 -15378 15654 -15352
rect 15626 -15379 15654 -15378
rect 15786 -15352 15814 -15351
rect 15786 -15378 15787 -15352
rect 15787 -15378 15813 -15352
rect 15813 -15378 15814 -15352
rect 15786 -15379 15814 -15378
rect 15946 -15352 15974 -15351
rect 15946 -15378 15947 -15352
rect 15947 -15378 15973 -15352
rect 15973 -15378 15974 -15352
rect 15946 -15379 15974 -15378
rect 16106 -15352 16134 -15351
rect 16106 -15378 16107 -15352
rect 16107 -15378 16133 -15352
rect 16133 -15378 16134 -15352
rect 16106 -15379 16134 -15378
rect 16266 -15352 16294 -15351
rect 16266 -15378 16267 -15352
rect 16267 -15378 16293 -15352
rect 16293 -15378 16294 -15352
rect 16266 -15379 16294 -15378
rect 16426 -15352 16454 -15351
rect 16426 -15378 16427 -15352
rect 16427 -15378 16453 -15352
rect 16453 -15378 16454 -15352
rect 16426 -15379 16454 -15378
rect 16586 -15352 16614 -15351
rect 16586 -15378 16587 -15352
rect 16587 -15378 16613 -15352
rect 16613 -15378 16614 -15352
rect 16586 -15379 16614 -15378
rect 16746 -15352 16774 -15351
rect 16746 -15378 16747 -15352
rect 16747 -15378 16773 -15352
rect 16773 -15378 16774 -15352
rect 16746 -15379 16774 -15378
rect 16906 -15352 16934 -15351
rect 16906 -15378 16907 -15352
rect 16907 -15378 16933 -15352
rect 16933 -15378 16934 -15352
rect 16906 -15379 16934 -15378
rect 17066 -15352 17094 -15351
rect 17066 -15378 17067 -15352
rect 17067 -15378 17093 -15352
rect 17093 -15378 17094 -15352
rect 17066 -15379 17094 -15378
rect 17226 -15352 17254 -15351
rect 17226 -15378 17227 -15352
rect 17227 -15378 17253 -15352
rect 17253 -15378 17254 -15352
rect 17226 -15379 17254 -15378
rect 17386 -15352 17414 -15351
rect 17386 -15378 17387 -15352
rect 17387 -15378 17413 -15352
rect 17413 -15378 17414 -15352
rect 17386 -15379 17414 -15378
rect 17546 -15352 17574 -15351
rect 17546 -15378 17547 -15352
rect 17547 -15378 17573 -15352
rect 17573 -15378 17574 -15352
rect 17546 -15379 17574 -15378
rect 17706 -15352 17734 -15351
rect 17706 -15378 17707 -15352
rect 17707 -15378 17733 -15352
rect 17733 -15378 17734 -15352
rect 17706 -15379 17734 -15378
rect 17866 -15352 17894 -15351
rect 17866 -15378 17867 -15352
rect 17867 -15378 17893 -15352
rect 17893 -15378 17894 -15352
rect 17866 -15379 17894 -15378
rect 18026 -15352 18054 -15351
rect 18026 -15378 18027 -15352
rect 18027 -15378 18053 -15352
rect 18053 -15378 18054 -15352
rect 18026 -15379 18054 -15378
rect 18186 -15352 18214 -15351
rect 18186 -15378 18187 -15352
rect 18187 -15378 18213 -15352
rect 18213 -15378 18214 -15352
rect 18186 -15379 18214 -15378
rect 18346 -15352 18374 -15351
rect 18346 -15378 18347 -15352
rect 18347 -15378 18373 -15352
rect 18373 -15378 18374 -15352
rect 18346 -15379 18374 -15378
rect 18506 -15352 18534 -15351
rect 18506 -15378 18507 -15352
rect 18507 -15378 18533 -15352
rect 18533 -15378 18534 -15352
rect 18506 -15379 18534 -15378
rect 18666 -15352 18694 -15351
rect 18666 -15378 18667 -15352
rect 18667 -15378 18693 -15352
rect 18693 -15378 18694 -15352
rect 18666 -15379 18694 -15378
rect 21306 -11624 21334 -11623
rect 21306 -11650 21307 -11624
rect 21307 -11650 21333 -11624
rect 21333 -11650 21334 -11624
rect 21306 -11651 21334 -11650
rect 21466 -11624 21494 -11623
rect 21466 -11650 21467 -11624
rect 21467 -11650 21493 -11624
rect 21493 -11650 21494 -11624
rect 21466 -11651 21494 -11650
rect 21626 -11624 21654 -11623
rect 21626 -11650 21627 -11624
rect 21627 -11650 21653 -11624
rect 21653 -11650 21654 -11624
rect 21626 -11651 21654 -11650
rect 21786 -11624 21814 -11623
rect 21786 -11650 21787 -11624
rect 21787 -11650 21813 -11624
rect 21813 -11650 21814 -11624
rect 21786 -11651 21814 -11650
rect 21946 -11624 21974 -11623
rect 21946 -11650 21947 -11624
rect 21947 -11650 21973 -11624
rect 21973 -11650 21974 -11624
rect 21946 -11651 21974 -11650
rect 22106 -11624 22134 -11623
rect 22106 -11650 22107 -11624
rect 22107 -11650 22133 -11624
rect 22133 -11650 22134 -11624
rect 22106 -11651 22134 -11650
rect 22266 -11624 22294 -11623
rect 22266 -11650 22267 -11624
rect 22267 -11650 22293 -11624
rect 22293 -11650 22294 -11624
rect 22266 -11651 22294 -11650
rect 22426 -11624 22454 -11623
rect 22426 -11650 22427 -11624
rect 22427 -11650 22453 -11624
rect 22453 -11650 22454 -11624
rect 22426 -11651 22454 -11650
rect 22586 -11624 22614 -11623
rect 22586 -11650 22587 -11624
rect 22587 -11650 22613 -11624
rect 22613 -11650 22614 -11624
rect 22586 -11651 22614 -11650
rect 22746 -11624 22774 -11623
rect 22746 -11650 22747 -11624
rect 22747 -11650 22773 -11624
rect 22773 -11650 22774 -11624
rect 22746 -11651 22774 -11650
rect 22906 -11624 22934 -11623
rect 22906 -11650 22907 -11624
rect 22907 -11650 22933 -11624
rect 22933 -11650 22934 -11624
rect 22906 -11651 22934 -11650
rect 23066 -11624 23094 -11623
rect 23066 -11650 23067 -11624
rect 23067 -11650 23093 -11624
rect 23093 -11650 23094 -11624
rect 23066 -11651 23094 -11650
rect 23226 -11624 23254 -11623
rect 23226 -11650 23227 -11624
rect 23227 -11650 23253 -11624
rect 23253 -11650 23254 -11624
rect 23226 -11651 23254 -11650
rect 23386 -11624 23414 -11623
rect 23386 -11650 23387 -11624
rect 23387 -11650 23413 -11624
rect 23413 -11650 23414 -11624
rect 23386 -11651 23414 -11650
rect 23546 -11624 23574 -11623
rect 23546 -11650 23547 -11624
rect 23547 -11650 23573 -11624
rect 23573 -11650 23574 -11624
rect 23546 -11651 23574 -11650
rect 23706 -11624 23734 -11623
rect 23706 -11650 23707 -11624
rect 23707 -11650 23733 -11624
rect 23733 -11650 23734 -11624
rect 23706 -11651 23734 -11650
rect 23866 -11624 23894 -11623
rect 23866 -11650 23867 -11624
rect 23867 -11650 23893 -11624
rect 23893 -11650 23894 -11624
rect 23866 -11651 23894 -11650
rect 24026 -11624 24054 -11623
rect 24026 -11650 24027 -11624
rect 24027 -11650 24053 -11624
rect 24053 -11650 24054 -11624
rect 24026 -11651 24054 -11650
rect 24186 -11624 24214 -11623
rect 24186 -11650 24187 -11624
rect 24187 -11650 24213 -11624
rect 24213 -11650 24214 -11624
rect 24186 -11651 24214 -11650
rect 24346 -11624 24374 -11623
rect 24346 -11650 24347 -11624
rect 24347 -11650 24373 -11624
rect 24373 -11650 24374 -11624
rect 24346 -11651 24374 -11650
rect 24506 -11624 24534 -11623
rect 24506 -11650 24507 -11624
rect 24507 -11650 24533 -11624
rect 24533 -11650 24534 -11624
rect 24506 -11651 24534 -11650
rect 24666 -11624 24694 -11623
rect 24666 -11650 24667 -11624
rect 24667 -11650 24693 -11624
rect 24693 -11650 24694 -11624
rect 24666 -11651 24694 -11650
rect 21121 -11727 21149 -11726
rect 21121 -11753 21122 -11727
rect 21122 -11753 21148 -11727
rect 21148 -11753 21149 -11727
rect 21121 -11754 21149 -11753
rect 24854 -11727 24882 -11726
rect 24854 -11753 24855 -11727
rect 24855 -11753 24881 -11727
rect 24881 -11753 24882 -11727
rect 24854 -11754 24882 -11753
rect 21121 -11887 21149 -11886
rect 21121 -11913 21122 -11887
rect 21122 -11913 21148 -11887
rect 21148 -11913 21149 -11887
rect 21121 -11914 21149 -11913
rect 21121 -12047 21149 -12046
rect 21121 -12073 21122 -12047
rect 21122 -12073 21148 -12047
rect 21148 -12073 21149 -12047
rect 21121 -12074 21149 -12073
rect 21121 -12207 21149 -12206
rect 21121 -12233 21122 -12207
rect 21122 -12233 21148 -12207
rect 21148 -12233 21149 -12207
rect 21121 -12234 21149 -12233
rect 21121 -12367 21149 -12366
rect 21121 -12393 21122 -12367
rect 21122 -12393 21148 -12367
rect 21148 -12393 21149 -12367
rect 21121 -12394 21149 -12393
rect 21121 -12527 21149 -12526
rect 21121 -12553 21122 -12527
rect 21122 -12553 21148 -12527
rect 21148 -12553 21149 -12527
rect 21121 -12554 21149 -12553
rect 21121 -12687 21149 -12686
rect 21121 -12713 21122 -12687
rect 21122 -12713 21148 -12687
rect 21148 -12713 21149 -12687
rect 21121 -12714 21149 -12713
rect 21121 -12847 21149 -12846
rect 21121 -12873 21122 -12847
rect 21122 -12873 21148 -12847
rect 21148 -12873 21149 -12847
rect 21121 -12874 21149 -12873
rect 21121 -13007 21149 -13006
rect 21121 -13033 21122 -13007
rect 21122 -13033 21148 -13007
rect 21148 -13033 21149 -13007
rect 21121 -13034 21149 -13033
rect 21121 -13167 21149 -13166
rect 21121 -13193 21122 -13167
rect 21122 -13193 21148 -13167
rect 21148 -13193 21149 -13167
rect 21121 -13194 21149 -13193
rect 21121 -13327 21149 -13326
rect 21121 -13353 21122 -13327
rect 21122 -13353 21148 -13327
rect 21148 -13353 21149 -13327
rect 21121 -13354 21149 -13353
rect 21121 -13487 21149 -13486
rect 21121 -13513 21122 -13487
rect 21122 -13513 21148 -13487
rect 21148 -13513 21149 -13487
rect 21121 -13514 21149 -13513
rect 21121 -13647 21149 -13646
rect 21121 -13673 21122 -13647
rect 21122 -13673 21148 -13647
rect 21148 -13673 21149 -13647
rect 21121 -13674 21149 -13673
rect 21121 -13807 21149 -13806
rect 21121 -13833 21122 -13807
rect 21122 -13833 21148 -13807
rect 21148 -13833 21149 -13807
rect 21121 -13834 21149 -13833
rect 21121 -13967 21149 -13966
rect 21121 -13993 21122 -13967
rect 21122 -13993 21148 -13967
rect 21148 -13993 21149 -13967
rect 21121 -13994 21149 -13993
rect 21121 -14127 21149 -14126
rect 21121 -14153 21122 -14127
rect 21122 -14153 21148 -14127
rect 21148 -14153 21149 -14127
rect 21121 -14154 21149 -14153
rect 21121 -14287 21149 -14286
rect 21121 -14313 21122 -14287
rect 21122 -14313 21148 -14287
rect 21148 -14313 21149 -14287
rect 21121 -14314 21149 -14313
rect 21121 -14447 21149 -14446
rect 21121 -14473 21122 -14447
rect 21122 -14473 21148 -14447
rect 21148 -14473 21149 -14447
rect 21121 -14474 21149 -14473
rect 21121 -14607 21149 -14606
rect 21121 -14633 21122 -14607
rect 21122 -14633 21148 -14607
rect 21148 -14633 21149 -14607
rect 21121 -14634 21149 -14633
rect 21121 -14767 21149 -14766
rect 21121 -14793 21122 -14767
rect 21122 -14793 21148 -14767
rect 21148 -14793 21149 -14767
rect 21121 -14794 21149 -14793
rect 21121 -14927 21149 -14926
rect 21121 -14953 21122 -14927
rect 21122 -14953 21148 -14927
rect 21148 -14953 21149 -14927
rect 21121 -14954 21149 -14953
rect 21121 -15087 21149 -15086
rect 21121 -15113 21122 -15087
rect 21122 -15113 21148 -15087
rect 21148 -15113 21149 -15087
rect 21121 -15114 21149 -15113
rect 24854 -11887 24882 -11886
rect 24854 -11913 24855 -11887
rect 24855 -11913 24881 -11887
rect 24881 -11913 24882 -11887
rect 24854 -11914 24882 -11913
rect 24854 -12047 24882 -12046
rect 24854 -12073 24855 -12047
rect 24855 -12073 24881 -12047
rect 24881 -12073 24882 -12047
rect 24854 -12074 24882 -12073
rect 24854 -12207 24882 -12206
rect 24854 -12233 24855 -12207
rect 24855 -12233 24881 -12207
rect 24881 -12233 24882 -12207
rect 24854 -12234 24882 -12233
rect 24854 -12367 24882 -12366
rect 24854 -12393 24855 -12367
rect 24855 -12393 24881 -12367
rect 24881 -12393 24882 -12367
rect 24854 -12394 24882 -12393
rect 24854 -12527 24882 -12526
rect 24854 -12553 24855 -12527
rect 24855 -12553 24881 -12527
rect 24881 -12553 24882 -12527
rect 24854 -12554 24882 -12553
rect 24854 -12687 24882 -12686
rect 24854 -12713 24855 -12687
rect 24855 -12713 24881 -12687
rect 24881 -12713 24882 -12687
rect 24854 -12714 24882 -12713
rect 24854 -12847 24882 -12846
rect 24854 -12873 24855 -12847
rect 24855 -12873 24881 -12847
rect 24881 -12873 24882 -12847
rect 24854 -12874 24882 -12873
rect 24854 -13007 24882 -13006
rect 24854 -13033 24855 -13007
rect 24855 -13033 24881 -13007
rect 24881 -13033 24882 -13007
rect 24854 -13034 24882 -13033
rect 24854 -13167 24882 -13166
rect 24854 -13193 24855 -13167
rect 24855 -13193 24881 -13167
rect 24881 -13193 24882 -13167
rect 24854 -13194 24882 -13193
rect 24854 -13327 24882 -13326
rect 24854 -13353 24855 -13327
rect 24855 -13353 24881 -13327
rect 24881 -13353 24882 -13327
rect 24854 -13354 24882 -13353
rect 24854 -13487 24882 -13486
rect 24854 -13513 24855 -13487
rect 24855 -13513 24881 -13487
rect 24881 -13513 24882 -13487
rect 24854 -13514 24882 -13513
rect 24854 -13647 24882 -13646
rect 24854 -13673 24855 -13647
rect 24855 -13673 24881 -13647
rect 24881 -13673 24882 -13647
rect 24854 -13674 24882 -13673
rect 24854 -13807 24882 -13806
rect 24854 -13833 24855 -13807
rect 24855 -13833 24881 -13807
rect 24881 -13833 24882 -13807
rect 24854 -13834 24882 -13833
rect 24854 -13967 24882 -13966
rect 24854 -13993 24855 -13967
rect 24855 -13993 24881 -13967
rect 24881 -13993 24882 -13967
rect 24854 -13994 24882 -13993
rect 24854 -14127 24882 -14126
rect 24854 -14153 24855 -14127
rect 24855 -14153 24881 -14127
rect 24881 -14153 24882 -14127
rect 24854 -14154 24882 -14153
rect 24854 -14287 24882 -14286
rect 24854 -14313 24855 -14287
rect 24855 -14313 24881 -14287
rect 24881 -14313 24882 -14287
rect 24854 -14314 24882 -14313
rect 24854 -14447 24882 -14446
rect 24854 -14473 24855 -14447
rect 24855 -14473 24881 -14447
rect 24881 -14473 24882 -14447
rect 24854 -14474 24882 -14473
rect 24854 -14607 24882 -14606
rect 24854 -14633 24855 -14607
rect 24855 -14633 24881 -14607
rect 24881 -14633 24882 -14607
rect 24854 -14634 24882 -14633
rect 24854 -14767 24882 -14766
rect 24854 -14793 24855 -14767
rect 24855 -14793 24881 -14767
rect 24881 -14793 24882 -14767
rect 24854 -14794 24882 -14793
rect 24854 -14927 24882 -14926
rect 24854 -14953 24855 -14927
rect 24855 -14953 24881 -14927
rect 24881 -14953 24882 -14927
rect 24854 -14954 24882 -14953
rect 24854 -15087 24882 -15086
rect 24854 -15113 24855 -15087
rect 24855 -15113 24881 -15087
rect 24881 -15113 24882 -15087
rect 24854 -15114 24882 -15113
rect 21121 -15247 21149 -15246
rect 21121 -15273 21122 -15247
rect 21122 -15273 21148 -15247
rect 21148 -15273 21149 -15247
rect 21121 -15274 21149 -15273
rect 24854 -15247 24882 -15246
rect 24854 -15273 24855 -15247
rect 24855 -15273 24881 -15247
rect 24881 -15273 24882 -15247
rect 24854 -15274 24882 -15273
rect 21306 -15352 21334 -15351
rect 21306 -15378 21307 -15352
rect 21307 -15378 21333 -15352
rect 21333 -15378 21334 -15352
rect 21306 -15379 21334 -15378
rect 21466 -15352 21494 -15351
rect 21466 -15378 21467 -15352
rect 21467 -15378 21493 -15352
rect 21493 -15378 21494 -15352
rect 21466 -15379 21494 -15378
rect 21626 -15352 21654 -15351
rect 21626 -15378 21627 -15352
rect 21627 -15378 21653 -15352
rect 21653 -15378 21654 -15352
rect 21626 -15379 21654 -15378
rect 21786 -15352 21814 -15351
rect 21786 -15378 21787 -15352
rect 21787 -15378 21813 -15352
rect 21813 -15378 21814 -15352
rect 21786 -15379 21814 -15378
rect 21946 -15352 21974 -15351
rect 21946 -15378 21947 -15352
rect 21947 -15378 21973 -15352
rect 21973 -15378 21974 -15352
rect 21946 -15379 21974 -15378
rect 22106 -15352 22134 -15351
rect 22106 -15378 22107 -15352
rect 22107 -15378 22133 -15352
rect 22133 -15378 22134 -15352
rect 22106 -15379 22134 -15378
rect 22266 -15352 22294 -15351
rect 22266 -15378 22267 -15352
rect 22267 -15378 22293 -15352
rect 22293 -15378 22294 -15352
rect 22266 -15379 22294 -15378
rect 22426 -15352 22454 -15351
rect 22426 -15378 22427 -15352
rect 22427 -15378 22453 -15352
rect 22453 -15378 22454 -15352
rect 22426 -15379 22454 -15378
rect 22586 -15352 22614 -15351
rect 22586 -15378 22587 -15352
rect 22587 -15378 22613 -15352
rect 22613 -15378 22614 -15352
rect 22586 -15379 22614 -15378
rect 22746 -15352 22774 -15351
rect 22746 -15378 22747 -15352
rect 22747 -15378 22773 -15352
rect 22773 -15378 22774 -15352
rect 22746 -15379 22774 -15378
rect 22906 -15352 22934 -15351
rect 22906 -15378 22907 -15352
rect 22907 -15378 22933 -15352
rect 22933 -15378 22934 -15352
rect 22906 -15379 22934 -15378
rect 23066 -15352 23094 -15351
rect 23066 -15378 23067 -15352
rect 23067 -15378 23093 -15352
rect 23093 -15378 23094 -15352
rect 23066 -15379 23094 -15378
rect 23226 -15352 23254 -15351
rect 23226 -15378 23227 -15352
rect 23227 -15378 23253 -15352
rect 23253 -15378 23254 -15352
rect 23226 -15379 23254 -15378
rect 23386 -15352 23414 -15351
rect 23386 -15378 23387 -15352
rect 23387 -15378 23413 -15352
rect 23413 -15378 23414 -15352
rect 23386 -15379 23414 -15378
rect 23546 -15352 23574 -15351
rect 23546 -15378 23547 -15352
rect 23547 -15378 23573 -15352
rect 23573 -15378 23574 -15352
rect 23546 -15379 23574 -15378
rect 23706 -15352 23734 -15351
rect 23706 -15378 23707 -15352
rect 23707 -15378 23733 -15352
rect 23733 -15378 23734 -15352
rect 23706 -15379 23734 -15378
rect 23866 -15352 23894 -15351
rect 23866 -15378 23867 -15352
rect 23867 -15378 23893 -15352
rect 23893 -15378 23894 -15352
rect 23866 -15379 23894 -15378
rect 24026 -15352 24054 -15351
rect 24026 -15378 24027 -15352
rect 24027 -15378 24053 -15352
rect 24053 -15378 24054 -15352
rect 24026 -15379 24054 -15378
rect 24186 -15352 24214 -15351
rect 24186 -15378 24187 -15352
rect 24187 -15378 24213 -15352
rect 24213 -15378 24214 -15352
rect 24186 -15379 24214 -15378
rect 24346 -15352 24374 -15351
rect 24346 -15378 24347 -15352
rect 24347 -15378 24373 -15352
rect 24373 -15378 24374 -15352
rect 24346 -15379 24374 -15378
rect 24506 -15352 24534 -15351
rect 24506 -15378 24507 -15352
rect 24507 -15378 24533 -15352
rect 24533 -15378 24534 -15352
rect 24506 -15379 24534 -15378
rect 24666 -15352 24694 -15351
rect 24666 -15378 24667 -15352
rect 24667 -15378 24693 -15352
rect 24693 -15378 24694 -15352
rect 24666 -15379 24694 -15378
<< metal3 >>
rect 3000 9381 7000 9500
rect 3000 9349 3304 9381
rect 3336 9349 3464 9381
rect 3496 9349 3624 9381
rect 3656 9349 3784 9381
rect 3816 9349 3944 9381
rect 3976 9349 4104 9381
rect 4136 9349 4264 9381
rect 4296 9349 4424 9381
rect 4456 9349 4584 9381
rect 4616 9349 4744 9381
rect 4776 9349 4904 9381
rect 4936 9349 5064 9381
rect 5096 9349 5224 9381
rect 5256 9349 5384 9381
rect 5416 9349 5544 9381
rect 5576 9349 5704 9381
rect 5736 9349 5864 9381
rect 5896 9349 6024 9381
rect 6056 9349 6184 9381
rect 6216 9349 6344 9381
rect 6376 9349 6504 9381
rect 6536 9349 6664 9381
rect 6696 9349 7000 9381
rect 3000 9276 7000 9349
rect 3000 9244 3116 9276
rect 3148 9244 6849 9276
rect 6881 9244 7000 9276
rect 3000 9230 7000 9244
rect 3000 9116 3270 9230
rect 3000 9084 3116 9116
rect 3148 9084 3270 9116
rect 3000 8956 3270 9084
rect 3000 8924 3116 8956
rect 3148 8924 3270 8956
rect 3000 8796 3270 8924
rect 3000 8764 3116 8796
rect 3148 8764 3270 8796
rect 3000 8636 3270 8764
rect 3000 8604 3116 8636
rect 3148 8604 3270 8636
rect 3000 8476 3270 8604
rect 3000 8444 3116 8476
rect 3148 8444 3270 8476
rect 3000 8316 3270 8444
rect 3000 8284 3116 8316
rect 3148 8284 3270 8316
rect 3000 8156 3270 8284
rect 3000 8124 3116 8156
rect 3148 8124 3270 8156
rect 3000 7996 3270 8124
rect 3000 7964 3116 7996
rect 3148 7964 3270 7996
rect 3000 7836 3270 7964
rect 3000 7804 3116 7836
rect 3148 7804 3270 7836
rect 3000 7676 3270 7804
rect 3000 7644 3116 7676
rect 3148 7644 3270 7676
rect 3000 7516 3270 7644
rect 3000 7484 3116 7516
rect 3148 7484 3270 7516
rect 3000 7356 3270 7484
rect 3000 7324 3116 7356
rect 3148 7324 3270 7356
rect 3000 7196 3270 7324
rect 3000 7164 3116 7196
rect 3148 7164 3270 7196
rect 3000 7036 3270 7164
rect 3000 7004 3116 7036
rect 3148 7004 3270 7036
rect 3000 6876 3270 7004
rect 3000 6844 3116 6876
rect 3148 6844 3270 6876
rect 3000 6716 3270 6844
rect 3000 6684 3116 6716
rect 3148 6684 3270 6716
rect 3000 6556 3270 6684
rect 3000 6524 3116 6556
rect 3148 6524 3270 6556
rect 3000 6396 3270 6524
rect 3000 6364 3116 6396
rect 3148 6364 3270 6396
rect 3000 6236 3270 6364
rect 3000 6204 3116 6236
rect 3148 6204 3270 6236
rect 3000 6076 3270 6204
rect 3000 6044 3116 6076
rect 3148 6044 3270 6076
rect 3000 5916 3270 6044
rect 3000 5884 3116 5916
rect 3148 5884 3270 5916
rect 3000 5770 3270 5884
rect 6730 9116 7000 9230
rect 6730 9084 6849 9116
rect 6881 9084 7000 9116
rect 6730 8956 7000 9084
rect 6730 8924 6849 8956
rect 6881 8924 7000 8956
rect 6730 8796 7000 8924
rect 6730 8764 6849 8796
rect 6881 8764 7000 8796
rect 6730 8636 7000 8764
rect 6730 8604 6849 8636
rect 6881 8604 7000 8636
rect 6730 8476 7000 8604
rect 6730 8444 6849 8476
rect 6881 8444 7000 8476
rect 6730 8316 7000 8444
rect 6730 8284 6849 8316
rect 6881 8284 7000 8316
rect 6730 8156 7000 8284
rect 6730 8124 6849 8156
rect 6881 8124 7000 8156
rect 6730 7996 7000 8124
rect 6730 7964 6849 7996
rect 6881 7964 7000 7996
rect 6730 7836 7000 7964
rect 6730 7804 6849 7836
rect 6881 7804 7000 7836
rect 6730 7676 7000 7804
rect 6730 7644 6849 7676
rect 6881 7644 7000 7676
rect 6730 7516 7000 7644
rect 6730 7484 6849 7516
rect 6881 7484 7000 7516
rect 6730 7356 7000 7484
rect 6730 7324 6849 7356
rect 6881 7324 7000 7356
rect 6730 7196 7000 7324
rect 6730 7164 6849 7196
rect 6881 7164 7000 7196
rect 6730 7036 7000 7164
rect 6730 7004 6849 7036
rect 6881 7004 7000 7036
rect 6730 6876 7000 7004
rect 6730 6844 6849 6876
rect 6881 6844 7000 6876
rect 6730 6716 7000 6844
rect 6730 6684 6849 6716
rect 6881 6684 7000 6716
rect 6730 6556 7000 6684
rect 6730 6524 6849 6556
rect 6881 6524 7000 6556
rect 6730 6396 7000 6524
rect 6730 6364 6849 6396
rect 6881 6364 7000 6396
rect 6730 6236 7000 6364
rect 6730 6204 6849 6236
rect 6881 6204 7000 6236
rect 6730 6076 7000 6204
rect 6730 6044 6849 6076
rect 6881 6044 7000 6076
rect 6730 5916 7000 6044
rect 6730 5884 6849 5916
rect 6881 5884 7000 5916
rect 6730 5770 7000 5884
rect 3000 5756 7000 5770
rect 3000 5724 3116 5756
rect 3148 5724 6849 5756
rect 6881 5724 7000 5756
rect 3000 5653 7000 5724
rect 3000 5621 3304 5653
rect 3336 5621 3464 5653
rect 3496 5621 3624 5653
rect 3656 5621 3784 5653
rect 3816 5621 3944 5653
rect 3976 5621 4104 5653
rect 4136 5621 4264 5653
rect 4296 5621 4424 5653
rect 4456 5621 4584 5653
rect 4616 5621 4744 5653
rect 4776 5621 4904 5653
rect 4936 5621 5064 5653
rect 5096 5621 5224 5653
rect 5256 5621 5384 5653
rect 5416 5621 5544 5653
rect 5576 5621 5704 5653
rect 5736 5621 5864 5653
rect 5896 5621 6024 5653
rect 6056 5621 6184 5653
rect 6216 5621 6344 5653
rect 6376 5621 6504 5653
rect 6536 5621 6664 5653
rect 6696 5621 7000 5653
rect 3000 5500 7000 5621
rect 9000 9381 13000 9500
rect 9000 9349 9304 9381
rect 9336 9349 9464 9381
rect 9496 9349 9624 9381
rect 9656 9349 9784 9381
rect 9816 9349 9944 9381
rect 9976 9349 10104 9381
rect 10136 9349 10264 9381
rect 10296 9349 10424 9381
rect 10456 9349 10584 9381
rect 10616 9349 10744 9381
rect 10776 9349 10904 9381
rect 10936 9349 11064 9381
rect 11096 9349 11224 9381
rect 11256 9349 11384 9381
rect 11416 9349 11544 9381
rect 11576 9349 11704 9381
rect 11736 9349 11864 9381
rect 11896 9349 12024 9381
rect 12056 9349 12184 9381
rect 12216 9349 12344 9381
rect 12376 9349 12504 9381
rect 12536 9349 12664 9381
rect 12696 9349 13000 9381
rect 9000 9276 13000 9349
rect 9000 9244 9116 9276
rect 9148 9244 12849 9276
rect 12881 9244 13000 9276
rect 9000 9230 13000 9244
rect 9000 9116 9270 9230
rect 9000 9084 9116 9116
rect 9148 9084 9270 9116
rect 9000 8956 9270 9084
rect 9000 8924 9116 8956
rect 9148 8924 9270 8956
rect 9000 8796 9270 8924
rect 9000 8764 9116 8796
rect 9148 8764 9270 8796
rect 9000 8636 9270 8764
rect 9000 8604 9116 8636
rect 9148 8604 9270 8636
rect 9000 8476 9270 8604
rect 9000 8444 9116 8476
rect 9148 8444 9270 8476
rect 9000 8316 9270 8444
rect 9000 8284 9116 8316
rect 9148 8284 9270 8316
rect 9000 8156 9270 8284
rect 9000 8124 9116 8156
rect 9148 8124 9270 8156
rect 9000 7996 9270 8124
rect 9000 7964 9116 7996
rect 9148 7964 9270 7996
rect 9000 7836 9270 7964
rect 9000 7804 9116 7836
rect 9148 7804 9270 7836
rect 9000 7676 9270 7804
rect 9000 7644 9116 7676
rect 9148 7644 9270 7676
rect 9000 7516 9270 7644
rect 9000 7484 9116 7516
rect 9148 7484 9270 7516
rect 9000 7356 9270 7484
rect 9000 7324 9116 7356
rect 9148 7324 9270 7356
rect 9000 7196 9270 7324
rect 9000 7164 9116 7196
rect 9148 7164 9270 7196
rect 9000 7036 9270 7164
rect 9000 7004 9116 7036
rect 9148 7004 9270 7036
rect 9000 6876 9270 7004
rect 9000 6844 9116 6876
rect 9148 6844 9270 6876
rect 9000 6716 9270 6844
rect 9000 6684 9116 6716
rect 9148 6684 9270 6716
rect 9000 6556 9270 6684
rect 9000 6524 9116 6556
rect 9148 6524 9270 6556
rect 9000 6396 9270 6524
rect 9000 6364 9116 6396
rect 9148 6364 9270 6396
rect 9000 6236 9270 6364
rect 9000 6204 9116 6236
rect 9148 6204 9270 6236
rect 9000 6076 9270 6204
rect 9000 6044 9116 6076
rect 9148 6044 9270 6076
rect 9000 5916 9270 6044
rect 9000 5884 9116 5916
rect 9148 5884 9270 5916
rect 9000 5770 9270 5884
rect 12730 9116 13000 9230
rect 12730 9084 12849 9116
rect 12881 9084 13000 9116
rect 12730 8956 13000 9084
rect 12730 8924 12849 8956
rect 12881 8924 13000 8956
rect 12730 8796 13000 8924
rect 12730 8764 12849 8796
rect 12881 8764 13000 8796
rect 12730 8636 13000 8764
rect 12730 8604 12849 8636
rect 12881 8604 13000 8636
rect 12730 8476 13000 8604
rect 12730 8444 12849 8476
rect 12881 8444 13000 8476
rect 12730 8316 13000 8444
rect 12730 8284 12849 8316
rect 12881 8284 13000 8316
rect 12730 8156 13000 8284
rect 12730 8124 12849 8156
rect 12881 8124 13000 8156
rect 12730 7996 13000 8124
rect 12730 7964 12849 7996
rect 12881 7964 13000 7996
rect 12730 7836 13000 7964
rect 12730 7804 12849 7836
rect 12881 7804 13000 7836
rect 12730 7676 13000 7804
rect 12730 7644 12849 7676
rect 12881 7644 13000 7676
rect 12730 7516 13000 7644
rect 12730 7484 12849 7516
rect 12881 7484 13000 7516
rect 12730 7356 13000 7484
rect 12730 7324 12849 7356
rect 12881 7324 13000 7356
rect 12730 7196 13000 7324
rect 12730 7164 12849 7196
rect 12881 7164 13000 7196
rect 12730 7036 13000 7164
rect 12730 7004 12849 7036
rect 12881 7004 13000 7036
rect 12730 6900 13000 7004
rect 15000 9381 19000 9500
rect 15000 9349 15304 9381
rect 15336 9349 15464 9381
rect 15496 9349 15624 9381
rect 15656 9349 15784 9381
rect 15816 9349 15944 9381
rect 15976 9349 16104 9381
rect 16136 9349 16264 9381
rect 16296 9349 16424 9381
rect 16456 9349 16584 9381
rect 16616 9349 16744 9381
rect 16776 9349 16904 9381
rect 16936 9349 17064 9381
rect 17096 9349 17224 9381
rect 17256 9349 17384 9381
rect 17416 9349 17544 9381
rect 17576 9349 17704 9381
rect 17736 9349 17864 9381
rect 17896 9349 18024 9381
rect 18056 9349 18184 9381
rect 18216 9349 18344 9381
rect 18376 9349 18504 9381
rect 18536 9349 18664 9381
rect 18696 9349 19000 9381
rect 15000 9276 19000 9349
rect 15000 9244 15116 9276
rect 15148 9244 18849 9276
rect 18881 9244 19000 9276
rect 15000 9230 19000 9244
rect 15000 9116 15270 9230
rect 15000 9084 15116 9116
rect 15148 9084 15270 9116
rect 15000 8956 15270 9084
rect 15000 8924 15116 8956
rect 15148 8924 15270 8956
rect 15000 8796 15270 8924
rect 15000 8764 15116 8796
rect 15148 8764 15270 8796
rect 15000 8636 15270 8764
rect 15000 8604 15116 8636
rect 15148 8604 15270 8636
rect 15000 8476 15270 8604
rect 15000 8444 15116 8476
rect 15148 8444 15270 8476
rect 15000 8316 15270 8444
rect 15000 8284 15116 8316
rect 15148 8284 15270 8316
rect 15000 8156 15270 8284
rect 15000 8124 15116 8156
rect 15148 8124 15270 8156
rect 15000 7996 15270 8124
rect 15000 7964 15116 7996
rect 15148 7964 15270 7996
rect 15000 7836 15270 7964
rect 15000 7804 15116 7836
rect 15148 7804 15270 7836
rect 15000 7676 15270 7804
rect 15000 7644 15116 7676
rect 15148 7644 15270 7676
rect 15000 7516 15270 7644
rect 15000 7484 15116 7516
rect 15148 7484 15270 7516
rect 15000 7356 15270 7484
rect 15000 7324 15116 7356
rect 15148 7324 15270 7356
rect 15000 7196 15270 7324
rect 15000 7164 15116 7196
rect 15148 7164 15270 7196
rect 15000 7036 15270 7164
rect 15000 7004 15116 7036
rect 15148 7004 15270 7036
rect 12730 6876 13880 6900
rect 12730 6844 12849 6876
rect 12881 6870 13880 6876
rect 12881 6844 13000 6870
rect 12730 6716 13000 6844
rect 12730 6684 12849 6716
rect 12881 6684 13000 6716
rect 12730 6556 13000 6684
rect 12730 6524 12849 6556
rect 12881 6524 13000 6556
rect 12730 6396 13000 6524
rect 12730 6364 12849 6396
rect 12881 6364 13000 6396
rect 12730 6236 13000 6364
rect 12730 6204 12849 6236
rect 12881 6204 13000 6236
rect 12730 6076 13000 6204
rect 12730 6044 12849 6076
rect 12881 6044 13000 6076
rect 12730 5916 13000 6044
rect 12730 5884 12849 5916
rect 12881 5884 13000 5916
rect 12730 5770 13000 5884
rect 9000 5756 13000 5770
rect 9000 5724 9116 5756
rect 9148 5724 12849 5756
rect 12881 5724 13000 5756
rect 9000 5653 13000 5724
rect 9000 5621 9304 5653
rect 9336 5621 9464 5653
rect 9496 5621 9624 5653
rect 9656 5621 9784 5653
rect 9816 5621 9944 5653
rect 9976 5621 10104 5653
rect 10136 5621 10264 5653
rect 10296 5621 10424 5653
rect 10456 5621 10584 5653
rect 10616 5621 10744 5653
rect 10776 5621 10904 5653
rect 10936 5621 11064 5653
rect 11096 5621 11224 5653
rect 11256 5621 11384 5653
rect 11416 5621 11544 5653
rect 11576 5621 11704 5653
rect 11736 5621 11864 5653
rect 11896 5621 12024 5653
rect 12056 5621 12184 5653
rect 12216 5621 12344 5653
rect 12376 5621 12504 5653
rect 12536 5621 12664 5653
rect 12696 5621 13000 5653
rect 9000 5500 13000 5621
rect 6625 5160 6665 5500
rect 13850 5360 13880 6870
rect 15000 6876 15270 7004
rect 15000 6844 15116 6876
rect 15148 6844 15270 6876
rect 15000 6716 15270 6844
rect 15000 6684 15116 6716
rect 15148 6684 15270 6716
rect 15000 6556 15270 6684
rect 15000 6524 15116 6556
rect 15148 6524 15270 6556
rect 15000 6396 15270 6524
rect 15000 6364 15116 6396
rect 15148 6364 15270 6396
rect 15000 6236 15270 6364
rect 15000 6204 15116 6236
rect 15148 6204 15270 6236
rect 15000 6076 15270 6204
rect 15000 6044 15116 6076
rect 15148 6044 15270 6076
rect 15000 5916 15270 6044
rect 15000 5884 15116 5916
rect 15148 5884 15270 5916
rect 15000 5770 15270 5884
rect 18730 9116 19000 9230
rect 18730 9084 18849 9116
rect 18881 9084 19000 9116
rect 18730 8956 19000 9084
rect 18730 8924 18849 8956
rect 18881 8924 19000 8956
rect 18730 8796 19000 8924
rect 18730 8764 18849 8796
rect 18881 8764 19000 8796
rect 18730 8636 19000 8764
rect 18730 8604 18849 8636
rect 18881 8604 19000 8636
rect 18730 8476 19000 8604
rect 18730 8444 18849 8476
rect 18881 8444 19000 8476
rect 18730 8316 19000 8444
rect 18730 8284 18849 8316
rect 18881 8284 19000 8316
rect 18730 8156 19000 8284
rect 18730 8124 18849 8156
rect 18881 8124 19000 8156
rect 18730 7996 19000 8124
rect 18730 7964 18849 7996
rect 18881 7964 19000 7996
rect 18730 7836 19000 7964
rect 18730 7804 18849 7836
rect 18881 7804 19000 7836
rect 18730 7676 19000 7804
rect 18730 7644 18849 7676
rect 18881 7644 19000 7676
rect 18730 7516 19000 7644
rect 18730 7484 18849 7516
rect 18881 7484 19000 7516
rect 18730 7356 19000 7484
rect 18730 7324 18849 7356
rect 18881 7324 19000 7356
rect 18730 7196 19000 7324
rect 18730 7164 18849 7196
rect 18881 7164 19000 7196
rect 18730 7036 19000 7164
rect 18730 7004 18849 7036
rect 18881 7004 19000 7036
rect 18730 6905 19000 7004
rect 21000 9381 25000 9500
rect 21000 9349 21304 9381
rect 21336 9349 21464 9381
rect 21496 9349 21624 9381
rect 21656 9349 21784 9381
rect 21816 9349 21944 9381
rect 21976 9349 22104 9381
rect 22136 9349 22264 9381
rect 22296 9349 22424 9381
rect 22456 9349 22584 9381
rect 22616 9349 22744 9381
rect 22776 9349 22904 9381
rect 22936 9349 23064 9381
rect 23096 9349 23224 9381
rect 23256 9349 23384 9381
rect 23416 9349 23544 9381
rect 23576 9349 23704 9381
rect 23736 9349 23864 9381
rect 23896 9349 24024 9381
rect 24056 9349 24184 9381
rect 24216 9349 24344 9381
rect 24376 9349 24504 9381
rect 24536 9349 24664 9381
rect 24696 9349 25000 9381
rect 21000 9276 25000 9349
rect 21000 9244 21116 9276
rect 21148 9244 24849 9276
rect 24881 9244 25000 9276
rect 21000 9230 25000 9244
rect 21000 9116 21270 9230
rect 21000 9084 21116 9116
rect 21148 9084 21270 9116
rect 21000 8956 21270 9084
rect 21000 8924 21116 8956
rect 21148 8924 21270 8956
rect 21000 8796 21270 8924
rect 21000 8764 21116 8796
rect 21148 8764 21270 8796
rect 21000 8636 21270 8764
rect 21000 8604 21116 8636
rect 21148 8604 21270 8636
rect 21000 8476 21270 8604
rect 21000 8444 21116 8476
rect 21148 8444 21270 8476
rect 21000 8316 21270 8444
rect 21000 8284 21116 8316
rect 21148 8284 21270 8316
rect 21000 8156 21270 8284
rect 21000 8124 21116 8156
rect 21148 8124 21270 8156
rect 21000 7996 21270 8124
rect 21000 7964 21116 7996
rect 21148 7964 21270 7996
rect 21000 7836 21270 7964
rect 21000 7804 21116 7836
rect 21148 7804 21270 7836
rect 21000 7676 21270 7804
rect 21000 7644 21116 7676
rect 21148 7644 21270 7676
rect 21000 7516 21270 7644
rect 21000 7484 21116 7516
rect 21148 7484 21270 7516
rect 21000 7356 21270 7484
rect 21000 7324 21116 7356
rect 21148 7324 21270 7356
rect 21000 7196 21270 7324
rect 21000 7164 21116 7196
rect 21148 7164 21270 7196
rect 21000 7036 21270 7164
rect 21000 7004 21116 7036
rect 21148 7004 21270 7036
rect 18730 6876 19770 6905
rect 21000 6900 21270 7004
rect 18730 6844 18849 6876
rect 18881 6875 19770 6876
rect 18881 6844 19000 6875
rect 18730 6716 19000 6844
rect 18730 6684 18849 6716
rect 18881 6684 19000 6716
rect 18730 6556 19000 6684
rect 18730 6524 18849 6556
rect 18881 6524 19000 6556
rect 18730 6396 19000 6524
rect 18730 6364 18849 6396
rect 18881 6364 19000 6396
rect 18730 6236 19000 6364
rect 18730 6204 18849 6236
rect 18881 6204 19000 6236
rect 18730 6076 19000 6204
rect 18730 6044 18849 6076
rect 18881 6044 19000 6076
rect 18730 5916 19000 6044
rect 18730 5884 18849 5916
rect 18881 5884 19000 5916
rect 18730 5770 19000 5884
rect 15000 5756 19000 5770
rect 15000 5724 15116 5756
rect 15148 5724 18849 5756
rect 18881 5724 19000 5756
rect 15000 5653 19000 5724
rect 15000 5621 15304 5653
rect 15336 5621 15464 5653
rect 15496 5621 15624 5653
rect 15656 5621 15784 5653
rect 15816 5621 15944 5653
rect 15976 5621 16104 5653
rect 16136 5621 16264 5653
rect 16296 5621 16424 5653
rect 16456 5621 16584 5653
rect 16616 5621 16744 5653
rect 16776 5621 16904 5653
rect 16936 5621 17064 5653
rect 17096 5621 17224 5653
rect 17256 5621 17384 5653
rect 17416 5621 17544 5653
rect 17576 5621 17704 5653
rect 17736 5621 17864 5653
rect 17896 5621 18024 5653
rect 18056 5621 18184 5653
rect 18216 5621 18344 5653
rect 18376 5621 18504 5653
rect 18536 5621 18664 5653
rect 18696 5621 19000 5653
rect 15000 5500 19000 5621
rect 13850 5330 19700 5360
rect 6625 5120 13455 5160
rect 3000 3381 7000 3500
rect 3000 3349 3304 3381
rect 3336 3349 3464 3381
rect 3496 3349 3624 3381
rect 3656 3349 3784 3381
rect 3816 3349 3944 3381
rect 3976 3349 4104 3381
rect 4136 3349 4264 3381
rect 4296 3349 4424 3381
rect 4456 3349 4584 3381
rect 4616 3349 4744 3381
rect 4776 3349 4904 3381
rect 4936 3349 5064 3381
rect 5096 3349 5224 3381
rect 5256 3349 5384 3381
rect 5416 3349 5544 3381
rect 5576 3349 5704 3381
rect 5736 3349 5864 3381
rect 5896 3349 6024 3381
rect 6056 3349 6184 3381
rect 6216 3349 6344 3381
rect 6376 3349 6504 3381
rect 6536 3349 6664 3381
rect 6696 3349 7000 3381
rect 3000 3276 7000 3349
rect 3000 3244 3116 3276
rect 3148 3244 6849 3276
rect 6881 3244 7000 3276
rect 3000 3230 7000 3244
rect 3000 3116 3270 3230
rect 3000 3084 3116 3116
rect 3148 3084 3270 3116
rect 3000 2956 3270 3084
rect 3000 2924 3116 2956
rect 3148 2924 3270 2956
rect 3000 2796 3270 2924
rect 3000 2764 3116 2796
rect 3148 2764 3270 2796
rect 3000 2636 3270 2764
rect 3000 2604 3116 2636
rect 3148 2604 3270 2636
rect 3000 2476 3270 2604
rect 3000 2444 3116 2476
rect 3148 2444 3270 2476
rect 3000 2316 3270 2444
rect 3000 2284 3116 2316
rect 3148 2284 3270 2316
rect 3000 2156 3270 2284
rect 3000 2124 3116 2156
rect 3148 2124 3270 2156
rect 3000 1996 3270 2124
rect 3000 1964 3116 1996
rect 3148 1964 3270 1996
rect 3000 1836 3270 1964
rect 3000 1804 3116 1836
rect 3148 1804 3270 1836
rect 3000 1676 3270 1804
rect 3000 1644 3116 1676
rect 3148 1644 3270 1676
rect 3000 1516 3270 1644
rect 3000 1484 3116 1516
rect 3148 1484 3270 1516
rect 3000 1356 3270 1484
rect 3000 1324 3116 1356
rect 3148 1324 3270 1356
rect 3000 1196 3270 1324
rect 3000 1164 3116 1196
rect 3148 1164 3270 1196
rect 3000 1036 3270 1164
rect 3000 1004 3116 1036
rect 3148 1004 3270 1036
rect 3000 876 3270 1004
rect 3000 844 3116 876
rect 3148 844 3270 876
rect 3000 716 3270 844
rect 3000 684 3116 716
rect 3148 684 3270 716
rect 3000 556 3270 684
rect 3000 524 3116 556
rect 3148 524 3270 556
rect 3000 396 3270 524
rect 3000 364 3116 396
rect 3148 364 3270 396
rect 3000 236 3270 364
rect 3000 204 3116 236
rect 3148 204 3270 236
rect 3000 76 3270 204
rect 3000 44 3116 76
rect 3148 44 3270 76
rect 3000 -84 3270 44
rect 3000 -116 3116 -84
rect 3148 -116 3270 -84
rect 3000 -230 3270 -116
rect 6730 3116 7000 3230
rect 6730 3084 6849 3116
rect 6881 3084 7000 3116
rect 6730 2956 7000 3084
rect 6730 2924 6849 2956
rect 6881 2924 7000 2956
rect 6730 2796 7000 2924
rect 6730 2764 6849 2796
rect 6881 2764 7000 2796
rect 6730 2636 7000 2764
rect 6730 2604 6849 2636
rect 6881 2604 7000 2636
rect 6730 2476 7000 2604
rect 6730 2444 6849 2476
rect 6881 2444 7000 2476
rect 6730 2316 7000 2444
rect 6730 2284 6849 2316
rect 6881 2284 7000 2316
rect 6730 2156 7000 2284
rect 6730 2124 6849 2156
rect 6881 2124 7000 2156
rect 6730 1996 7000 2124
rect 6730 1964 6849 1996
rect 6881 1964 7000 1996
rect 6730 1836 7000 1964
rect 6730 1804 6849 1836
rect 6881 1804 7000 1836
rect 6730 1676 7000 1804
rect 6730 1644 6849 1676
rect 6881 1644 7000 1676
rect 6730 1516 7000 1644
rect 6730 1484 6849 1516
rect 6881 1484 7000 1516
rect 6730 1356 7000 1484
rect 6730 1324 6849 1356
rect 6881 1324 7000 1356
rect 6730 1196 7000 1324
rect 6730 1164 6849 1196
rect 6881 1164 7000 1196
rect 6730 1036 7000 1164
rect 6730 1004 6849 1036
rect 6881 1004 7000 1036
rect 6730 876 7000 1004
rect 6730 844 6849 876
rect 6881 844 7000 876
rect 6730 716 7000 844
rect 6730 684 6849 716
rect 6881 684 7000 716
rect 6730 556 7000 684
rect 6730 524 6849 556
rect 6881 524 7000 556
rect 6730 396 7000 524
rect 6730 364 6849 396
rect 6881 364 7000 396
rect 6730 236 7000 364
rect 6730 204 6849 236
rect 6881 204 7000 236
rect 6730 76 7000 204
rect 6730 44 6849 76
rect 6881 44 7000 76
rect 6730 -84 7000 44
rect 6730 -116 6849 -84
rect 6881 -116 7000 -84
rect 6730 -230 7000 -116
rect 3000 -244 7000 -230
rect 3000 -276 3116 -244
rect 3148 -276 6849 -244
rect 6881 -276 7000 -244
rect 3000 -347 7000 -276
rect 3000 -379 3304 -347
rect 3336 -379 3464 -347
rect 3496 -379 3624 -347
rect 3656 -379 3784 -347
rect 3816 -379 3944 -347
rect 3976 -379 4104 -347
rect 4136 -379 4264 -347
rect 4296 -379 4424 -347
rect 4456 -379 4584 -347
rect 4616 -379 4744 -347
rect 4776 -379 4904 -347
rect 4936 -379 5064 -347
rect 5096 -379 5224 -347
rect 5256 -379 5384 -347
rect 5416 -379 5544 -347
rect 5576 -379 5704 -347
rect 5736 -379 5864 -347
rect 5896 -379 6024 -347
rect 6056 -379 6184 -347
rect 6216 -379 6344 -347
rect 6376 -379 6504 -347
rect 6536 -379 6664 -347
rect 6696 -379 7000 -347
rect 3000 -500 7000 -379
rect 9000 3381 13000 3500
rect 9000 3349 9304 3381
rect 9336 3349 9464 3381
rect 9496 3349 9624 3381
rect 9656 3349 9784 3381
rect 9816 3349 9944 3381
rect 9976 3349 10104 3381
rect 10136 3349 10264 3381
rect 10296 3349 10424 3381
rect 10456 3349 10584 3381
rect 10616 3349 10744 3381
rect 10776 3349 10904 3381
rect 10936 3349 11064 3381
rect 11096 3349 11224 3381
rect 11256 3349 11384 3381
rect 11416 3349 11544 3381
rect 11576 3349 11704 3381
rect 11736 3349 11864 3381
rect 11896 3349 12024 3381
rect 12056 3349 12184 3381
rect 12216 3349 12344 3381
rect 12376 3349 12504 3381
rect 12536 3349 12664 3381
rect 12696 3349 13000 3381
rect 9000 3276 13000 3349
rect 9000 3244 9116 3276
rect 9148 3244 12849 3276
rect 12881 3244 13000 3276
rect 9000 3230 13000 3244
rect 9000 3116 9270 3230
rect 9000 3084 9116 3116
rect 9148 3084 9270 3116
rect 9000 2956 9270 3084
rect 9000 2924 9116 2956
rect 9148 2924 9270 2956
rect 9000 2796 9270 2924
rect 9000 2764 9116 2796
rect 9148 2764 9270 2796
rect 9000 2636 9270 2764
rect 9000 2604 9116 2636
rect 9148 2604 9270 2636
rect 9000 2476 9270 2604
rect 9000 2444 9116 2476
rect 9148 2444 9270 2476
rect 9000 2316 9270 2444
rect 9000 2284 9116 2316
rect 9148 2284 9270 2316
rect 9000 2156 9270 2284
rect 9000 2124 9116 2156
rect 9148 2124 9270 2156
rect 9000 1996 9270 2124
rect 9000 1964 9116 1996
rect 9148 1964 9270 1996
rect 9000 1836 9270 1964
rect 9000 1804 9116 1836
rect 9148 1804 9270 1836
rect 9000 1676 9270 1804
rect 9000 1644 9116 1676
rect 9148 1644 9270 1676
rect 9000 1516 9270 1644
rect 9000 1484 9116 1516
rect 9148 1484 9270 1516
rect 9000 1356 9270 1484
rect 9000 1324 9116 1356
rect 9148 1324 9270 1356
rect 9000 1196 9270 1324
rect 9000 1164 9116 1196
rect 9148 1164 9270 1196
rect 9000 1036 9270 1164
rect 9000 1004 9116 1036
rect 9148 1004 9270 1036
rect 9000 876 9270 1004
rect 9000 844 9116 876
rect 9148 844 9270 876
rect 9000 716 9270 844
rect 9000 684 9116 716
rect 9148 684 9270 716
rect 9000 556 9270 684
rect 9000 524 9116 556
rect 9148 524 9270 556
rect 9000 396 9270 524
rect 9000 364 9116 396
rect 9148 364 9270 396
rect 9000 236 9270 364
rect 9000 204 9116 236
rect 9148 204 9270 236
rect 9000 76 9270 204
rect 9000 44 9116 76
rect 9148 44 9270 76
rect 9000 -84 9270 44
rect 9000 -116 9116 -84
rect 9148 -116 9270 -84
rect 9000 -230 9270 -116
rect 12730 3116 13000 3230
rect 12730 3084 12849 3116
rect 12881 3084 13000 3116
rect 12730 2956 13000 3084
rect 12730 2924 12849 2956
rect 12881 2924 13000 2956
rect 12730 2796 13000 2924
rect 12730 2764 12849 2796
rect 12881 2764 13000 2796
rect 12730 2636 13000 2764
rect 12730 2604 12849 2636
rect 12881 2604 13000 2636
rect 12730 2476 13000 2604
rect 12730 2444 12849 2476
rect 12881 2444 13000 2476
rect 12730 2316 13000 2444
rect 12730 2284 12849 2316
rect 12881 2284 13000 2316
rect 12730 2156 13000 2284
rect 12730 2124 12849 2156
rect 12881 2124 13000 2156
rect 12730 1996 13000 2124
rect 12730 1964 12849 1996
rect 12881 1964 13000 1996
rect 12730 1836 13000 1964
rect 12730 1804 12849 1836
rect 12881 1804 13000 1836
rect 12730 1715 13000 1804
rect 13415 1835 13455 5120
rect 15000 3381 19000 3500
rect 15000 3349 15304 3381
rect 15336 3349 15464 3381
rect 15496 3349 15624 3381
rect 15656 3349 15784 3381
rect 15816 3349 15944 3381
rect 15976 3349 16104 3381
rect 16136 3349 16264 3381
rect 16296 3349 16424 3381
rect 16456 3349 16584 3381
rect 16616 3349 16744 3381
rect 16776 3349 16904 3381
rect 16936 3349 17064 3381
rect 17096 3349 17224 3381
rect 17256 3349 17384 3381
rect 17416 3349 17544 3381
rect 17576 3349 17704 3381
rect 17736 3349 17864 3381
rect 17896 3349 18024 3381
rect 18056 3349 18184 3381
rect 18216 3349 18344 3381
rect 18376 3349 18504 3381
rect 18536 3349 18664 3381
rect 18696 3349 19000 3381
rect 15000 3276 19000 3349
rect 15000 3244 15116 3276
rect 15148 3244 18849 3276
rect 18881 3244 19000 3276
rect 15000 3230 19000 3244
rect 15000 3116 15270 3230
rect 15000 3084 15116 3116
rect 15148 3084 15270 3116
rect 15000 2956 15270 3084
rect 15000 2924 15116 2956
rect 15148 2924 15270 2956
rect 15000 2796 15270 2924
rect 15000 2764 15116 2796
rect 15148 2764 15270 2796
rect 15000 2636 15270 2764
rect 15000 2604 15116 2636
rect 15148 2604 15270 2636
rect 15000 2476 15270 2604
rect 15000 2444 15116 2476
rect 15148 2444 15270 2476
rect 15000 2316 15270 2444
rect 15000 2284 15116 2316
rect 15148 2284 15270 2316
rect 15000 2156 15270 2284
rect 15000 2124 15116 2156
rect 15148 2124 15270 2156
rect 15000 1996 15270 2124
rect 15000 1964 15116 1996
rect 15148 1964 15270 1996
rect 15000 1836 15270 1964
rect 13415 1795 14800 1835
rect 12730 1676 14700 1715
rect 12730 1644 12849 1676
rect 12881 1675 14700 1676
rect 12881 1644 13000 1675
rect 12730 1516 13000 1644
rect 12730 1484 12849 1516
rect 12881 1484 13000 1516
rect 12730 1356 13000 1484
rect 12730 1324 12849 1356
rect 12881 1324 13000 1356
rect 12730 1196 13000 1324
rect 12730 1164 12849 1196
rect 12881 1164 13000 1196
rect 12730 1036 13000 1164
rect 12730 1004 12849 1036
rect 12881 1004 13000 1036
rect 12730 876 13000 1004
rect 12730 844 12849 876
rect 12881 844 13000 876
rect 12730 716 13000 844
rect 12730 684 12849 716
rect 12881 684 13000 716
rect 12730 556 13000 684
rect 12730 524 12849 556
rect 12881 524 13000 556
rect 12730 396 13000 524
rect 12730 364 12849 396
rect 12881 364 13000 396
rect 12730 236 13000 364
rect 12730 204 12849 236
rect 12881 204 13000 236
rect 12730 76 13000 204
rect 12730 44 12849 76
rect 12881 44 13000 76
rect 12730 -84 13000 44
rect 12730 -116 12849 -84
rect 12881 -116 13000 -84
rect 12730 -230 13000 -116
rect 9000 -244 13000 -230
rect 9000 -276 9116 -244
rect 9148 -276 12849 -244
rect 12881 -276 13000 -244
rect 9000 -347 13000 -276
rect 9000 -379 9304 -347
rect 9336 -379 9464 -347
rect 9496 -379 9624 -347
rect 9656 -379 9784 -347
rect 9816 -379 9944 -347
rect 9976 -379 10104 -347
rect 10136 -379 10264 -347
rect 10296 -379 10424 -347
rect 10456 -379 10584 -347
rect 10616 -379 10744 -347
rect 10776 -379 10904 -347
rect 10936 -379 11064 -347
rect 11096 -379 11224 -347
rect 11256 -379 11384 -347
rect 11416 -379 11544 -347
rect 11576 -379 11704 -347
rect 11736 -379 11864 -347
rect 11896 -379 12024 -347
rect 12056 -379 12184 -347
rect 12216 -379 12344 -347
rect 12376 -379 12504 -347
rect 12536 -379 12664 -347
rect 12696 -379 13000 -347
rect 9000 -500 13000 -379
rect 14660 -660 14700 1675
rect 14760 -560 14800 1795
rect 15000 1804 15116 1836
rect 15148 1804 15270 1836
rect 15000 1676 15270 1804
rect 15000 1644 15116 1676
rect 15148 1644 15270 1676
rect 15000 1516 15270 1644
rect 15000 1484 15116 1516
rect 15148 1484 15270 1516
rect 15000 1356 15270 1484
rect 15000 1324 15116 1356
rect 15148 1324 15270 1356
rect 15000 1196 15270 1324
rect 15000 1164 15116 1196
rect 15148 1164 15270 1196
rect 15000 1036 15270 1164
rect 15000 1004 15116 1036
rect 15148 1004 15270 1036
rect 15000 876 15270 1004
rect 15000 844 15116 876
rect 15148 844 15270 876
rect 15000 716 15270 844
rect 15000 684 15116 716
rect 15148 684 15270 716
rect 15000 556 15270 684
rect 15000 524 15116 556
rect 15148 524 15270 556
rect 15000 396 15270 524
rect 15000 364 15116 396
rect 15148 364 15270 396
rect 15000 236 15270 364
rect 15000 204 15116 236
rect 15148 204 15270 236
rect 15000 76 15270 204
rect 15000 44 15116 76
rect 15148 44 15270 76
rect 15000 -84 15270 44
rect 15000 -116 15116 -84
rect 15148 -116 15270 -84
rect 15000 -230 15270 -116
rect 18730 3116 19000 3230
rect 18730 3084 18849 3116
rect 18881 3084 19000 3116
rect 18730 2956 19000 3084
rect 18730 2924 18849 2956
rect 18881 2924 19000 2956
rect 18730 2796 19000 2924
rect 18730 2764 18849 2796
rect 18881 2764 19000 2796
rect 18730 2636 19000 2764
rect 18730 2604 18849 2636
rect 18881 2604 19000 2636
rect 18730 2476 19000 2604
rect 18730 2444 18849 2476
rect 18881 2444 19000 2476
rect 18730 2316 19000 2444
rect 18730 2284 18849 2316
rect 18881 2284 19000 2316
rect 18730 2156 19000 2284
rect 18730 2124 18849 2156
rect 18881 2124 19000 2156
rect 18730 1996 19000 2124
rect 18730 1964 18849 1996
rect 18881 1964 19000 1996
rect 18730 1836 19000 1964
rect 18730 1804 18849 1836
rect 18881 1804 19000 1836
rect 18730 1676 19000 1804
rect 18730 1644 18849 1676
rect 18881 1644 19000 1676
rect 18730 1516 19000 1644
rect 18730 1484 18849 1516
rect 18881 1484 19000 1516
rect 18730 1356 19000 1484
rect 18730 1324 18849 1356
rect 18881 1324 19000 1356
rect 18730 1196 19000 1324
rect 18730 1164 18849 1196
rect 18881 1164 19000 1196
rect 18730 1036 19000 1164
rect 18730 1004 18849 1036
rect 18881 1004 19000 1036
rect 18730 876 19000 1004
rect 18730 844 18849 876
rect 18881 844 19000 876
rect 18730 716 19000 844
rect 18730 684 18849 716
rect 18881 684 19000 716
rect 18730 556 19000 684
rect 18730 524 18849 556
rect 18881 524 19000 556
rect 18730 396 19000 524
rect 18730 364 18849 396
rect 18881 364 19000 396
rect 18730 236 19000 364
rect 18730 204 18849 236
rect 18881 204 19000 236
rect 18730 76 19000 204
rect 18730 44 18849 76
rect 18881 44 19000 76
rect 18730 -84 19000 44
rect 18730 -116 18849 -84
rect 18881 -116 19000 -84
rect 18730 -230 19000 -116
rect 15000 -244 19000 -230
rect 15000 -276 15116 -244
rect 15148 -276 18849 -244
rect 18881 -276 19000 -244
rect 15000 -347 19000 -276
rect 15000 -379 15304 -347
rect 15336 -379 15464 -347
rect 15496 -379 15624 -347
rect 15656 -379 15784 -347
rect 15816 -379 15944 -347
rect 15976 -379 16104 -347
rect 16136 -379 16264 -347
rect 16296 -379 16424 -347
rect 16456 -379 16584 -347
rect 16616 -379 16744 -347
rect 16776 -379 16904 -347
rect 16936 -379 17064 -347
rect 17096 -379 17224 -347
rect 17256 -379 17384 -347
rect 17416 -379 17544 -347
rect 17576 -379 17704 -347
rect 17736 -379 17864 -347
rect 17896 -379 18024 -347
rect 18056 -379 18184 -347
rect 18216 -379 18344 -347
rect 18376 -379 18504 -347
rect 18536 -379 18664 -347
rect 18696 -379 19000 -347
rect 15000 -500 19000 -379
rect 14760 -600 15940 -560
rect 14660 -700 15835 -660
rect 15795 -2225 15835 -700
rect 15900 -2065 15940 -600
rect 19670 -625 19700 5330
rect 19430 -630 19700 -625
rect 19430 -690 19440 -630
rect 19480 -690 19700 -630
rect 19430 -695 19700 -690
rect 19670 -1015 19700 -695
rect 19740 -955 19770 6875
rect 19805 6876 21270 6900
rect 19805 6870 21116 6876
rect 19805 -895 19835 6870
rect 21000 6844 21116 6870
rect 21148 6844 21270 6876
rect 21000 6716 21270 6844
rect 21000 6684 21116 6716
rect 21148 6684 21270 6716
rect 21000 6556 21270 6684
rect 21000 6524 21116 6556
rect 21148 6524 21270 6556
rect 21000 6396 21270 6524
rect 21000 6364 21116 6396
rect 21148 6364 21270 6396
rect 21000 6236 21270 6364
rect 21000 6204 21116 6236
rect 21148 6204 21270 6236
rect 21000 6076 21270 6204
rect 21000 6044 21116 6076
rect 21148 6044 21270 6076
rect 21000 5916 21270 6044
rect 21000 5884 21116 5916
rect 21148 5884 21270 5916
rect 21000 5770 21270 5884
rect 24730 9116 25000 9230
rect 24730 9084 24849 9116
rect 24881 9084 25000 9116
rect 24730 8956 25000 9084
rect 24730 8924 24849 8956
rect 24881 8924 25000 8956
rect 24730 8796 25000 8924
rect 24730 8764 24849 8796
rect 24881 8764 25000 8796
rect 24730 8636 25000 8764
rect 24730 8604 24849 8636
rect 24881 8604 25000 8636
rect 24730 8476 25000 8604
rect 24730 8444 24849 8476
rect 24881 8444 25000 8476
rect 24730 8316 25000 8444
rect 24730 8284 24849 8316
rect 24881 8284 25000 8316
rect 24730 8156 25000 8284
rect 24730 8124 24849 8156
rect 24881 8124 25000 8156
rect 24730 7996 25000 8124
rect 24730 7964 24849 7996
rect 24881 7964 25000 7996
rect 24730 7836 25000 7964
rect 24730 7804 24849 7836
rect 24881 7804 25000 7836
rect 24730 7676 25000 7804
rect 24730 7644 24849 7676
rect 24881 7644 25000 7676
rect 24730 7516 25000 7644
rect 24730 7484 24849 7516
rect 24881 7484 25000 7516
rect 24730 7356 25000 7484
rect 24730 7324 24849 7356
rect 24881 7324 25000 7356
rect 24730 7196 25000 7324
rect 24730 7164 24849 7196
rect 24881 7164 25000 7196
rect 24730 7036 25000 7164
rect 24730 7004 24849 7036
rect 24881 7004 25000 7036
rect 24730 6876 25000 7004
rect 24730 6844 24849 6876
rect 24881 6844 25000 6876
rect 24730 6716 25000 6844
rect 24730 6684 24849 6716
rect 24881 6684 25000 6716
rect 24730 6556 25000 6684
rect 24730 6524 24849 6556
rect 24881 6524 25000 6556
rect 24730 6396 25000 6524
rect 24730 6364 24849 6396
rect 24881 6364 25000 6396
rect 24730 6236 25000 6364
rect 24730 6204 24849 6236
rect 24881 6204 25000 6236
rect 24730 6076 25000 6204
rect 24730 6044 24849 6076
rect 24881 6044 25000 6076
rect 24730 5916 25000 6044
rect 24730 5884 24849 5916
rect 24881 5884 25000 5916
rect 24730 5770 25000 5884
rect 21000 5756 25000 5770
rect 21000 5724 21116 5756
rect 21148 5724 24849 5756
rect 24881 5724 25000 5756
rect 21000 5653 25000 5724
rect 21000 5621 21304 5653
rect 21336 5621 21464 5653
rect 21496 5621 21624 5653
rect 21656 5621 21784 5653
rect 21816 5621 21944 5653
rect 21976 5621 22104 5653
rect 22136 5621 22264 5653
rect 22296 5621 22424 5653
rect 22456 5621 22584 5653
rect 22616 5621 22744 5653
rect 22776 5621 22904 5653
rect 22936 5621 23064 5653
rect 23096 5621 23224 5653
rect 23256 5621 23384 5653
rect 23416 5621 23544 5653
rect 23576 5621 23704 5653
rect 23736 5621 23864 5653
rect 23896 5621 24024 5653
rect 24056 5621 24184 5653
rect 24216 5621 24344 5653
rect 24376 5621 24504 5653
rect 24536 5621 24664 5653
rect 24696 5621 25000 5653
rect 21000 5500 25000 5621
rect 21000 3381 25000 3500
rect 21000 3349 21304 3381
rect 21336 3349 21464 3381
rect 21496 3349 21624 3381
rect 21656 3349 21784 3381
rect 21816 3349 21944 3381
rect 21976 3349 22104 3381
rect 22136 3349 22264 3381
rect 22296 3349 22424 3381
rect 22456 3349 22584 3381
rect 22616 3349 22744 3381
rect 22776 3349 22904 3381
rect 22936 3349 23064 3381
rect 23096 3349 23224 3381
rect 23256 3349 23384 3381
rect 23416 3349 23544 3381
rect 23576 3349 23704 3381
rect 23736 3349 23864 3381
rect 23896 3349 24024 3381
rect 24056 3349 24184 3381
rect 24216 3349 24344 3381
rect 24376 3349 24504 3381
rect 24536 3349 24664 3381
rect 24696 3349 25000 3381
rect 21000 3276 25000 3349
rect 21000 3244 21116 3276
rect 21148 3244 24849 3276
rect 24881 3244 25000 3276
rect 21000 3230 25000 3244
rect 21000 3116 21270 3230
rect 21000 3084 21116 3116
rect 21148 3084 21270 3116
rect 21000 2956 21270 3084
rect 21000 2924 21116 2956
rect 21148 2924 21270 2956
rect 21000 2796 21270 2924
rect 21000 2764 21116 2796
rect 21148 2764 21270 2796
rect 21000 2636 21270 2764
rect 21000 2604 21116 2636
rect 21148 2604 21270 2636
rect 21000 2476 21270 2604
rect 21000 2444 21116 2476
rect 21148 2444 21270 2476
rect 21000 2316 21270 2444
rect 21000 2284 21116 2316
rect 21148 2284 21270 2316
rect 21000 2156 21270 2284
rect 21000 2124 21116 2156
rect 21148 2124 21270 2156
rect 21000 1996 21270 2124
rect 21000 1964 21116 1996
rect 21148 1964 21270 1996
rect 21000 1836 21270 1964
rect 21000 1804 21116 1836
rect 21148 1804 21270 1836
rect 21000 1676 21270 1804
rect 21000 1644 21116 1676
rect 21148 1644 21270 1676
rect 21000 1516 21270 1644
rect 21000 1484 21116 1516
rect 21148 1484 21270 1516
rect 21000 1356 21270 1484
rect 21000 1324 21116 1356
rect 21148 1324 21270 1356
rect 21000 1196 21270 1324
rect 21000 1164 21116 1196
rect 21148 1164 21270 1196
rect 21000 1036 21270 1164
rect 21000 1004 21116 1036
rect 21148 1004 21270 1036
rect 21000 876 21270 1004
rect 21000 844 21116 876
rect 21148 844 21270 876
rect 21000 716 21270 844
rect 21000 684 21116 716
rect 21148 684 21270 716
rect 21000 556 21270 684
rect 21000 524 21116 556
rect 21148 524 21270 556
rect 21000 396 21270 524
rect 21000 364 21116 396
rect 21148 364 21270 396
rect 21000 236 21270 364
rect 21000 204 21116 236
rect 21148 204 21270 236
rect 21000 76 21270 204
rect 21000 44 21116 76
rect 21148 44 21270 76
rect 21000 -84 21270 44
rect 21000 -116 21116 -84
rect 21148 -116 21270 -84
rect 21000 -230 21270 -116
rect 24730 3116 25000 3230
rect 24730 3084 24849 3116
rect 24881 3084 25000 3116
rect 24730 2956 25000 3084
rect 24730 2924 24849 2956
rect 24881 2924 25000 2956
rect 24730 2796 25000 2924
rect 24730 2764 24849 2796
rect 24881 2764 25000 2796
rect 24730 2636 25000 2764
rect 24730 2604 24849 2636
rect 24881 2604 25000 2636
rect 24730 2476 25000 2604
rect 24730 2444 24849 2476
rect 24881 2444 25000 2476
rect 24730 2316 25000 2444
rect 24730 2284 24849 2316
rect 24881 2284 25000 2316
rect 24730 2156 25000 2284
rect 24730 2124 24849 2156
rect 24881 2124 25000 2156
rect 24730 1996 25000 2124
rect 24730 1964 24849 1996
rect 24881 1964 25000 1996
rect 24730 1836 25000 1964
rect 24730 1804 24849 1836
rect 24881 1804 25000 1836
rect 24730 1676 25000 1804
rect 24730 1644 24849 1676
rect 24881 1644 25000 1676
rect 24730 1516 25000 1644
rect 24730 1484 24849 1516
rect 24881 1484 25000 1516
rect 24730 1356 25000 1484
rect 24730 1324 24849 1356
rect 24881 1324 25000 1356
rect 24730 1196 25000 1324
rect 24730 1164 24849 1196
rect 24881 1164 25000 1196
rect 24730 1036 25000 1164
rect 24730 1004 24849 1036
rect 24881 1004 25000 1036
rect 24730 876 25000 1004
rect 24730 844 24849 876
rect 24881 844 25000 876
rect 24730 716 25000 844
rect 24730 684 24849 716
rect 24881 684 25000 716
rect 24730 556 25000 684
rect 24730 524 24849 556
rect 24881 524 25000 556
rect 24730 396 25000 524
rect 24730 364 24849 396
rect 24881 364 25000 396
rect 24730 236 25000 364
rect 24730 204 24849 236
rect 24881 204 25000 236
rect 24730 76 25000 204
rect 24730 44 24849 76
rect 24881 44 25000 76
rect 24730 -84 25000 44
rect 24730 -116 24849 -84
rect 24881 -116 25000 -84
rect 24730 -230 25000 -116
rect 21000 -244 25000 -230
rect 21000 -276 21116 -244
rect 21148 -276 24849 -244
rect 24881 -276 25000 -244
rect 21000 -347 25000 -276
rect 21000 -379 21304 -347
rect 21336 -379 21464 -347
rect 21496 -379 21624 -347
rect 21656 -379 21784 -347
rect 21816 -379 21944 -347
rect 21976 -379 22104 -347
rect 22136 -379 22264 -347
rect 22296 -379 22424 -347
rect 22456 -379 22584 -347
rect 22616 -379 22744 -347
rect 22776 -379 22904 -347
rect 22936 -379 23064 -347
rect 23096 -379 23224 -347
rect 23256 -379 23384 -347
rect 23416 -379 23544 -347
rect 23576 -379 23704 -347
rect 23736 -379 23864 -347
rect 23896 -379 24024 -347
rect 24056 -379 24184 -347
rect 24216 -379 24344 -347
rect 24376 -379 24504 -347
rect 24536 -379 24664 -347
rect 24696 -379 25000 -347
rect 21000 -500 25000 -379
rect 19805 -925 20135 -895
rect 19740 -985 20070 -955
rect 19670 -1045 20000 -1015
rect 19970 -1210 20000 -1045
rect 20040 -1135 20070 -985
rect 20030 -1140 20070 -1135
rect 20030 -1170 20035 -1140
rect 20065 -1170 20070 -1140
rect 20030 -1175 20070 -1170
rect 20105 -1205 20135 -925
rect 19960 -1215 20000 -1210
rect 19960 -1245 19965 -1215
rect 19995 -1245 20000 -1215
rect 20065 -1210 20135 -1205
rect 20065 -1240 20070 -1210
rect 20100 -1240 20135 -1210
rect 20065 -1245 20135 -1240
rect 19960 -1250 20000 -1245
rect 16315 -1870 17520 -1830
rect 16315 -2065 16355 -1870
rect 15900 -2070 16355 -2065
rect 15900 -2100 16155 -2070
rect 16225 -2100 16355 -2070
rect 15900 -2105 16355 -2100
rect 16420 -1950 17440 -1910
rect 16420 -2225 16460 -1950
rect 15795 -2230 16460 -2225
rect 15795 -2260 16295 -2230
rect 16365 -2260 16460 -2230
rect 15795 -2265 16460 -2260
rect 17400 -2570 17440 -1950
rect 17480 -2495 17520 -1870
rect 17480 -2535 18070 -2495
rect 17400 -2610 17970 -2570
rect 17930 -2675 17970 -2610
rect 18030 -2675 18070 -2535
rect 9930 -3465 9970 -3325
rect 10030 -3390 10070 -3325
rect 10030 -3430 10600 -3390
rect 9930 -3505 10520 -3465
rect 10480 -4130 10520 -3505
rect 10560 -4050 10600 -3430
rect 11540 -3740 12205 -3735
rect 11540 -3770 11635 -3740
rect 11705 -3770 12205 -3740
rect 11540 -3775 12205 -3770
rect 11540 -4050 11580 -3775
rect 10560 -4090 11580 -4050
rect 11645 -3900 12100 -3895
rect 11645 -3930 11775 -3900
rect 11845 -3930 12100 -3900
rect 11645 -3935 12100 -3930
rect 11645 -4130 11685 -3935
rect 10480 -4170 11685 -4130
rect 8300 -4755 8340 -4750
rect 8165 -4760 8235 -4755
rect 8165 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8165 -4795 8235 -4790
rect 8300 -4785 8305 -4755
rect 8335 -4785 8340 -4755
rect 8300 -4790 8340 -4785
rect 3000 -5621 7000 -5500
rect 3000 -5653 3304 -5621
rect 3336 -5653 3464 -5621
rect 3496 -5653 3624 -5621
rect 3656 -5653 3784 -5621
rect 3816 -5653 3944 -5621
rect 3976 -5653 4104 -5621
rect 4136 -5653 4264 -5621
rect 4296 -5653 4424 -5621
rect 4456 -5653 4584 -5621
rect 4616 -5653 4744 -5621
rect 4776 -5653 4904 -5621
rect 4936 -5653 5064 -5621
rect 5096 -5653 5224 -5621
rect 5256 -5653 5384 -5621
rect 5416 -5653 5544 -5621
rect 5576 -5653 5704 -5621
rect 5736 -5653 5864 -5621
rect 5896 -5653 6024 -5621
rect 6056 -5653 6184 -5621
rect 6216 -5653 6344 -5621
rect 6376 -5653 6504 -5621
rect 6536 -5653 6664 -5621
rect 6696 -5653 7000 -5621
rect 3000 -5724 7000 -5653
rect 3000 -5756 3119 -5724
rect 3151 -5756 6852 -5724
rect 6884 -5756 7000 -5724
rect 3000 -5770 7000 -5756
rect 3000 -5884 3270 -5770
rect 3000 -5916 3119 -5884
rect 3151 -5916 3270 -5884
rect 3000 -6044 3270 -5916
rect 3000 -6076 3119 -6044
rect 3151 -6076 3270 -6044
rect 3000 -6204 3270 -6076
rect 3000 -6236 3119 -6204
rect 3151 -6236 3270 -6204
rect 3000 -6364 3270 -6236
rect 3000 -6396 3119 -6364
rect 3151 -6396 3270 -6364
rect 3000 -6524 3270 -6396
rect 3000 -6556 3119 -6524
rect 3151 -6556 3270 -6524
rect 3000 -6684 3270 -6556
rect 3000 -6716 3119 -6684
rect 3151 -6716 3270 -6684
rect 3000 -6844 3270 -6716
rect 3000 -6876 3119 -6844
rect 3151 -6876 3270 -6844
rect 3000 -7004 3270 -6876
rect 3000 -7036 3119 -7004
rect 3151 -7036 3270 -7004
rect 3000 -7164 3270 -7036
rect 3000 -7196 3119 -7164
rect 3151 -7196 3270 -7164
rect 3000 -7324 3270 -7196
rect 3000 -7356 3119 -7324
rect 3151 -7356 3270 -7324
rect 3000 -7484 3270 -7356
rect 3000 -7516 3119 -7484
rect 3151 -7516 3270 -7484
rect 3000 -7644 3270 -7516
rect 3000 -7676 3119 -7644
rect 3151 -7676 3270 -7644
rect 3000 -7804 3270 -7676
rect 3000 -7836 3119 -7804
rect 3151 -7836 3270 -7804
rect 3000 -7964 3270 -7836
rect 3000 -7996 3119 -7964
rect 3151 -7996 3270 -7964
rect 3000 -8124 3270 -7996
rect 3000 -8156 3119 -8124
rect 3151 -8156 3270 -8124
rect 3000 -8284 3270 -8156
rect 3000 -8316 3119 -8284
rect 3151 -8316 3270 -8284
rect 3000 -8444 3270 -8316
rect 3000 -8476 3119 -8444
rect 3151 -8476 3270 -8444
rect 3000 -8604 3270 -8476
rect 3000 -8636 3119 -8604
rect 3151 -8636 3270 -8604
rect 3000 -8764 3270 -8636
rect 3000 -8796 3119 -8764
rect 3151 -8796 3270 -8764
rect 3000 -8924 3270 -8796
rect 3000 -8956 3119 -8924
rect 3151 -8956 3270 -8924
rect 3000 -9084 3270 -8956
rect 3000 -9116 3119 -9084
rect 3151 -9116 3270 -9084
rect 3000 -9230 3270 -9116
rect 6730 -5884 7000 -5770
rect 6730 -5916 6852 -5884
rect 6884 -5916 7000 -5884
rect 6730 -6044 7000 -5916
rect 6730 -6076 6852 -6044
rect 6884 -6076 7000 -6044
rect 6730 -6204 7000 -6076
rect 6730 -6236 6852 -6204
rect 6884 -6236 7000 -6204
rect 6730 -6364 7000 -6236
rect 6730 -6396 6852 -6364
rect 6884 -6396 7000 -6364
rect 6730 -6524 7000 -6396
rect 6730 -6556 6852 -6524
rect 6884 -6556 7000 -6524
rect 6730 -6684 7000 -6556
rect 6730 -6716 6852 -6684
rect 6884 -6716 7000 -6684
rect 6730 -6844 7000 -6716
rect 6730 -6876 6852 -6844
rect 6884 -6876 7000 -6844
rect 6730 -7004 7000 -6876
rect 6730 -7036 6852 -7004
rect 6884 -7036 7000 -7004
rect 6730 -7164 7000 -7036
rect 6730 -7196 6852 -7164
rect 6884 -7196 7000 -7164
rect 6730 -7324 7000 -7196
rect 6730 -7356 6852 -7324
rect 6884 -7356 7000 -7324
rect 6730 -7484 7000 -7356
rect 6730 -7516 6852 -7484
rect 6884 -7516 7000 -7484
rect 6730 -7644 7000 -7516
rect 6730 -7676 6852 -7644
rect 6884 -7676 7000 -7644
rect 6730 -7804 7000 -7676
rect 6730 -7836 6852 -7804
rect 6884 -7836 7000 -7804
rect 6730 -7964 7000 -7836
rect 6730 -7996 6852 -7964
rect 6884 -7996 7000 -7964
rect 6730 -8124 7000 -7996
rect 6730 -8156 6852 -8124
rect 6884 -8156 7000 -8124
rect 6730 -8284 7000 -8156
rect 6730 -8316 6852 -8284
rect 6884 -8316 7000 -8284
rect 6730 -8444 7000 -8316
rect 6730 -8476 6852 -8444
rect 6884 -8476 7000 -8444
rect 6730 -8604 7000 -8476
rect 6730 -8636 6852 -8604
rect 6884 -8636 7000 -8604
rect 6730 -8764 7000 -8636
rect 6730 -8796 6852 -8764
rect 6884 -8796 7000 -8764
rect 6730 -8924 7000 -8796
rect 6730 -8956 6852 -8924
rect 6884 -8956 7000 -8924
rect 6730 -9084 7000 -8956
rect 6730 -9116 6852 -9084
rect 6884 -9116 7000 -9084
rect 6730 -9230 7000 -9116
rect 3000 -9244 7000 -9230
rect 3000 -9276 3119 -9244
rect 3151 -9276 6852 -9244
rect 6884 -9276 7000 -9244
rect 3000 -9349 7000 -9276
rect 3000 -9381 3304 -9349
rect 3336 -9381 3464 -9349
rect 3496 -9381 3624 -9349
rect 3656 -9381 3784 -9349
rect 3816 -9381 3944 -9349
rect 3976 -9381 4104 -9349
rect 4136 -9381 4264 -9349
rect 4296 -9381 4424 -9349
rect 4456 -9381 4584 -9349
rect 4616 -9381 4744 -9349
rect 4776 -9381 4904 -9349
rect 4936 -9381 5064 -9349
rect 5096 -9381 5224 -9349
rect 5256 -9381 5384 -9349
rect 5416 -9381 5544 -9349
rect 5576 -9381 5704 -9349
rect 5736 -9381 5864 -9349
rect 5896 -9381 6024 -9349
rect 6056 -9381 6184 -9349
rect 6216 -9381 6344 -9349
rect 6376 -9381 6504 -9349
rect 6536 -9381 6664 -9349
rect 6696 -9381 7000 -9349
rect 3000 -9500 7000 -9381
rect 3000 -11621 7000 -11500
rect 3000 -11653 3304 -11621
rect 3336 -11653 3464 -11621
rect 3496 -11653 3624 -11621
rect 3656 -11653 3784 -11621
rect 3816 -11653 3944 -11621
rect 3976 -11653 4104 -11621
rect 4136 -11653 4264 -11621
rect 4296 -11653 4424 -11621
rect 4456 -11653 4584 -11621
rect 4616 -11653 4744 -11621
rect 4776 -11653 4904 -11621
rect 4936 -11653 5064 -11621
rect 5096 -11653 5224 -11621
rect 5256 -11653 5384 -11621
rect 5416 -11653 5544 -11621
rect 5576 -11653 5704 -11621
rect 5736 -11653 5864 -11621
rect 5896 -11653 6024 -11621
rect 6056 -11653 6184 -11621
rect 6216 -11653 6344 -11621
rect 6376 -11653 6504 -11621
rect 6536 -11653 6664 -11621
rect 6696 -11653 7000 -11621
rect 3000 -11724 7000 -11653
rect 3000 -11756 3119 -11724
rect 3151 -11756 6852 -11724
rect 6884 -11756 7000 -11724
rect 3000 -11770 7000 -11756
rect 3000 -11884 3270 -11770
rect 3000 -11916 3119 -11884
rect 3151 -11916 3270 -11884
rect 3000 -12044 3270 -11916
rect 3000 -12076 3119 -12044
rect 3151 -12076 3270 -12044
rect 3000 -12204 3270 -12076
rect 3000 -12236 3119 -12204
rect 3151 -12236 3270 -12204
rect 3000 -12364 3270 -12236
rect 3000 -12396 3119 -12364
rect 3151 -12396 3270 -12364
rect 3000 -12524 3270 -12396
rect 3000 -12556 3119 -12524
rect 3151 -12556 3270 -12524
rect 3000 -12684 3270 -12556
rect 3000 -12716 3119 -12684
rect 3151 -12716 3270 -12684
rect 3000 -12844 3270 -12716
rect 3000 -12876 3119 -12844
rect 3151 -12876 3270 -12844
rect 3000 -13004 3270 -12876
rect 3000 -13036 3119 -13004
rect 3151 -13036 3270 -13004
rect 3000 -13164 3270 -13036
rect 3000 -13196 3119 -13164
rect 3151 -13196 3270 -13164
rect 3000 -13324 3270 -13196
rect 3000 -13356 3119 -13324
rect 3151 -13356 3270 -13324
rect 3000 -13484 3270 -13356
rect 3000 -13516 3119 -13484
rect 3151 -13516 3270 -13484
rect 3000 -13644 3270 -13516
rect 3000 -13676 3119 -13644
rect 3151 -13676 3270 -13644
rect 3000 -13804 3270 -13676
rect 3000 -13836 3119 -13804
rect 3151 -13836 3270 -13804
rect 3000 -13964 3270 -13836
rect 3000 -13996 3119 -13964
rect 3151 -13996 3270 -13964
rect 3000 -14124 3270 -13996
rect 3000 -14156 3119 -14124
rect 3151 -14156 3270 -14124
rect 3000 -14284 3270 -14156
rect 3000 -14316 3119 -14284
rect 3151 -14316 3270 -14284
rect 3000 -14444 3270 -14316
rect 3000 -14476 3119 -14444
rect 3151 -14476 3270 -14444
rect 3000 -14604 3270 -14476
rect 3000 -14636 3119 -14604
rect 3151 -14636 3270 -14604
rect 3000 -14764 3270 -14636
rect 3000 -14796 3119 -14764
rect 3151 -14796 3270 -14764
rect 3000 -14924 3270 -14796
rect 3000 -14956 3119 -14924
rect 3151 -14956 3270 -14924
rect 3000 -15084 3270 -14956
rect 3000 -15116 3119 -15084
rect 3151 -15116 3270 -15084
rect 3000 -15230 3270 -15116
rect 6730 -11884 7000 -11770
rect 6730 -11916 6852 -11884
rect 6884 -11916 7000 -11884
rect 6730 -12044 7000 -11916
rect 6730 -12076 6852 -12044
rect 6884 -12076 7000 -12044
rect 6730 -12204 7000 -12076
rect 6730 -12236 6852 -12204
rect 6884 -12236 7000 -12204
rect 6730 -12364 7000 -12236
rect 6730 -12396 6852 -12364
rect 6884 -12396 7000 -12364
rect 6730 -12524 7000 -12396
rect 6730 -12556 6852 -12524
rect 6884 -12556 7000 -12524
rect 6730 -12684 7000 -12556
rect 6730 -12716 6852 -12684
rect 6884 -12716 7000 -12684
rect 6730 -12844 7000 -12716
rect 6730 -12876 6852 -12844
rect 6884 -12870 7000 -12844
rect 8165 -12870 8195 -4795
rect 6884 -12876 8195 -12870
rect 6730 -12900 8195 -12876
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 8230 -12875 8260 -4865
rect 8300 -5305 8330 -4790
rect 8300 -5310 8570 -5305
rect 8300 -5370 8520 -5310
rect 8560 -5370 8570 -5310
rect 8300 -5375 8570 -5370
rect 8300 -11330 8330 -5375
rect 12060 -5400 12100 -3935
rect 12165 -5300 12205 -3775
rect 12165 -5340 13340 -5300
rect 12060 -5440 13240 -5400
rect 9000 -5621 13000 -5500
rect 9000 -5653 9304 -5621
rect 9336 -5653 9464 -5621
rect 9496 -5653 9624 -5621
rect 9656 -5653 9784 -5621
rect 9816 -5653 9944 -5621
rect 9976 -5653 10104 -5621
rect 10136 -5653 10264 -5621
rect 10296 -5653 10424 -5621
rect 10456 -5653 10584 -5621
rect 10616 -5653 10744 -5621
rect 10776 -5653 10904 -5621
rect 10936 -5653 11064 -5621
rect 11096 -5653 11224 -5621
rect 11256 -5653 11384 -5621
rect 11416 -5653 11544 -5621
rect 11576 -5653 11704 -5621
rect 11736 -5653 11864 -5621
rect 11896 -5653 12024 -5621
rect 12056 -5653 12184 -5621
rect 12216 -5653 12344 -5621
rect 12376 -5653 12504 -5621
rect 12536 -5653 12664 -5621
rect 12696 -5653 13000 -5621
rect 9000 -5724 13000 -5653
rect 9000 -5756 9119 -5724
rect 9151 -5756 12852 -5724
rect 12884 -5756 13000 -5724
rect 9000 -5770 13000 -5756
rect 9000 -5884 9270 -5770
rect 9000 -5916 9119 -5884
rect 9151 -5916 9270 -5884
rect 9000 -6044 9270 -5916
rect 9000 -6076 9119 -6044
rect 9151 -6076 9270 -6044
rect 9000 -6204 9270 -6076
rect 9000 -6236 9119 -6204
rect 9151 -6236 9270 -6204
rect 9000 -6364 9270 -6236
rect 9000 -6396 9119 -6364
rect 9151 -6396 9270 -6364
rect 9000 -6524 9270 -6396
rect 9000 -6556 9119 -6524
rect 9151 -6556 9270 -6524
rect 9000 -6684 9270 -6556
rect 9000 -6716 9119 -6684
rect 9151 -6716 9270 -6684
rect 9000 -6844 9270 -6716
rect 9000 -6876 9119 -6844
rect 9151 -6876 9270 -6844
rect 9000 -7004 9270 -6876
rect 9000 -7036 9119 -7004
rect 9151 -7036 9270 -7004
rect 9000 -7164 9270 -7036
rect 9000 -7196 9119 -7164
rect 9151 -7196 9270 -7164
rect 9000 -7324 9270 -7196
rect 9000 -7356 9119 -7324
rect 9151 -7356 9270 -7324
rect 9000 -7484 9270 -7356
rect 9000 -7516 9119 -7484
rect 9151 -7516 9270 -7484
rect 9000 -7644 9270 -7516
rect 9000 -7676 9119 -7644
rect 9151 -7676 9270 -7644
rect 9000 -7804 9270 -7676
rect 9000 -7836 9119 -7804
rect 9151 -7836 9270 -7804
rect 9000 -7964 9270 -7836
rect 9000 -7996 9119 -7964
rect 9151 -7996 9270 -7964
rect 9000 -8124 9270 -7996
rect 9000 -8156 9119 -8124
rect 9151 -8156 9270 -8124
rect 9000 -8284 9270 -8156
rect 9000 -8316 9119 -8284
rect 9151 -8316 9270 -8284
rect 9000 -8444 9270 -8316
rect 9000 -8476 9119 -8444
rect 9151 -8476 9270 -8444
rect 9000 -8604 9270 -8476
rect 9000 -8636 9119 -8604
rect 9151 -8636 9270 -8604
rect 9000 -8764 9270 -8636
rect 9000 -8796 9119 -8764
rect 9151 -8796 9270 -8764
rect 9000 -8924 9270 -8796
rect 9000 -8956 9119 -8924
rect 9151 -8956 9270 -8924
rect 9000 -9084 9270 -8956
rect 9000 -9116 9119 -9084
rect 9151 -9116 9270 -9084
rect 9000 -9230 9270 -9116
rect 12730 -5884 13000 -5770
rect 12730 -5916 12852 -5884
rect 12884 -5916 13000 -5884
rect 12730 -6044 13000 -5916
rect 12730 -6076 12852 -6044
rect 12884 -6076 13000 -6044
rect 12730 -6204 13000 -6076
rect 12730 -6236 12852 -6204
rect 12884 -6236 13000 -6204
rect 12730 -6364 13000 -6236
rect 12730 -6396 12852 -6364
rect 12884 -6396 13000 -6364
rect 12730 -6524 13000 -6396
rect 12730 -6556 12852 -6524
rect 12884 -6556 13000 -6524
rect 12730 -6684 13000 -6556
rect 12730 -6716 12852 -6684
rect 12884 -6716 13000 -6684
rect 12730 -6844 13000 -6716
rect 12730 -6876 12852 -6844
rect 12884 -6876 13000 -6844
rect 12730 -7004 13000 -6876
rect 12730 -7036 12852 -7004
rect 12884 -7036 13000 -7004
rect 12730 -7164 13000 -7036
rect 12730 -7196 12852 -7164
rect 12884 -7196 13000 -7164
rect 12730 -7324 13000 -7196
rect 12730 -7356 12852 -7324
rect 12884 -7356 13000 -7324
rect 12730 -7484 13000 -7356
rect 12730 -7516 12852 -7484
rect 12884 -7516 13000 -7484
rect 12730 -7644 13000 -7516
rect 12730 -7676 12852 -7644
rect 12884 -7676 13000 -7644
rect 12730 -7804 13000 -7676
rect 12730 -7836 12852 -7804
rect 12884 -7836 13000 -7804
rect 13200 -7795 13240 -5440
rect 13300 -7675 13340 -5340
rect 15000 -5621 19000 -5500
rect 15000 -5653 15304 -5621
rect 15336 -5653 15464 -5621
rect 15496 -5653 15624 -5621
rect 15656 -5653 15784 -5621
rect 15816 -5653 15944 -5621
rect 15976 -5653 16104 -5621
rect 16136 -5653 16264 -5621
rect 16296 -5653 16424 -5621
rect 16456 -5653 16584 -5621
rect 16616 -5653 16744 -5621
rect 16776 -5653 16904 -5621
rect 16936 -5653 17064 -5621
rect 17096 -5653 17224 -5621
rect 17256 -5653 17384 -5621
rect 17416 -5653 17544 -5621
rect 17576 -5653 17704 -5621
rect 17736 -5653 17864 -5621
rect 17896 -5653 18024 -5621
rect 18056 -5653 18184 -5621
rect 18216 -5653 18344 -5621
rect 18376 -5653 18504 -5621
rect 18536 -5653 18664 -5621
rect 18696 -5653 19000 -5621
rect 15000 -5724 19000 -5653
rect 15000 -5756 15119 -5724
rect 15151 -5756 18852 -5724
rect 18884 -5756 19000 -5724
rect 15000 -5770 19000 -5756
rect 15000 -5884 15270 -5770
rect 15000 -5916 15119 -5884
rect 15151 -5916 15270 -5884
rect 15000 -6044 15270 -5916
rect 15000 -6076 15119 -6044
rect 15151 -6076 15270 -6044
rect 15000 -6204 15270 -6076
rect 15000 -6236 15119 -6204
rect 15151 -6236 15270 -6204
rect 15000 -6364 15270 -6236
rect 15000 -6396 15119 -6364
rect 15151 -6396 15270 -6364
rect 15000 -6524 15270 -6396
rect 15000 -6556 15119 -6524
rect 15151 -6556 15270 -6524
rect 15000 -6684 15270 -6556
rect 15000 -6716 15119 -6684
rect 15151 -6716 15270 -6684
rect 15000 -6844 15270 -6716
rect 15000 -6876 15119 -6844
rect 15151 -6876 15270 -6844
rect 15000 -7004 15270 -6876
rect 15000 -7036 15119 -7004
rect 15151 -7036 15270 -7004
rect 15000 -7164 15270 -7036
rect 15000 -7196 15119 -7164
rect 15151 -7196 15270 -7164
rect 15000 -7324 15270 -7196
rect 15000 -7356 15119 -7324
rect 15151 -7356 15270 -7324
rect 15000 -7484 15270 -7356
rect 15000 -7516 15119 -7484
rect 15151 -7516 15270 -7484
rect 15000 -7644 15270 -7516
rect 15000 -7675 15119 -7644
rect 13300 -7676 15119 -7675
rect 15151 -7676 15270 -7644
rect 13300 -7715 15270 -7676
rect 13200 -7835 14585 -7795
rect 12730 -7964 13000 -7836
rect 12730 -7996 12852 -7964
rect 12884 -7996 13000 -7964
rect 12730 -8124 13000 -7996
rect 12730 -8156 12852 -8124
rect 12884 -8156 13000 -8124
rect 12730 -8284 13000 -8156
rect 12730 -8316 12852 -8284
rect 12884 -8316 13000 -8284
rect 12730 -8444 13000 -8316
rect 12730 -8476 12852 -8444
rect 12884 -8476 13000 -8444
rect 12730 -8604 13000 -8476
rect 12730 -8636 12852 -8604
rect 12884 -8636 13000 -8604
rect 12730 -8764 13000 -8636
rect 12730 -8796 12852 -8764
rect 12884 -8796 13000 -8764
rect 12730 -8924 13000 -8796
rect 12730 -8956 12852 -8924
rect 12884 -8956 13000 -8924
rect 12730 -9084 13000 -8956
rect 12730 -9116 12852 -9084
rect 12884 -9116 13000 -9084
rect 12730 -9230 13000 -9116
rect 9000 -9244 13000 -9230
rect 9000 -9276 9119 -9244
rect 9151 -9276 12852 -9244
rect 12884 -9276 13000 -9244
rect 9000 -9349 13000 -9276
rect 9000 -9381 9304 -9349
rect 9336 -9381 9464 -9349
rect 9496 -9381 9624 -9349
rect 9656 -9381 9784 -9349
rect 9816 -9381 9944 -9349
rect 9976 -9381 10104 -9349
rect 10136 -9381 10264 -9349
rect 10296 -9381 10424 -9349
rect 10456 -9381 10584 -9349
rect 10616 -9381 10744 -9349
rect 10776 -9381 10904 -9349
rect 10936 -9381 11064 -9349
rect 11096 -9381 11224 -9349
rect 11256 -9381 11384 -9349
rect 11416 -9381 11544 -9349
rect 11576 -9381 11704 -9349
rect 11736 -9381 11864 -9349
rect 11896 -9381 12024 -9349
rect 12056 -9381 12184 -9349
rect 12216 -9381 12344 -9349
rect 12376 -9381 12504 -9349
rect 12536 -9381 12664 -9349
rect 12696 -9381 13000 -9349
rect 9000 -9500 13000 -9381
rect 14545 -11120 14585 -7835
rect 15000 -7804 15270 -7715
rect 15000 -7836 15119 -7804
rect 15151 -7836 15270 -7804
rect 15000 -7964 15270 -7836
rect 15000 -7996 15119 -7964
rect 15151 -7996 15270 -7964
rect 15000 -8124 15270 -7996
rect 15000 -8156 15119 -8124
rect 15151 -8156 15270 -8124
rect 15000 -8284 15270 -8156
rect 15000 -8316 15119 -8284
rect 15151 -8316 15270 -8284
rect 15000 -8444 15270 -8316
rect 15000 -8476 15119 -8444
rect 15151 -8476 15270 -8444
rect 15000 -8604 15270 -8476
rect 15000 -8636 15119 -8604
rect 15151 -8636 15270 -8604
rect 15000 -8764 15270 -8636
rect 15000 -8796 15119 -8764
rect 15151 -8796 15270 -8764
rect 15000 -8924 15270 -8796
rect 15000 -8956 15119 -8924
rect 15151 -8956 15270 -8924
rect 15000 -9084 15270 -8956
rect 15000 -9116 15119 -9084
rect 15151 -9116 15270 -9084
rect 15000 -9230 15270 -9116
rect 18730 -5884 19000 -5770
rect 18730 -5916 18852 -5884
rect 18884 -5916 19000 -5884
rect 18730 -6044 19000 -5916
rect 18730 -6076 18852 -6044
rect 18884 -6076 19000 -6044
rect 18730 -6204 19000 -6076
rect 18730 -6236 18852 -6204
rect 18884 -6236 19000 -6204
rect 18730 -6364 19000 -6236
rect 18730 -6396 18852 -6364
rect 18884 -6396 19000 -6364
rect 18730 -6524 19000 -6396
rect 18730 -6556 18852 -6524
rect 18884 -6556 19000 -6524
rect 18730 -6684 19000 -6556
rect 18730 -6716 18852 -6684
rect 18884 -6716 19000 -6684
rect 18730 -6844 19000 -6716
rect 18730 -6876 18852 -6844
rect 18884 -6876 19000 -6844
rect 18730 -7004 19000 -6876
rect 18730 -7036 18852 -7004
rect 18884 -7036 19000 -7004
rect 18730 -7164 19000 -7036
rect 18730 -7196 18852 -7164
rect 18884 -7196 19000 -7164
rect 18730 -7324 19000 -7196
rect 18730 -7356 18852 -7324
rect 18884 -7356 19000 -7324
rect 18730 -7484 19000 -7356
rect 18730 -7516 18852 -7484
rect 18884 -7516 19000 -7484
rect 18730 -7644 19000 -7516
rect 18730 -7676 18852 -7644
rect 18884 -7676 19000 -7644
rect 18730 -7804 19000 -7676
rect 18730 -7836 18852 -7804
rect 18884 -7836 19000 -7804
rect 18730 -7964 19000 -7836
rect 18730 -7996 18852 -7964
rect 18884 -7996 19000 -7964
rect 18730 -8124 19000 -7996
rect 18730 -8156 18852 -8124
rect 18884 -8156 19000 -8124
rect 18730 -8284 19000 -8156
rect 18730 -8316 18852 -8284
rect 18884 -8316 19000 -8284
rect 18730 -8444 19000 -8316
rect 18730 -8476 18852 -8444
rect 18884 -8476 19000 -8444
rect 18730 -8604 19000 -8476
rect 18730 -8636 18852 -8604
rect 18884 -8636 19000 -8604
rect 18730 -8764 19000 -8636
rect 18730 -8796 18852 -8764
rect 18884 -8796 19000 -8764
rect 18730 -8924 19000 -8796
rect 18730 -8956 18852 -8924
rect 18884 -8956 19000 -8924
rect 18730 -9084 19000 -8956
rect 18730 -9116 18852 -9084
rect 18884 -9116 19000 -9084
rect 18730 -9230 19000 -9116
rect 15000 -9244 19000 -9230
rect 15000 -9276 15119 -9244
rect 15151 -9276 18852 -9244
rect 18884 -9276 19000 -9244
rect 15000 -9349 19000 -9276
rect 15000 -9381 15304 -9349
rect 15336 -9381 15464 -9349
rect 15496 -9381 15624 -9349
rect 15656 -9381 15784 -9349
rect 15816 -9381 15944 -9349
rect 15976 -9381 16104 -9349
rect 16136 -9381 16264 -9349
rect 16296 -9381 16424 -9349
rect 16456 -9381 16584 -9349
rect 16616 -9381 16744 -9349
rect 16776 -9381 16904 -9349
rect 16936 -9381 17064 -9349
rect 17096 -9381 17224 -9349
rect 17256 -9381 17384 -9349
rect 17416 -9381 17544 -9349
rect 17576 -9381 17704 -9349
rect 17736 -9381 17864 -9349
rect 17896 -9381 18024 -9349
rect 18056 -9381 18184 -9349
rect 18216 -9381 18344 -9349
rect 18376 -9381 18504 -9349
rect 18536 -9381 18664 -9349
rect 18696 -9381 19000 -9349
rect 15000 -9500 19000 -9381
rect 21000 -5621 25000 -5500
rect 21000 -5653 21304 -5621
rect 21336 -5653 21464 -5621
rect 21496 -5653 21624 -5621
rect 21656 -5653 21784 -5621
rect 21816 -5653 21944 -5621
rect 21976 -5653 22104 -5621
rect 22136 -5653 22264 -5621
rect 22296 -5653 22424 -5621
rect 22456 -5653 22584 -5621
rect 22616 -5653 22744 -5621
rect 22776 -5653 22904 -5621
rect 22936 -5653 23064 -5621
rect 23096 -5653 23224 -5621
rect 23256 -5653 23384 -5621
rect 23416 -5653 23544 -5621
rect 23576 -5653 23704 -5621
rect 23736 -5653 23864 -5621
rect 23896 -5653 24024 -5621
rect 24056 -5653 24184 -5621
rect 24216 -5653 24344 -5621
rect 24376 -5653 24504 -5621
rect 24536 -5653 24664 -5621
rect 24696 -5653 25000 -5621
rect 21000 -5724 25000 -5653
rect 21000 -5756 21119 -5724
rect 21151 -5756 24852 -5724
rect 24884 -5756 25000 -5724
rect 21000 -5770 25000 -5756
rect 21000 -5884 21270 -5770
rect 21000 -5916 21119 -5884
rect 21151 -5916 21270 -5884
rect 21000 -6044 21270 -5916
rect 21000 -6076 21119 -6044
rect 21151 -6076 21270 -6044
rect 21000 -6204 21270 -6076
rect 21000 -6236 21119 -6204
rect 21151 -6236 21270 -6204
rect 21000 -6364 21270 -6236
rect 21000 -6396 21119 -6364
rect 21151 -6396 21270 -6364
rect 21000 -6524 21270 -6396
rect 21000 -6556 21119 -6524
rect 21151 -6556 21270 -6524
rect 21000 -6684 21270 -6556
rect 21000 -6716 21119 -6684
rect 21151 -6716 21270 -6684
rect 21000 -6844 21270 -6716
rect 21000 -6876 21119 -6844
rect 21151 -6876 21270 -6844
rect 21000 -7004 21270 -6876
rect 21000 -7036 21119 -7004
rect 21151 -7036 21270 -7004
rect 21000 -7164 21270 -7036
rect 21000 -7196 21119 -7164
rect 21151 -7196 21270 -7164
rect 21000 -7324 21270 -7196
rect 21000 -7356 21119 -7324
rect 21151 -7356 21270 -7324
rect 21000 -7484 21270 -7356
rect 21000 -7516 21119 -7484
rect 21151 -7516 21270 -7484
rect 21000 -7644 21270 -7516
rect 21000 -7676 21119 -7644
rect 21151 -7676 21270 -7644
rect 21000 -7804 21270 -7676
rect 21000 -7836 21119 -7804
rect 21151 -7836 21270 -7804
rect 21000 -7964 21270 -7836
rect 21000 -7996 21119 -7964
rect 21151 -7996 21270 -7964
rect 21000 -8124 21270 -7996
rect 21000 -8156 21119 -8124
rect 21151 -8156 21270 -8124
rect 21000 -8284 21270 -8156
rect 21000 -8316 21119 -8284
rect 21151 -8316 21270 -8284
rect 21000 -8444 21270 -8316
rect 21000 -8476 21119 -8444
rect 21151 -8476 21270 -8444
rect 21000 -8604 21270 -8476
rect 21000 -8636 21119 -8604
rect 21151 -8636 21270 -8604
rect 21000 -8764 21270 -8636
rect 21000 -8796 21119 -8764
rect 21151 -8796 21270 -8764
rect 21000 -8924 21270 -8796
rect 21000 -8956 21119 -8924
rect 21151 -8956 21270 -8924
rect 21000 -9084 21270 -8956
rect 21000 -9116 21119 -9084
rect 21151 -9116 21270 -9084
rect 21000 -9230 21270 -9116
rect 24730 -5884 25000 -5770
rect 24730 -5916 24852 -5884
rect 24884 -5916 25000 -5884
rect 24730 -6044 25000 -5916
rect 24730 -6076 24852 -6044
rect 24884 -6076 25000 -6044
rect 24730 -6204 25000 -6076
rect 24730 -6236 24852 -6204
rect 24884 -6236 25000 -6204
rect 24730 -6364 25000 -6236
rect 24730 -6396 24852 -6364
rect 24884 -6396 25000 -6364
rect 24730 -6524 25000 -6396
rect 24730 -6556 24852 -6524
rect 24884 -6556 25000 -6524
rect 24730 -6684 25000 -6556
rect 24730 -6716 24852 -6684
rect 24884 -6716 25000 -6684
rect 24730 -6844 25000 -6716
rect 24730 -6876 24852 -6844
rect 24884 -6876 25000 -6844
rect 24730 -7004 25000 -6876
rect 24730 -7036 24852 -7004
rect 24884 -7036 25000 -7004
rect 24730 -7164 25000 -7036
rect 24730 -7196 24852 -7164
rect 24884 -7196 25000 -7164
rect 24730 -7324 25000 -7196
rect 24730 -7356 24852 -7324
rect 24884 -7356 25000 -7324
rect 24730 -7484 25000 -7356
rect 24730 -7516 24852 -7484
rect 24884 -7516 25000 -7484
rect 24730 -7644 25000 -7516
rect 24730 -7676 24852 -7644
rect 24884 -7676 25000 -7644
rect 24730 -7804 25000 -7676
rect 24730 -7836 24852 -7804
rect 24884 -7836 25000 -7804
rect 24730 -7964 25000 -7836
rect 24730 -7996 24852 -7964
rect 24884 -7996 25000 -7964
rect 24730 -8124 25000 -7996
rect 24730 -8156 24852 -8124
rect 24884 -8156 25000 -8124
rect 24730 -8284 25000 -8156
rect 24730 -8316 24852 -8284
rect 24884 -8316 25000 -8284
rect 24730 -8444 25000 -8316
rect 24730 -8476 24852 -8444
rect 24884 -8476 25000 -8444
rect 24730 -8604 25000 -8476
rect 24730 -8636 24852 -8604
rect 24884 -8636 25000 -8604
rect 24730 -8764 25000 -8636
rect 24730 -8796 24852 -8764
rect 24884 -8796 25000 -8764
rect 24730 -8924 25000 -8796
rect 24730 -8956 24852 -8924
rect 24884 -8956 25000 -8924
rect 24730 -9084 25000 -8956
rect 24730 -9116 24852 -9084
rect 24884 -9116 25000 -9084
rect 24730 -9230 25000 -9116
rect 21000 -9244 25000 -9230
rect 21000 -9276 21119 -9244
rect 21151 -9276 24852 -9244
rect 24884 -9276 25000 -9244
rect 21000 -9349 25000 -9276
rect 21000 -9381 21304 -9349
rect 21336 -9381 21464 -9349
rect 21496 -9381 21624 -9349
rect 21656 -9381 21784 -9349
rect 21816 -9381 21944 -9349
rect 21976 -9381 22104 -9349
rect 22136 -9381 22264 -9349
rect 22296 -9381 22424 -9349
rect 22456 -9381 22584 -9349
rect 22616 -9381 22744 -9349
rect 22776 -9381 22904 -9349
rect 22936 -9381 23064 -9349
rect 23096 -9381 23224 -9349
rect 23256 -9381 23384 -9349
rect 23416 -9381 23544 -9349
rect 23576 -9381 23704 -9349
rect 23736 -9381 23864 -9349
rect 23896 -9381 24024 -9349
rect 24056 -9381 24184 -9349
rect 24216 -9381 24344 -9349
rect 24376 -9381 24504 -9349
rect 24536 -9381 24664 -9349
rect 24696 -9381 25000 -9349
rect 21000 -9500 25000 -9381
rect 14545 -11160 21375 -11120
rect 8300 -11360 14150 -11330
rect 9000 -11621 13000 -11500
rect 9000 -11653 9304 -11621
rect 9336 -11653 9464 -11621
rect 9496 -11653 9624 -11621
rect 9656 -11653 9784 -11621
rect 9816 -11653 9944 -11621
rect 9976 -11653 10104 -11621
rect 10136 -11653 10264 -11621
rect 10296 -11653 10424 -11621
rect 10456 -11653 10584 -11621
rect 10616 -11653 10744 -11621
rect 10776 -11653 10904 -11621
rect 10936 -11653 11064 -11621
rect 11096 -11653 11224 -11621
rect 11256 -11653 11384 -11621
rect 11416 -11653 11544 -11621
rect 11576 -11653 11704 -11621
rect 11736 -11653 11864 -11621
rect 11896 -11653 12024 -11621
rect 12056 -11653 12184 -11621
rect 12216 -11653 12344 -11621
rect 12376 -11653 12504 -11621
rect 12536 -11653 12664 -11621
rect 12696 -11653 13000 -11621
rect 9000 -11724 13000 -11653
rect 9000 -11756 9119 -11724
rect 9151 -11756 12852 -11724
rect 12884 -11756 13000 -11724
rect 9000 -11770 13000 -11756
rect 9000 -11884 9270 -11770
rect 9000 -11916 9119 -11884
rect 9151 -11916 9270 -11884
rect 9000 -12044 9270 -11916
rect 9000 -12076 9119 -12044
rect 9151 -12076 9270 -12044
rect 9000 -12204 9270 -12076
rect 9000 -12236 9119 -12204
rect 9151 -12236 9270 -12204
rect 9000 -12364 9270 -12236
rect 9000 -12396 9119 -12364
rect 9151 -12396 9270 -12364
rect 9000 -12524 9270 -12396
rect 9000 -12556 9119 -12524
rect 9151 -12556 9270 -12524
rect 9000 -12684 9270 -12556
rect 9000 -12716 9119 -12684
rect 9151 -12716 9270 -12684
rect 9000 -12844 9270 -12716
rect 9000 -12875 9119 -12844
rect 8230 -12876 9119 -12875
rect 9151 -12876 9270 -12844
rect 6730 -13004 7000 -12900
rect 8230 -12905 9270 -12876
rect 6730 -13036 6852 -13004
rect 6884 -13036 7000 -13004
rect 6730 -13164 7000 -13036
rect 6730 -13196 6852 -13164
rect 6884 -13196 7000 -13164
rect 6730 -13324 7000 -13196
rect 6730 -13356 6852 -13324
rect 6884 -13356 7000 -13324
rect 6730 -13484 7000 -13356
rect 6730 -13516 6852 -13484
rect 6884 -13516 7000 -13484
rect 6730 -13644 7000 -13516
rect 6730 -13676 6852 -13644
rect 6884 -13676 7000 -13644
rect 6730 -13804 7000 -13676
rect 6730 -13836 6852 -13804
rect 6884 -13836 7000 -13804
rect 6730 -13964 7000 -13836
rect 6730 -13996 6852 -13964
rect 6884 -13996 7000 -13964
rect 6730 -14124 7000 -13996
rect 6730 -14156 6852 -14124
rect 6884 -14156 7000 -14124
rect 6730 -14284 7000 -14156
rect 6730 -14316 6852 -14284
rect 6884 -14316 7000 -14284
rect 6730 -14444 7000 -14316
rect 6730 -14476 6852 -14444
rect 6884 -14476 7000 -14444
rect 6730 -14604 7000 -14476
rect 6730 -14636 6852 -14604
rect 6884 -14636 7000 -14604
rect 6730 -14764 7000 -14636
rect 6730 -14796 6852 -14764
rect 6884 -14796 7000 -14764
rect 6730 -14924 7000 -14796
rect 6730 -14956 6852 -14924
rect 6884 -14956 7000 -14924
rect 6730 -15084 7000 -14956
rect 6730 -15116 6852 -15084
rect 6884 -15116 7000 -15084
rect 6730 -15230 7000 -15116
rect 3000 -15244 7000 -15230
rect 3000 -15276 3119 -15244
rect 3151 -15276 6852 -15244
rect 6884 -15276 7000 -15244
rect 3000 -15349 7000 -15276
rect 3000 -15381 3304 -15349
rect 3336 -15381 3464 -15349
rect 3496 -15381 3624 -15349
rect 3656 -15381 3784 -15349
rect 3816 -15381 3944 -15349
rect 3976 -15381 4104 -15349
rect 4136 -15381 4264 -15349
rect 4296 -15381 4424 -15349
rect 4456 -15381 4584 -15349
rect 4616 -15381 4744 -15349
rect 4776 -15381 4904 -15349
rect 4936 -15381 5064 -15349
rect 5096 -15381 5224 -15349
rect 5256 -15381 5384 -15349
rect 5416 -15381 5544 -15349
rect 5576 -15381 5704 -15349
rect 5736 -15381 5864 -15349
rect 5896 -15381 6024 -15349
rect 6056 -15381 6184 -15349
rect 6216 -15381 6344 -15349
rect 6376 -15381 6504 -15349
rect 6536 -15381 6664 -15349
rect 6696 -15381 7000 -15349
rect 3000 -15500 7000 -15381
rect 9000 -13004 9270 -12905
rect 9000 -13036 9119 -13004
rect 9151 -13036 9270 -13004
rect 9000 -13164 9270 -13036
rect 9000 -13196 9119 -13164
rect 9151 -13196 9270 -13164
rect 9000 -13324 9270 -13196
rect 9000 -13356 9119 -13324
rect 9151 -13356 9270 -13324
rect 9000 -13484 9270 -13356
rect 9000 -13516 9119 -13484
rect 9151 -13516 9270 -13484
rect 9000 -13644 9270 -13516
rect 9000 -13676 9119 -13644
rect 9151 -13676 9270 -13644
rect 9000 -13804 9270 -13676
rect 9000 -13836 9119 -13804
rect 9151 -13836 9270 -13804
rect 9000 -13964 9270 -13836
rect 9000 -13996 9119 -13964
rect 9151 -13996 9270 -13964
rect 9000 -14124 9270 -13996
rect 9000 -14156 9119 -14124
rect 9151 -14156 9270 -14124
rect 9000 -14284 9270 -14156
rect 9000 -14316 9119 -14284
rect 9151 -14316 9270 -14284
rect 9000 -14444 9270 -14316
rect 9000 -14476 9119 -14444
rect 9151 -14476 9270 -14444
rect 9000 -14604 9270 -14476
rect 9000 -14636 9119 -14604
rect 9151 -14636 9270 -14604
rect 9000 -14764 9270 -14636
rect 9000 -14796 9119 -14764
rect 9151 -14796 9270 -14764
rect 9000 -14924 9270 -14796
rect 9000 -14956 9119 -14924
rect 9151 -14956 9270 -14924
rect 9000 -15084 9270 -14956
rect 9000 -15116 9119 -15084
rect 9151 -15116 9270 -15084
rect 9000 -15230 9270 -15116
rect 12730 -11884 13000 -11770
rect 12730 -11916 12852 -11884
rect 12884 -11916 13000 -11884
rect 12730 -12044 13000 -11916
rect 12730 -12076 12852 -12044
rect 12884 -12076 13000 -12044
rect 12730 -12204 13000 -12076
rect 12730 -12236 12852 -12204
rect 12884 -12236 13000 -12204
rect 12730 -12364 13000 -12236
rect 12730 -12396 12852 -12364
rect 12884 -12396 13000 -12364
rect 12730 -12524 13000 -12396
rect 12730 -12556 12852 -12524
rect 12884 -12556 13000 -12524
rect 12730 -12684 13000 -12556
rect 12730 -12716 12852 -12684
rect 12884 -12716 13000 -12684
rect 12730 -12844 13000 -12716
rect 12730 -12876 12852 -12844
rect 12884 -12876 13000 -12844
rect 12730 -13004 13000 -12876
rect 14120 -12870 14150 -11360
rect 21335 -11500 21375 -11160
rect 15000 -11621 19000 -11500
rect 15000 -11653 15304 -11621
rect 15336 -11653 15464 -11621
rect 15496 -11653 15624 -11621
rect 15656 -11653 15784 -11621
rect 15816 -11653 15944 -11621
rect 15976 -11653 16104 -11621
rect 16136 -11653 16264 -11621
rect 16296 -11653 16424 -11621
rect 16456 -11653 16584 -11621
rect 16616 -11653 16744 -11621
rect 16776 -11653 16904 -11621
rect 16936 -11653 17064 -11621
rect 17096 -11653 17224 -11621
rect 17256 -11653 17384 -11621
rect 17416 -11653 17544 -11621
rect 17576 -11653 17704 -11621
rect 17736 -11653 17864 -11621
rect 17896 -11653 18024 -11621
rect 18056 -11653 18184 -11621
rect 18216 -11653 18344 -11621
rect 18376 -11653 18504 -11621
rect 18536 -11653 18664 -11621
rect 18696 -11653 19000 -11621
rect 15000 -11724 19000 -11653
rect 15000 -11756 15119 -11724
rect 15151 -11756 18852 -11724
rect 18884 -11756 19000 -11724
rect 15000 -11770 19000 -11756
rect 15000 -11884 15270 -11770
rect 15000 -11916 15119 -11884
rect 15151 -11916 15270 -11884
rect 15000 -12044 15270 -11916
rect 15000 -12076 15119 -12044
rect 15151 -12076 15270 -12044
rect 15000 -12204 15270 -12076
rect 15000 -12236 15119 -12204
rect 15151 -12236 15270 -12204
rect 15000 -12364 15270 -12236
rect 15000 -12396 15119 -12364
rect 15151 -12396 15270 -12364
rect 15000 -12524 15270 -12396
rect 15000 -12556 15119 -12524
rect 15151 -12556 15270 -12524
rect 15000 -12684 15270 -12556
rect 15000 -12716 15119 -12684
rect 15151 -12716 15270 -12684
rect 15000 -12844 15270 -12716
rect 15000 -12870 15119 -12844
rect 14120 -12876 15119 -12870
rect 15151 -12876 15270 -12844
rect 14120 -12900 15270 -12876
rect 12730 -13036 12852 -13004
rect 12884 -13036 13000 -13004
rect 12730 -13164 13000 -13036
rect 12730 -13196 12852 -13164
rect 12884 -13196 13000 -13164
rect 12730 -13324 13000 -13196
rect 12730 -13356 12852 -13324
rect 12884 -13356 13000 -13324
rect 12730 -13484 13000 -13356
rect 12730 -13516 12852 -13484
rect 12884 -13516 13000 -13484
rect 12730 -13644 13000 -13516
rect 12730 -13676 12852 -13644
rect 12884 -13676 13000 -13644
rect 12730 -13804 13000 -13676
rect 12730 -13836 12852 -13804
rect 12884 -13836 13000 -13804
rect 12730 -13964 13000 -13836
rect 12730 -13996 12852 -13964
rect 12884 -13996 13000 -13964
rect 12730 -14124 13000 -13996
rect 12730 -14156 12852 -14124
rect 12884 -14156 13000 -14124
rect 12730 -14284 13000 -14156
rect 12730 -14316 12852 -14284
rect 12884 -14316 13000 -14284
rect 12730 -14444 13000 -14316
rect 12730 -14476 12852 -14444
rect 12884 -14476 13000 -14444
rect 12730 -14604 13000 -14476
rect 12730 -14636 12852 -14604
rect 12884 -14636 13000 -14604
rect 12730 -14764 13000 -14636
rect 12730 -14796 12852 -14764
rect 12884 -14796 13000 -14764
rect 12730 -14924 13000 -14796
rect 12730 -14956 12852 -14924
rect 12884 -14956 13000 -14924
rect 12730 -15084 13000 -14956
rect 12730 -15116 12852 -15084
rect 12884 -15116 13000 -15084
rect 12730 -15230 13000 -15116
rect 9000 -15244 13000 -15230
rect 9000 -15276 9119 -15244
rect 9151 -15276 12852 -15244
rect 12884 -15276 13000 -15244
rect 9000 -15349 13000 -15276
rect 9000 -15381 9304 -15349
rect 9336 -15381 9464 -15349
rect 9496 -15381 9624 -15349
rect 9656 -15381 9784 -15349
rect 9816 -15381 9944 -15349
rect 9976 -15381 10104 -15349
rect 10136 -15381 10264 -15349
rect 10296 -15381 10424 -15349
rect 10456 -15381 10584 -15349
rect 10616 -15381 10744 -15349
rect 10776 -15381 10904 -15349
rect 10936 -15381 11064 -15349
rect 11096 -15381 11224 -15349
rect 11256 -15381 11384 -15349
rect 11416 -15381 11544 -15349
rect 11576 -15381 11704 -15349
rect 11736 -15381 11864 -15349
rect 11896 -15381 12024 -15349
rect 12056 -15381 12184 -15349
rect 12216 -15381 12344 -15349
rect 12376 -15381 12504 -15349
rect 12536 -15381 12664 -15349
rect 12696 -15381 13000 -15349
rect 9000 -15500 13000 -15381
rect 15000 -13004 15270 -12900
rect 15000 -13036 15119 -13004
rect 15151 -13036 15270 -13004
rect 15000 -13164 15270 -13036
rect 15000 -13196 15119 -13164
rect 15151 -13196 15270 -13164
rect 15000 -13324 15270 -13196
rect 15000 -13356 15119 -13324
rect 15151 -13356 15270 -13324
rect 15000 -13484 15270 -13356
rect 15000 -13516 15119 -13484
rect 15151 -13516 15270 -13484
rect 15000 -13644 15270 -13516
rect 15000 -13676 15119 -13644
rect 15151 -13676 15270 -13644
rect 15000 -13804 15270 -13676
rect 15000 -13836 15119 -13804
rect 15151 -13836 15270 -13804
rect 15000 -13964 15270 -13836
rect 15000 -13996 15119 -13964
rect 15151 -13996 15270 -13964
rect 15000 -14124 15270 -13996
rect 15000 -14156 15119 -14124
rect 15151 -14156 15270 -14124
rect 15000 -14284 15270 -14156
rect 15000 -14316 15119 -14284
rect 15151 -14316 15270 -14284
rect 15000 -14444 15270 -14316
rect 15000 -14476 15119 -14444
rect 15151 -14476 15270 -14444
rect 15000 -14604 15270 -14476
rect 15000 -14636 15119 -14604
rect 15151 -14636 15270 -14604
rect 15000 -14764 15270 -14636
rect 15000 -14796 15119 -14764
rect 15151 -14796 15270 -14764
rect 15000 -14924 15270 -14796
rect 15000 -14956 15119 -14924
rect 15151 -14956 15270 -14924
rect 15000 -15084 15270 -14956
rect 15000 -15116 15119 -15084
rect 15151 -15116 15270 -15084
rect 15000 -15230 15270 -15116
rect 18730 -11884 19000 -11770
rect 18730 -11916 18852 -11884
rect 18884 -11916 19000 -11884
rect 18730 -12044 19000 -11916
rect 18730 -12076 18852 -12044
rect 18884 -12076 19000 -12044
rect 18730 -12204 19000 -12076
rect 18730 -12236 18852 -12204
rect 18884 -12236 19000 -12204
rect 18730 -12364 19000 -12236
rect 18730 -12396 18852 -12364
rect 18884 -12396 19000 -12364
rect 18730 -12524 19000 -12396
rect 18730 -12556 18852 -12524
rect 18884 -12556 19000 -12524
rect 18730 -12684 19000 -12556
rect 18730 -12716 18852 -12684
rect 18884 -12716 19000 -12684
rect 18730 -12844 19000 -12716
rect 18730 -12876 18852 -12844
rect 18884 -12876 19000 -12844
rect 18730 -13004 19000 -12876
rect 18730 -13036 18852 -13004
rect 18884 -13036 19000 -13004
rect 18730 -13164 19000 -13036
rect 18730 -13196 18852 -13164
rect 18884 -13196 19000 -13164
rect 18730 -13324 19000 -13196
rect 18730 -13356 18852 -13324
rect 18884 -13356 19000 -13324
rect 18730 -13484 19000 -13356
rect 18730 -13516 18852 -13484
rect 18884 -13516 19000 -13484
rect 18730 -13644 19000 -13516
rect 18730 -13676 18852 -13644
rect 18884 -13676 19000 -13644
rect 18730 -13804 19000 -13676
rect 18730 -13836 18852 -13804
rect 18884 -13836 19000 -13804
rect 18730 -13964 19000 -13836
rect 18730 -13996 18852 -13964
rect 18884 -13996 19000 -13964
rect 18730 -14124 19000 -13996
rect 18730 -14156 18852 -14124
rect 18884 -14156 19000 -14124
rect 18730 -14284 19000 -14156
rect 18730 -14316 18852 -14284
rect 18884 -14316 19000 -14284
rect 18730 -14444 19000 -14316
rect 18730 -14476 18852 -14444
rect 18884 -14476 19000 -14444
rect 18730 -14604 19000 -14476
rect 18730 -14636 18852 -14604
rect 18884 -14636 19000 -14604
rect 18730 -14764 19000 -14636
rect 18730 -14796 18852 -14764
rect 18884 -14796 19000 -14764
rect 18730 -14924 19000 -14796
rect 18730 -14956 18852 -14924
rect 18884 -14956 19000 -14924
rect 18730 -15084 19000 -14956
rect 18730 -15116 18852 -15084
rect 18884 -15116 19000 -15084
rect 18730 -15230 19000 -15116
rect 15000 -15244 19000 -15230
rect 15000 -15276 15119 -15244
rect 15151 -15276 18852 -15244
rect 18884 -15276 19000 -15244
rect 15000 -15349 19000 -15276
rect 15000 -15381 15304 -15349
rect 15336 -15381 15464 -15349
rect 15496 -15381 15624 -15349
rect 15656 -15381 15784 -15349
rect 15816 -15381 15944 -15349
rect 15976 -15381 16104 -15349
rect 16136 -15381 16264 -15349
rect 16296 -15381 16424 -15349
rect 16456 -15381 16584 -15349
rect 16616 -15381 16744 -15349
rect 16776 -15381 16904 -15349
rect 16936 -15381 17064 -15349
rect 17096 -15381 17224 -15349
rect 17256 -15381 17384 -15349
rect 17416 -15381 17544 -15349
rect 17576 -15381 17704 -15349
rect 17736 -15381 17864 -15349
rect 17896 -15381 18024 -15349
rect 18056 -15381 18184 -15349
rect 18216 -15381 18344 -15349
rect 18376 -15381 18504 -15349
rect 18536 -15381 18664 -15349
rect 18696 -15381 19000 -15349
rect 15000 -15500 19000 -15381
rect 21000 -11621 25000 -11500
rect 21000 -11653 21304 -11621
rect 21336 -11653 21464 -11621
rect 21496 -11653 21624 -11621
rect 21656 -11653 21784 -11621
rect 21816 -11653 21944 -11621
rect 21976 -11653 22104 -11621
rect 22136 -11653 22264 -11621
rect 22296 -11653 22424 -11621
rect 22456 -11653 22584 -11621
rect 22616 -11653 22744 -11621
rect 22776 -11653 22904 -11621
rect 22936 -11653 23064 -11621
rect 23096 -11653 23224 -11621
rect 23256 -11653 23384 -11621
rect 23416 -11653 23544 -11621
rect 23576 -11653 23704 -11621
rect 23736 -11653 23864 -11621
rect 23896 -11653 24024 -11621
rect 24056 -11653 24184 -11621
rect 24216 -11653 24344 -11621
rect 24376 -11653 24504 -11621
rect 24536 -11653 24664 -11621
rect 24696 -11653 25000 -11621
rect 21000 -11724 25000 -11653
rect 21000 -11756 21119 -11724
rect 21151 -11756 24852 -11724
rect 24884 -11756 25000 -11724
rect 21000 -11770 25000 -11756
rect 21000 -11884 21270 -11770
rect 21000 -11916 21119 -11884
rect 21151 -11916 21270 -11884
rect 21000 -12044 21270 -11916
rect 21000 -12076 21119 -12044
rect 21151 -12076 21270 -12044
rect 21000 -12204 21270 -12076
rect 21000 -12236 21119 -12204
rect 21151 -12236 21270 -12204
rect 21000 -12364 21270 -12236
rect 21000 -12396 21119 -12364
rect 21151 -12396 21270 -12364
rect 21000 -12524 21270 -12396
rect 21000 -12556 21119 -12524
rect 21151 -12556 21270 -12524
rect 21000 -12684 21270 -12556
rect 21000 -12716 21119 -12684
rect 21151 -12716 21270 -12684
rect 21000 -12844 21270 -12716
rect 21000 -12876 21119 -12844
rect 21151 -12876 21270 -12844
rect 21000 -13004 21270 -12876
rect 21000 -13036 21119 -13004
rect 21151 -13036 21270 -13004
rect 21000 -13164 21270 -13036
rect 21000 -13196 21119 -13164
rect 21151 -13196 21270 -13164
rect 21000 -13324 21270 -13196
rect 21000 -13356 21119 -13324
rect 21151 -13356 21270 -13324
rect 21000 -13484 21270 -13356
rect 21000 -13516 21119 -13484
rect 21151 -13516 21270 -13484
rect 21000 -13644 21270 -13516
rect 21000 -13676 21119 -13644
rect 21151 -13676 21270 -13644
rect 21000 -13804 21270 -13676
rect 21000 -13836 21119 -13804
rect 21151 -13836 21270 -13804
rect 21000 -13964 21270 -13836
rect 21000 -13996 21119 -13964
rect 21151 -13996 21270 -13964
rect 21000 -14124 21270 -13996
rect 21000 -14156 21119 -14124
rect 21151 -14156 21270 -14124
rect 21000 -14284 21270 -14156
rect 21000 -14316 21119 -14284
rect 21151 -14316 21270 -14284
rect 21000 -14444 21270 -14316
rect 21000 -14476 21119 -14444
rect 21151 -14476 21270 -14444
rect 21000 -14604 21270 -14476
rect 21000 -14636 21119 -14604
rect 21151 -14636 21270 -14604
rect 21000 -14764 21270 -14636
rect 21000 -14796 21119 -14764
rect 21151 -14796 21270 -14764
rect 21000 -14924 21270 -14796
rect 21000 -14956 21119 -14924
rect 21151 -14956 21270 -14924
rect 21000 -15084 21270 -14956
rect 21000 -15116 21119 -15084
rect 21151 -15116 21270 -15084
rect 21000 -15230 21270 -15116
rect 24730 -11884 25000 -11770
rect 24730 -11916 24852 -11884
rect 24884 -11916 25000 -11884
rect 24730 -12044 25000 -11916
rect 24730 -12076 24852 -12044
rect 24884 -12076 25000 -12044
rect 24730 -12204 25000 -12076
rect 24730 -12236 24852 -12204
rect 24884 -12236 25000 -12204
rect 24730 -12364 25000 -12236
rect 24730 -12396 24852 -12364
rect 24884 -12396 25000 -12364
rect 24730 -12524 25000 -12396
rect 24730 -12556 24852 -12524
rect 24884 -12556 25000 -12524
rect 24730 -12684 25000 -12556
rect 24730 -12716 24852 -12684
rect 24884 -12716 25000 -12684
rect 24730 -12844 25000 -12716
rect 24730 -12876 24852 -12844
rect 24884 -12876 25000 -12844
rect 24730 -13004 25000 -12876
rect 24730 -13036 24852 -13004
rect 24884 -13036 25000 -13004
rect 24730 -13164 25000 -13036
rect 24730 -13196 24852 -13164
rect 24884 -13196 25000 -13164
rect 24730 -13324 25000 -13196
rect 24730 -13356 24852 -13324
rect 24884 -13356 25000 -13324
rect 24730 -13484 25000 -13356
rect 24730 -13516 24852 -13484
rect 24884 -13516 25000 -13484
rect 24730 -13644 25000 -13516
rect 24730 -13676 24852 -13644
rect 24884 -13676 25000 -13644
rect 24730 -13804 25000 -13676
rect 24730 -13836 24852 -13804
rect 24884 -13836 25000 -13804
rect 24730 -13964 25000 -13836
rect 24730 -13996 24852 -13964
rect 24884 -13996 25000 -13964
rect 24730 -14124 25000 -13996
rect 24730 -14156 24852 -14124
rect 24884 -14156 25000 -14124
rect 24730 -14284 25000 -14156
rect 24730 -14316 24852 -14284
rect 24884 -14316 25000 -14284
rect 24730 -14444 25000 -14316
rect 24730 -14476 24852 -14444
rect 24884 -14476 25000 -14444
rect 24730 -14604 25000 -14476
rect 24730 -14636 24852 -14604
rect 24884 -14636 25000 -14604
rect 24730 -14764 25000 -14636
rect 24730 -14796 24852 -14764
rect 24884 -14796 25000 -14764
rect 24730 -14924 25000 -14796
rect 24730 -14956 24852 -14924
rect 24884 -14956 25000 -14924
rect 24730 -15084 25000 -14956
rect 24730 -15116 24852 -15084
rect 24884 -15116 25000 -15084
rect 24730 -15230 25000 -15116
rect 21000 -15244 25000 -15230
rect 21000 -15276 21119 -15244
rect 21151 -15276 24852 -15244
rect 24884 -15276 25000 -15244
rect 21000 -15349 25000 -15276
rect 21000 -15381 21304 -15349
rect 21336 -15381 21464 -15349
rect 21496 -15381 21624 -15349
rect 21656 -15381 21784 -15349
rect 21816 -15381 21944 -15349
rect 21976 -15381 22104 -15349
rect 22136 -15381 22264 -15349
rect 22296 -15381 22424 -15349
rect 22456 -15381 22584 -15349
rect 22616 -15381 22744 -15349
rect 22776 -15381 22904 -15349
rect 22936 -15381 23064 -15349
rect 23096 -15381 23224 -15349
rect 23256 -15381 23384 -15349
rect 23416 -15381 23544 -15349
rect 23576 -15381 23704 -15349
rect 23736 -15381 23864 -15349
rect 23896 -15381 24024 -15349
rect 24056 -15381 24184 -15349
rect 24216 -15381 24344 -15349
rect 24376 -15381 24504 -15349
rect 24536 -15381 24664 -15349
rect 24696 -15381 25000 -15349
rect 21000 -15500 25000 -15381
<< via3 >>
rect 3304 9379 3336 9381
rect 3304 9351 3306 9379
rect 3306 9351 3334 9379
rect 3334 9351 3336 9379
rect 3304 9349 3336 9351
rect 3464 9379 3496 9381
rect 3464 9351 3466 9379
rect 3466 9351 3494 9379
rect 3494 9351 3496 9379
rect 3464 9349 3496 9351
rect 3624 9379 3656 9381
rect 3624 9351 3626 9379
rect 3626 9351 3654 9379
rect 3654 9351 3656 9379
rect 3624 9349 3656 9351
rect 3784 9379 3816 9381
rect 3784 9351 3786 9379
rect 3786 9351 3814 9379
rect 3814 9351 3816 9379
rect 3784 9349 3816 9351
rect 3944 9379 3976 9381
rect 3944 9351 3946 9379
rect 3946 9351 3974 9379
rect 3974 9351 3976 9379
rect 3944 9349 3976 9351
rect 4104 9379 4136 9381
rect 4104 9351 4106 9379
rect 4106 9351 4134 9379
rect 4134 9351 4136 9379
rect 4104 9349 4136 9351
rect 4264 9379 4296 9381
rect 4264 9351 4266 9379
rect 4266 9351 4294 9379
rect 4294 9351 4296 9379
rect 4264 9349 4296 9351
rect 4424 9379 4456 9381
rect 4424 9351 4426 9379
rect 4426 9351 4454 9379
rect 4454 9351 4456 9379
rect 4424 9349 4456 9351
rect 4584 9379 4616 9381
rect 4584 9351 4586 9379
rect 4586 9351 4614 9379
rect 4614 9351 4616 9379
rect 4584 9349 4616 9351
rect 4744 9379 4776 9381
rect 4744 9351 4746 9379
rect 4746 9351 4774 9379
rect 4774 9351 4776 9379
rect 4744 9349 4776 9351
rect 4904 9379 4936 9381
rect 4904 9351 4906 9379
rect 4906 9351 4934 9379
rect 4934 9351 4936 9379
rect 4904 9349 4936 9351
rect 5064 9379 5096 9381
rect 5064 9351 5066 9379
rect 5066 9351 5094 9379
rect 5094 9351 5096 9379
rect 5064 9349 5096 9351
rect 5224 9379 5256 9381
rect 5224 9351 5226 9379
rect 5226 9351 5254 9379
rect 5254 9351 5256 9379
rect 5224 9349 5256 9351
rect 5384 9379 5416 9381
rect 5384 9351 5386 9379
rect 5386 9351 5414 9379
rect 5414 9351 5416 9379
rect 5384 9349 5416 9351
rect 5544 9379 5576 9381
rect 5544 9351 5546 9379
rect 5546 9351 5574 9379
rect 5574 9351 5576 9379
rect 5544 9349 5576 9351
rect 5704 9379 5736 9381
rect 5704 9351 5706 9379
rect 5706 9351 5734 9379
rect 5734 9351 5736 9379
rect 5704 9349 5736 9351
rect 5864 9379 5896 9381
rect 5864 9351 5866 9379
rect 5866 9351 5894 9379
rect 5894 9351 5896 9379
rect 5864 9349 5896 9351
rect 6024 9379 6056 9381
rect 6024 9351 6026 9379
rect 6026 9351 6054 9379
rect 6054 9351 6056 9379
rect 6024 9349 6056 9351
rect 6184 9379 6216 9381
rect 6184 9351 6186 9379
rect 6186 9351 6214 9379
rect 6214 9351 6216 9379
rect 6184 9349 6216 9351
rect 6344 9379 6376 9381
rect 6344 9351 6346 9379
rect 6346 9351 6374 9379
rect 6374 9351 6376 9379
rect 6344 9349 6376 9351
rect 6504 9379 6536 9381
rect 6504 9351 6506 9379
rect 6506 9351 6534 9379
rect 6534 9351 6536 9379
rect 6504 9349 6536 9351
rect 6664 9379 6696 9381
rect 6664 9351 6666 9379
rect 6666 9351 6694 9379
rect 6694 9351 6696 9379
rect 6664 9349 6696 9351
rect 3116 9274 3148 9276
rect 3116 9246 3118 9274
rect 3118 9246 3146 9274
rect 3146 9246 3148 9274
rect 3116 9244 3148 9246
rect 6849 9274 6881 9276
rect 6849 9246 6851 9274
rect 6851 9246 6879 9274
rect 6879 9246 6881 9274
rect 6849 9244 6881 9246
rect 3116 9114 3148 9116
rect 3116 9086 3118 9114
rect 3118 9086 3146 9114
rect 3146 9086 3148 9114
rect 3116 9084 3148 9086
rect 3116 8954 3148 8956
rect 3116 8926 3118 8954
rect 3118 8926 3146 8954
rect 3146 8926 3148 8954
rect 3116 8924 3148 8926
rect 3116 8794 3148 8796
rect 3116 8766 3118 8794
rect 3118 8766 3146 8794
rect 3146 8766 3148 8794
rect 3116 8764 3148 8766
rect 3116 8634 3148 8636
rect 3116 8606 3118 8634
rect 3118 8606 3146 8634
rect 3146 8606 3148 8634
rect 3116 8604 3148 8606
rect 3116 8474 3148 8476
rect 3116 8446 3118 8474
rect 3118 8446 3146 8474
rect 3146 8446 3148 8474
rect 3116 8444 3148 8446
rect 3116 8314 3148 8316
rect 3116 8286 3118 8314
rect 3118 8286 3146 8314
rect 3146 8286 3148 8314
rect 3116 8284 3148 8286
rect 3116 8154 3148 8156
rect 3116 8126 3118 8154
rect 3118 8126 3146 8154
rect 3146 8126 3148 8154
rect 3116 8124 3148 8126
rect 3116 7994 3148 7996
rect 3116 7966 3118 7994
rect 3118 7966 3146 7994
rect 3146 7966 3148 7994
rect 3116 7964 3148 7966
rect 3116 7834 3148 7836
rect 3116 7806 3118 7834
rect 3118 7806 3146 7834
rect 3146 7806 3148 7834
rect 3116 7804 3148 7806
rect 3116 7674 3148 7676
rect 3116 7646 3118 7674
rect 3118 7646 3146 7674
rect 3146 7646 3148 7674
rect 3116 7644 3148 7646
rect 3116 7514 3148 7516
rect 3116 7486 3118 7514
rect 3118 7486 3146 7514
rect 3146 7486 3148 7514
rect 3116 7484 3148 7486
rect 3116 7354 3148 7356
rect 3116 7326 3118 7354
rect 3118 7326 3146 7354
rect 3146 7326 3148 7354
rect 3116 7324 3148 7326
rect 3116 7194 3148 7196
rect 3116 7166 3118 7194
rect 3118 7166 3146 7194
rect 3146 7166 3148 7194
rect 3116 7164 3148 7166
rect 3116 7034 3148 7036
rect 3116 7006 3118 7034
rect 3118 7006 3146 7034
rect 3146 7006 3148 7034
rect 3116 7004 3148 7006
rect 3116 6874 3148 6876
rect 3116 6846 3118 6874
rect 3118 6846 3146 6874
rect 3146 6846 3148 6874
rect 3116 6844 3148 6846
rect 3116 6714 3148 6716
rect 3116 6686 3118 6714
rect 3118 6686 3146 6714
rect 3146 6686 3148 6714
rect 3116 6684 3148 6686
rect 3116 6554 3148 6556
rect 3116 6526 3118 6554
rect 3118 6526 3146 6554
rect 3146 6526 3148 6554
rect 3116 6524 3148 6526
rect 3116 6394 3148 6396
rect 3116 6366 3118 6394
rect 3118 6366 3146 6394
rect 3146 6366 3148 6394
rect 3116 6364 3148 6366
rect 3116 6234 3148 6236
rect 3116 6206 3118 6234
rect 3118 6206 3146 6234
rect 3146 6206 3148 6234
rect 3116 6204 3148 6206
rect 3116 6074 3148 6076
rect 3116 6046 3118 6074
rect 3118 6046 3146 6074
rect 3146 6046 3148 6074
rect 3116 6044 3148 6046
rect 3116 5914 3148 5916
rect 3116 5886 3118 5914
rect 3118 5886 3146 5914
rect 3146 5886 3148 5914
rect 3116 5884 3148 5886
rect 6849 9114 6881 9116
rect 6849 9086 6851 9114
rect 6851 9086 6879 9114
rect 6879 9086 6881 9114
rect 6849 9084 6881 9086
rect 6849 8954 6881 8956
rect 6849 8926 6851 8954
rect 6851 8926 6879 8954
rect 6879 8926 6881 8954
rect 6849 8924 6881 8926
rect 6849 8794 6881 8796
rect 6849 8766 6851 8794
rect 6851 8766 6879 8794
rect 6879 8766 6881 8794
rect 6849 8764 6881 8766
rect 6849 8634 6881 8636
rect 6849 8606 6851 8634
rect 6851 8606 6879 8634
rect 6879 8606 6881 8634
rect 6849 8604 6881 8606
rect 6849 8474 6881 8476
rect 6849 8446 6851 8474
rect 6851 8446 6879 8474
rect 6879 8446 6881 8474
rect 6849 8444 6881 8446
rect 6849 8314 6881 8316
rect 6849 8286 6851 8314
rect 6851 8286 6879 8314
rect 6879 8286 6881 8314
rect 6849 8284 6881 8286
rect 6849 8154 6881 8156
rect 6849 8126 6851 8154
rect 6851 8126 6879 8154
rect 6879 8126 6881 8154
rect 6849 8124 6881 8126
rect 6849 7994 6881 7996
rect 6849 7966 6851 7994
rect 6851 7966 6879 7994
rect 6879 7966 6881 7994
rect 6849 7964 6881 7966
rect 6849 7834 6881 7836
rect 6849 7806 6851 7834
rect 6851 7806 6879 7834
rect 6879 7806 6881 7834
rect 6849 7804 6881 7806
rect 6849 7674 6881 7676
rect 6849 7646 6851 7674
rect 6851 7646 6879 7674
rect 6879 7646 6881 7674
rect 6849 7644 6881 7646
rect 6849 7514 6881 7516
rect 6849 7486 6851 7514
rect 6851 7486 6879 7514
rect 6879 7486 6881 7514
rect 6849 7484 6881 7486
rect 6849 7354 6881 7356
rect 6849 7326 6851 7354
rect 6851 7326 6879 7354
rect 6879 7326 6881 7354
rect 6849 7324 6881 7326
rect 6849 7194 6881 7196
rect 6849 7166 6851 7194
rect 6851 7166 6879 7194
rect 6879 7166 6881 7194
rect 6849 7164 6881 7166
rect 6849 7034 6881 7036
rect 6849 7006 6851 7034
rect 6851 7006 6879 7034
rect 6879 7006 6881 7034
rect 6849 7004 6881 7006
rect 6849 6874 6881 6876
rect 6849 6846 6851 6874
rect 6851 6846 6879 6874
rect 6879 6846 6881 6874
rect 6849 6844 6881 6846
rect 6849 6714 6881 6716
rect 6849 6686 6851 6714
rect 6851 6686 6879 6714
rect 6879 6686 6881 6714
rect 6849 6684 6881 6686
rect 6849 6554 6881 6556
rect 6849 6526 6851 6554
rect 6851 6526 6879 6554
rect 6879 6526 6881 6554
rect 6849 6524 6881 6526
rect 6849 6394 6881 6396
rect 6849 6366 6851 6394
rect 6851 6366 6879 6394
rect 6879 6366 6881 6394
rect 6849 6364 6881 6366
rect 6849 6234 6881 6236
rect 6849 6206 6851 6234
rect 6851 6206 6879 6234
rect 6879 6206 6881 6234
rect 6849 6204 6881 6206
rect 6849 6074 6881 6076
rect 6849 6046 6851 6074
rect 6851 6046 6879 6074
rect 6879 6046 6881 6074
rect 6849 6044 6881 6046
rect 6849 5914 6881 5916
rect 6849 5886 6851 5914
rect 6851 5886 6879 5914
rect 6879 5886 6881 5914
rect 6849 5884 6881 5886
rect 3116 5754 3148 5756
rect 3116 5726 3118 5754
rect 3118 5726 3146 5754
rect 3146 5726 3148 5754
rect 3116 5724 3148 5726
rect 6849 5754 6881 5756
rect 6849 5726 6851 5754
rect 6851 5726 6879 5754
rect 6879 5726 6881 5754
rect 6849 5724 6881 5726
rect 3304 5651 3336 5653
rect 3304 5623 3306 5651
rect 3306 5623 3334 5651
rect 3334 5623 3336 5651
rect 3304 5621 3336 5623
rect 3464 5651 3496 5653
rect 3464 5623 3466 5651
rect 3466 5623 3494 5651
rect 3494 5623 3496 5651
rect 3464 5621 3496 5623
rect 3624 5651 3656 5653
rect 3624 5623 3626 5651
rect 3626 5623 3654 5651
rect 3654 5623 3656 5651
rect 3624 5621 3656 5623
rect 3784 5651 3816 5653
rect 3784 5623 3786 5651
rect 3786 5623 3814 5651
rect 3814 5623 3816 5651
rect 3784 5621 3816 5623
rect 3944 5651 3976 5653
rect 3944 5623 3946 5651
rect 3946 5623 3974 5651
rect 3974 5623 3976 5651
rect 3944 5621 3976 5623
rect 4104 5651 4136 5653
rect 4104 5623 4106 5651
rect 4106 5623 4134 5651
rect 4134 5623 4136 5651
rect 4104 5621 4136 5623
rect 4264 5651 4296 5653
rect 4264 5623 4266 5651
rect 4266 5623 4294 5651
rect 4294 5623 4296 5651
rect 4264 5621 4296 5623
rect 4424 5651 4456 5653
rect 4424 5623 4426 5651
rect 4426 5623 4454 5651
rect 4454 5623 4456 5651
rect 4424 5621 4456 5623
rect 4584 5651 4616 5653
rect 4584 5623 4586 5651
rect 4586 5623 4614 5651
rect 4614 5623 4616 5651
rect 4584 5621 4616 5623
rect 4744 5651 4776 5653
rect 4744 5623 4746 5651
rect 4746 5623 4774 5651
rect 4774 5623 4776 5651
rect 4744 5621 4776 5623
rect 4904 5651 4936 5653
rect 4904 5623 4906 5651
rect 4906 5623 4934 5651
rect 4934 5623 4936 5651
rect 4904 5621 4936 5623
rect 5064 5651 5096 5653
rect 5064 5623 5066 5651
rect 5066 5623 5094 5651
rect 5094 5623 5096 5651
rect 5064 5621 5096 5623
rect 5224 5651 5256 5653
rect 5224 5623 5226 5651
rect 5226 5623 5254 5651
rect 5254 5623 5256 5651
rect 5224 5621 5256 5623
rect 5384 5651 5416 5653
rect 5384 5623 5386 5651
rect 5386 5623 5414 5651
rect 5414 5623 5416 5651
rect 5384 5621 5416 5623
rect 5544 5651 5576 5653
rect 5544 5623 5546 5651
rect 5546 5623 5574 5651
rect 5574 5623 5576 5651
rect 5544 5621 5576 5623
rect 5704 5651 5736 5653
rect 5704 5623 5706 5651
rect 5706 5623 5734 5651
rect 5734 5623 5736 5651
rect 5704 5621 5736 5623
rect 5864 5651 5896 5653
rect 5864 5623 5866 5651
rect 5866 5623 5894 5651
rect 5894 5623 5896 5651
rect 5864 5621 5896 5623
rect 6024 5651 6056 5653
rect 6024 5623 6026 5651
rect 6026 5623 6054 5651
rect 6054 5623 6056 5651
rect 6024 5621 6056 5623
rect 6184 5651 6216 5653
rect 6184 5623 6186 5651
rect 6186 5623 6214 5651
rect 6214 5623 6216 5651
rect 6184 5621 6216 5623
rect 6344 5651 6376 5653
rect 6344 5623 6346 5651
rect 6346 5623 6374 5651
rect 6374 5623 6376 5651
rect 6344 5621 6376 5623
rect 6504 5651 6536 5653
rect 6504 5623 6506 5651
rect 6506 5623 6534 5651
rect 6534 5623 6536 5651
rect 6504 5621 6536 5623
rect 6664 5651 6696 5653
rect 6664 5623 6666 5651
rect 6666 5623 6694 5651
rect 6694 5623 6696 5651
rect 6664 5621 6696 5623
rect 9304 9379 9336 9381
rect 9304 9351 9306 9379
rect 9306 9351 9334 9379
rect 9334 9351 9336 9379
rect 9304 9349 9336 9351
rect 9464 9379 9496 9381
rect 9464 9351 9466 9379
rect 9466 9351 9494 9379
rect 9494 9351 9496 9379
rect 9464 9349 9496 9351
rect 9624 9379 9656 9381
rect 9624 9351 9626 9379
rect 9626 9351 9654 9379
rect 9654 9351 9656 9379
rect 9624 9349 9656 9351
rect 9784 9379 9816 9381
rect 9784 9351 9786 9379
rect 9786 9351 9814 9379
rect 9814 9351 9816 9379
rect 9784 9349 9816 9351
rect 9944 9379 9976 9381
rect 9944 9351 9946 9379
rect 9946 9351 9974 9379
rect 9974 9351 9976 9379
rect 9944 9349 9976 9351
rect 10104 9379 10136 9381
rect 10104 9351 10106 9379
rect 10106 9351 10134 9379
rect 10134 9351 10136 9379
rect 10104 9349 10136 9351
rect 10264 9379 10296 9381
rect 10264 9351 10266 9379
rect 10266 9351 10294 9379
rect 10294 9351 10296 9379
rect 10264 9349 10296 9351
rect 10424 9379 10456 9381
rect 10424 9351 10426 9379
rect 10426 9351 10454 9379
rect 10454 9351 10456 9379
rect 10424 9349 10456 9351
rect 10584 9379 10616 9381
rect 10584 9351 10586 9379
rect 10586 9351 10614 9379
rect 10614 9351 10616 9379
rect 10584 9349 10616 9351
rect 10744 9379 10776 9381
rect 10744 9351 10746 9379
rect 10746 9351 10774 9379
rect 10774 9351 10776 9379
rect 10744 9349 10776 9351
rect 10904 9379 10936 9381
rect 10904 9351 10906 9379
rect 10906 9351 10934 9379
rect 10934 9351 10936 9379
rect 10904 9349 10936 9351
rect 11064 9379 11096 9381
rect 11064 9351 11066 9379
rect 11066 9351 11094 9379
rect 11094 9351 11096 9379
rect 11064 9349 11096 9351
rect 11224 9379 11256 9381
rect 11224 9351 11226 9379
rect 11226 9351 11254 9379
rect 11254 9351 11256 9379
rect 11224 9349 11256 9351
rect 11384 9379 11416 9381
rect 11384 9351 11386 9379
rect 11386 9351 11414 9379
rect 11414 9351 11416 9379
rect 11384 9349 11416 9351
rect 11544 9379 11576 9381
rect 11544 9351 11546 9379
rect 11546 9351 11574 9379
rect 11574 9351 11576 9379
rect 11544 9349 11576 9351
rect 11704 9379 11736 9381
rect 11704 9351 11706 9379
rect 11706 9351 11734 9379
rect 11734 9351 11736 9379
rect 11704 9349 11736 9351
rect 11864 9379 11896 9381
rect 11864 9351 11866 9379
rect 11866 9351 11894 9379
rect 11894 9351 11896 9379
rect 11864 9349 11896 9351
rect 12024 9379 12056 9381
rect 12024 9351 12026 9379
rect 12026 9351 12054 9379
rect 12054 9351 12056 9379
rect 12024 9349 12056 9351
rect 12184 9379 12216 9381
rect 12184 9351 12186 9379
rect 12186 9351 12214 9379
rect 12214 9351 12216 9379
rect 12184 9349 12216 9351
rect 12344 9379 12376 9381
rect 12344 9351 12346 9379
rect 12346 9351 12374 9379
rect 12374 9351 12376 9379
rect 12344 9349 12376 9351
rect 12504 9379 12536 9381
rect 12504 9351 12506 9379
rect 12506 9351 12534 9379
rect 12534 9351 12536 9379
rect 12504 9349 12536 9351
rect 12664 9379 12696 9381
rect 12664 9351 12666 9379
rect 12666 9351 12694 9379
rect 12694 9351 12696 9379
rect 12664 9349 12696 9351
rect 9116 9274 9148 9276
rect 9116 9246 9118 9274
rect 9118 9246 9146 9274
rect 9146 9246 9148 9274
rect 9116 9244 9148 9246
rect 12849 9274 12881 9276
rect 12849 9246 12851 9274
rect 12851 9246 12879 9274
rect 12879 9246 12881 9274
rect 12849 9244 12881 9246
rect 9116 9114 9148 9116
rect 9116 9086 9118 9114
rect 9118 9086 9146 9114
rect 9146 9086 9148 9114
rect 9116 9084 9148 9086
rect 9116 8954 9148 8956
rect 9116 8926 9118 8954
rect 9118 8926 9146 8954
rect 9146 8926 9148 8954
rect 9116 8924 9148 8926
rect 9116 8794 9148 8796
rect 9116 8766 9118 8794
rect 9118 8766 9146 8794
rect 9146 8766 9148 8794
rect 9116 8764 9148 8766
rect 9116 8634 9148 8636
rect 9116 8606 9118 8634
rect 9118 8606 9146 8634
rect 9146 8606 9148 8634
rect 9116 8604 9148 8606
rect 9116 8474 9148 8476
rect 9116 8446 9118 8474
rect 9118 8446 9146 8474
rect 9146 8446 9148 8474
rect 9116 8444 9148 8446
rect 9116 8314 9148 8316
rect 9116 8286 9118 8314
rect 9118 8286 9146 8314
rect 9146 8286 9148 8314
rect 9116 8284 9148 8286
rect 9116 8154 9148 8156
rect 9116 8126 9118 8154
rect 9118 8126 9146 8154
rect 9146 8126 9148 8154
rect 9116 8124 9148 8126
rect 9116 7994 9148 7996
rect 9116 7966 9118 7994
rect 9118 7966 9146 7994
rect 9146 7966 9148 7994
rect 9116 7964 9148 7966
rect 9116 7834 9148 7836
rect 9116 7806 9118 7834
rect 9118 7806 9146 7834
rect 9146 7806 9148 7834
rect 9116 7804 9148 7806
rect 9116 7674 9148 7676
rect 9116 7646 9118 7674
rect 9118 7646 9146 7674
rect 9146 7646 9148 7674
rect 9116 7644 9148 7646
rect 9116 7514 9148 7516
rect 9116 7486 9118 7514
rect 9118 7486 9146 7514
rect 9146 7486 9148 7514
rect 9116 7484 9148 7486
rect 9116 7354 9148 7356
rect 9116 7326 9118 7354
rect 9118 7326 9146 7354
rect 9146 7326 9148 7354
rect 9116 7324 9148 7326
rect 9116 7194 9148 7196
rect 9116 7166 9118 7194
rect 9118 7166 9146 7194
rect 9146 7166 9148 7194
rect 9116 7164 9148 7166
rect 9116 7034 9148 7036
rect 9116 7006 9118 7034
rect 9118 7006 9146 7034
rect 9146 7006 9148 7034
rect 9116 7004 9148 7006
rect 9116 6874 9148 6876
rect 9116 6846 9118 6874
rect 9118 6846 9146 6874
rect 9146 6846 9148 6874
rect 9116 6844 9148 6846
rect 9116 6714 9148 6716
rect 9116 6686 9118 6714
rect 9118 6686 9146 6714
rect 9146 6686 9148 6714
rect 9116 6684 9148 6686
rect 9116 6554 9148 6556
rect 9116 6526 9118 6554
rect 9118 6526 9146 6554
rect 9146 6526 9148 6554
rect 9116 6524 9148 6526
rect 9116 6394 9148 6396
rect 9116 6366 9118 6394
rect 9118 6366 9146 6394
rect 9146 6366 9148 6394
rect 9116 6364 9148 6366
rect 9116 6234 9148 6236
rect 9116 6206 9118 6234
rect 9118 6206 9146 6234
rect 9146 6206 9148 6234
rect 9116 6204 9148 6206
rect 9116 6074 9148 6076
rect 9116 6046 9118 6074
rect 9118 6046 9146 6074
rect 9146 6046 9148 6074
rect 9116 6044 9148 6046
rect 9116 5914 9148 5916
rect 9116 5886 9118 5914
rect 9118 5886 9146 5914
rect 9146 5886 9148 5914
rect 9116 5884 9148 5886
rect 12849 9114 12881 9116
rect 12849 9086 12851 9114
rect 12851 9086 12879 9114
rect 12879 9086 12881 9114
rect 12849 9084 12881 9086
rect 12849 8954 12881 8956
rect 12849 8926 12851 8954
rect 12851 8926 12879 8954
rect 12879 8926 12881 8954
rect 12849 8924 12881 8926
rect 12849 8794 12881 8796
rect 12849 8766 12851 8794
rect 12851 8766 12879 8794
rect 12879 8766 12881 8794
rect 12849 8764 12881 8766
rect 12849 8634 12881 8636
rect 12849 8606 12851 8634
rect 12851 8606 12879 8634
rect 12879 8606 12881 8634
rect 12849 8604 12881 8606
rect 12849 8474 12881 8476
rect 12849 8446 12851 8474
rect 12851 8446 12879 8474
rect 12879 8446 12881 8474
rect 12849 8444 12881 8446
rect 12849 8314 12881 8316
rect 12849 8286 12851 8314
rect 12851 8286 12879 8314
rect 12879 8286 12881 8314
rect 12849 8284 12881 8286
rect 12849 8154 12881 8156
rect 12849 8126 12851 8154
rect 12851 8126 12879 8154
rect 12879 8126 12881 8154
rect 12849 8124 12881 8126
rect 12849 7994 12881 7996
rect 12849 7966 12851 7994
rect 12851 7966 12879 7994
rect 12879 7966 12881 7994
rect 12849 7964 12881 7966
rect 12849 7834 12881 7836
rect 12849 7806 12851 7834
rect 12851 7806 12879 7834
rect 12879 7806 12881 7834
rect 12849 7804 12881 7806
rect 12849 7674 12881 7676
rect 12849 7646 12851 7674
rect 12851 7646 12879 7674
rect 12879 7646 12881 7674
rect 12849 7644 12881 7646
rect 12849 7514 12881 7516
rect 12849 7486 12851 7514
rect 12851 7486 12879 7514
rect 12879 7486 12881 7514
rect 12849 7484 12881 7486
rect 12849 7354 12881 7356
rect 12849 7326 12851 7354
rect 12851 7326 12879 7354
rect 12879 7326 12881 7354
rect 12849 7324 12881 7326
rect 12849 7194 12881 7196
rect 12849 7166 12851 7194
rect 12851 7166 12879 7194
rect 12879 7166 12881 7194
rect 12849 7164 12881 7166
rect 12849 7034 12881 7036
rect 12849 7006 12851 7034
rect 12851 7006 12879 7034
rect 12879 7006 12881 7034
rect 12849 7004 12881 7006
rect 15304 9379 15336 9381
rect 15304 9351 15306 9379
rect 15306 9351 15334 9379
rect 15334 9351 15336 9379
rect 15304 9349 15336 9351
rect 15464 9379 15496 9381
rect 15464 9351 15466 9379
rect 15466 9351 15494 9379
rect 15494 9351 15496 9379
rect 15464 9349 15496 9351
rect 15624 9379 15656 9381
rect 15624 9351 15626 9379
rect 15626 9351 15654 9379
rect 15654 9351 15656 9379
rect 15624 9349 15656 9351
rect 15784 9379 15816 9381
rect 15784 9351 15786 9379
rect 15786 9351 15814 9379
rect 15814 9351 15816 9379
rect 15784 9349 15816 9351
rect 15944 9379 15976 9381
rect 15944 9351 15946 9379
rect 15946 9351 15974 9379
rect 15974 9351 15976 9379
rect 15944 9349 15976 9351
rect 16104 9379 16136 9381
rect 16104 9351 16106 9379
rect 16106 9351 16134 9379
rect 16134 9351 16136 9379
rect 16104 9349 16136 9351
rect 16264 9379 16296 9381
rect 16264 9351 16266 9379
rect 16266 9351 16294 9379
rect 16294 9351 16296 9379
rect 16264 9349 16296 9351
rect 16424 9379 16456 9381
rect 16424 9351 16426 9379
rect 16426 9351 16454 9379
rect 16454 9351 16456 9379
rect 16424 9349 16456 9351
rect 16584 9379 16616 9381
rect 16584 9351 16586 9379
rect 16586 9351 16614 9379
rect 16614 9351 16616 9379
rect 16584 9349 16616 9351
rect 16744 9379 16776 9381
rect 16744 9351 16746 9379
rect 16746 9351 16774 9379
rect 16774 9351 16776 9379
rect 16744 9349 16776 9351
rect 16904 9379 16936 9381
rect 16904 9351 16906 9379
rect 16906 9351 16934 9379
rect 16934 9351 16936 9379
rect 16904 9349 16936 9351
rect 17064 9379 17096 9381
rect 17064 9351 17066 9379
rect 17066 9351 17094 9379
rect 17094 9351 17096 9379
rect 17064 9349 17096 9351
rect 17224 9379 17256 9381
rect 17224 9351 17226 9379
rect 17226 9351 17254 9379
rect 17254 9351 17256 9379
rect 17224 9349 17256 9351
rect 17384 9379 17416 9381
rect 17384 9351 17386 9379
rect 17386 9351 17414 9379
rect 17414 9351 17416 9379
rect 17384 9349 17416 9351
rect 17544 9379 17576 9381
rect 17544 9351 17546 9379
rect 17546 9351 17574 9379
rect 17574 9351 17576 9379
rect 17544 9349 17576 9351
rect 17704 9379 17736 9381
rect 17704 9351 17706 9379
rect 17706 9351 17734 9379
rect 17734 9351 17736 9379
rect 17704 9349 17736 9351
rect 17864 9379 17896 9381
rect 17864 9351 17866 9379
rect 17866 9351 17894 9379
rect 17894 9351 17896 9379
rect 17864 9349 17896 9351
rect 18024 9379 18056 9381
rect 18024 9351 18026 9379
rect 18026 9351 18054 9379
rect 18054 9351 18056 9379
rect 18024 9349 18056 9351
rect 18184 9379 18216 9381
rect 18184 9351 18186 9379
rect 18186 9351 18214 9379
rect 18214 9351 18216 9379
rect 18184 9349 18216 9351
rect 18344 9379 18376 9381
rect 18344 9351 18346 9379
rect 18346 9351 18374 9379
rect 18374 9351 18376 9379
rect 18344 9349 18376 9351
rect 18504 9379 18536 9381
rect 18504 9351 18506 9379
rect 18506 9351 18534 9379
rect 18534 9351 18536 9379
rect 18504 9349 18536 9351
rect 18664 9379 18696 9381
rect 18664 9351 18666 9379
rect 18666 9351 18694 9379
rect 18694 9351 18696 9379
rect 18664 9349 18696 9351
rect 15116 9274 15148 9276
rect 15116 9246 15118 9274
rect 15118 9246 15146 9274
rect 15146 9246 15148 9274
rect 15116 9244 15148 9246
rect 18849 9274 18881 9276
rect 18849 9246 18851 9274
rect 18851 9246 18879 9274
rect 18879 9246 18881 9274
rect 18849 9244 18881 9246
rect 15116 9114 15148 9116
rect 15116 9086 15118 9114
rect 15118 9086 15146 9114
rect 15146 9086 15148 9114
rect 15116 9084 15148 9086
rect 15116 8954 15148 8956
rect 15116 8926 15118 8954
rect 15118 8926 15146 8954
rect 15146 8926 15148 8954
rect 15116 8924 15148 8926
rect 15116 8794 15148 8796
rect 15116 8766 15118 8794
rect 15118 8766 15146 8794
rect 15146 8766 15148 8794
rect 15116 8764 15148 8766
rect 15116 8634 15148 8636
rect 15116 8606 15118 8634
rect 15118 8606 15146 8634
rect 15146 8606 15148 8634
rect 15116 8604 15148 8606
rect 15116 8474 15148 8476
rect 15116 8446 15118 8474
rect 15118 8446 15146 8474
rect 15146 8446 15148 8474
rect 15116 8444 15148 8446
rect 15116 8314 15148 8316
rect 15116 8286 15118 8314
rect 15118 8286 15146 8314
rect 15146 8286 15148 8314
rect 15116 8284 15148 8286
rect 15116 8154 15148 8156
rect 15116 8126 15118 8154
rect 15118 8126 15146 8154
rect 15146 8126 15148 8154
rect 15116 8124 15148 8126
rect 15116 7994 15148 7996
rect 15116 7966 15118 7994
rect 15118 7966 15146 7994
rect 15146 7966 15148 7994
rect 15116 7964 15148 7966
rect 15116 7834 15148 7836
rect 15116 7806 15118 7834
rect 15118 7806 15146 7834
rect 15146 7806 15148 7834
rect 15116 7804 15148 7806
rect 15116 7674 15148 7676
rect 15116 7646 15118 7674
rect 15118 7646 15146 7674
rect 15146 7646 15148 7674
rect 15116 7644 15148 7646
rect 15116 7514 15148 7516
rect 15116 7486 15118 7514
rect 15118 7486 15146 7514
rect 15146 7486 15148 7514
rect 15116 7484 15148 7486
rect 15116 7354 15148 7356
rect 15116 7326 15118 7354
rect 15118 7326 15146 7354
rect 15146 7326 15148 7354
rect 15116 7324 15148 7326
rect 15116 7194 15148 7196
rect 15116 7166 15118 7194
rect 15118 7166 15146 7194
rect 15146 7166 15148 7194
rect 15116 7164 15148 7166
rect 15116 7034 15148 7036
rect 15116 7006 15118 7034
rect 15118 7006 15146 7034
rect 15146 7006 15148 7034
rect 15116 7004 15148 7006
rect 12849 6874 12881 6876
rect 12849 6846 12851 6874
rect 12851 6846 12879 6874
rect 12879 6846 12881 6874
rect 12849 6844 12881 6846
rect 12849 6714 12881 6716
rect 12849 6686 12851 6714
rect 12851 6686 12879 6714
rect 12879 6686 12881 6714
rect 12849 6684 12881 6686
rect 12849 6554 12881 6556
rect 12849 6526 12851 6554
rect 12851 6526 12879 6554
rect 12879 6526 12881 6554
rect 12849 6524 12881 6526
rect 12849 6394 12881 6396
rect 12849 6366 12851 6394
rect 12851 6366 12879 6394
rect 12879 6366 12881 6394
rect 12849 6364 12881 6366
rect 12849 6234 12881 6236
rect 12849 6206 12851 6234
rect 12851 6206 12879 6234
rect 12879 6206 12881 6234
rect 12849 6204 12881 6206
rect 12849 6074 12881 6076
rect 12849 6046 12851 6074
rect 12851 6046 12879 6074
rect 12879 6046 12881 6074
rect 12849 6044 12881 6046
rect 12849 5914 12881 5916
rect 12849 5886 12851 5914
rect 12851 5886 12879 5914
rect 12879 5886 12881 5914
rect 12849 5884 12881 5886
rect 9116 5754 9148 5756
rect 9116 5726 9118 5754
rect 9118 5726 9146 5754
rect 9146 5726 9148 5754
rect 9116 5724 9148 5726
rect 12849 5754 12881 5756
rect 12849 5726 12851 5754
rect 12851 5726 12879 5754
rect 12879 5726 12881 5754
rect 12849 5724 12881 5726
rect 9304 5651 9336 5653
rect 9304 5623 9306 5651
rect 9306 5623 9334 5651
rect 9334 5623 9336 5651
rect 9304 5621 9336 5623
rect 9464 5651 9496 5653
rect 9464 5623 9466 5651
rect 9466 5623 9494 5651
rect 9494 5623 9496 5651
rect 9464 5621 9496 5623
rect 9624 5651 9656 5653
rect 9624 5623 9626 5651
rect 9626 5623 9654 5651
rect 9654 5623 9656 5651
rect 9624 5621 9656 5623
rect 9784 5651 9816 5653
rect 9784 5623 9786 5651
rect 9786 5623 9814 5651
rect 9814 5623 9816 5651
rect 9784 5621 9816 5623
rect 9944 5651 9976 5653
rect 9944 5623 9946 5651
rect 9946 5623 9974 5651
rect 9974 5623 9976 5651
rect 9944 5621 9976 5623
rect 10104 5651 10136 5653
rect 10104 5623 10106 5651
rect 10106 5623 10134 5651
rect 10134 5623 10136 5651
rect 10104 5621 10136 5623
rect 10264 5651 10296 5653
rect 10264 5623 10266 5651
rect 10266 5623 10294 5651
rect 10294 5623 10296 5651
rect 10264 5621 10296 5623
rect 10424 5651 10456 5653
rect 10424 5623 10426 5651
rect 10426 5623 10454 5651
rect 10454 5623 10456 5651
rect 10424 5621 10456 5623
rect 10584 5651 10616 5653
rect 10584 5623 10586 5651
rect 10586 5623 10614 5651
rect 10614 5623 10616 5651
rect 10584 5621 10616 5623
rect 10744 5651 10776 5653
rect 10744 5623 10746 5651
rect 10746 5623 10774 5651
rect 10774 5623 10776 5651
rect 10744 5621 10776 5623
rect 10904 5651 10936 5653
rect 10904 5623 10906 5651
rect 10906 5623 10934 5651
rect 10934 5623 10936 5651
rect 10904 5621 10936 5623
rect 11064 5651 11096 5653
rect 11064 5623 11066 5651
rect 11066 5623 11094 5651
rect 11094 5623 11096 5651
rect 11064 5621 11096 5623
rect 11224 5651 11256 5653
rect 11224 5623 11226 5651
rect 11226 5623 11254 5651
rect 11254 5623 11256 5651
rect 11224 5621 11256 5623
rect 11384 5651 11416 5653
rect 11384 5623 11386 5651
rect 11386 5623 11414 5651
rect 11414 5623 11416 5651
rect 11384 5621 11416 5623
rect 11544 5651 11576 5653
rect 11544 5623 11546 5651
rect 11546 5623 11574 5651
rect 11574 5623 11576 5651
rect 11544 5621 11576 5623
rect 11704 5651 11736 5653
rect 11704 5623 11706 5651
rect 11706 5623 11734 5651
rect 11734 5623 11736 5651
rect 11704 5621 11736 5623
rect 11864 5651 11896 5653
rect 11864 5623 11866 5651
rect 11866 5623 11894 5651
rect 11894 5623 11896 5651
rect 11864 5621 11896 5623
rect 12024 5651 12056 5653
rect 12024 5623 12026 5651
rect 12026 5623 12054 5651
rect 12054 5623 12056 5651
rect 12024 5621 12056 5623
rect 12184 5651 12216 5653
rect 12184 5623 12186 5651
rect 12186 5623 12214 5651
rect 12214 5623 12216 5651
rect 12184 5621 12216 5623
rect 12344 5651 12376 5653
rect 12344 5623 12346 5651
rect 12346 5623 12374 5651
rect 12374 5623 12376 5651
rect 12344 5621 12376 5623
rect 12504 5651 12536 5653
rect 12504 5623 12506 5651
rect 12506 5623 12534 5651
rect 12534 5623 12536 5651
rect 12504 5621 12536 5623
rect 12664 5651 12696 5653
rect 12664 5623 12666 5651
rect 12666 5623 12694 5651
rect 12694 5623 12696 5651
rect 12664 5621 12696 5623
rect 15116 6874 15148 6876
rect 15116 6846 15118 6874
rect 15118 6846 15146 6874
rect 15146 6846 15148 6874
rect 15116 6844 15148 6846
rect 15116 6714 15148 6716
rect 15116 6686 15118 6714
rect 15118 6686 15146 6714
rect 15146 6686 15148 6714
rect 15116 6684 15148 6686
rect 15116 6554 15148 6556
rect 15116 6526 15118 6554
rect 15118 6526 15146 6554
rect 15146 6526 15148 6554
rect 15116 6524 15148 6526
rect 15116 6394 15148 6396
rect 15116 6366 15118 6394
rect 15118 6366 15146 6394
rect 15146 6366 15148 6394
rect 15116 6364 15148 6366
rect 15116 6234 15148 6236
rect 15116 6206 15118 6234
rect 15118 6206 15146 6234
rect 15146 6206 15148 6234
rect 15116 6204 15148 6206
rect 15116 6074 15148 6076
rect 15116 6046 15118 6074
rect 15118 6046 15146 6074
rect 15146 6046 15148 6074
rect 15116 6044 15148 6046
rect 15116 5914 15148 5916
rect 15116 5886 15118 5914
rect 15118 5886 15146 5914
rect 15146 5886 15148 5914
rect 15116 5884 15148 5886
rect 18849 9114 18881 9116
rect 18849 9086 18851 9114
rect 18851 9086 18879 9114
rect 18879 9086 18881 9114
rect 18849 9084 18881 9086
rect 18849 8954 18881 8956
rect 18849 8926 18851 8954
rect 18851 8926 18879 8954
rect 18879 8926 18881 8954
rect 18849 8924 18881 8926
rect 18849 8794 18881 8796
rect 18849 8766 18851 8794
rect 18851 8766 18879 8794
rect 18879 8766 18881 8794
rect 18849 8764 18881 8766
rect 18849 8634 18881 8636
rect 18849 8606 18851 8634
rect 18851 8606 18879 8634
rect 18879 8606 18881 8634
rect 18849 8604 18881 8606
rect 18849 8474 18881 8476
rect 18849 8446 18851 8474
rect 18851 8446 18879 8474
rect 18879 8446 18881 8474
rect 18849 8444 18881 8446
rect 18849 8314 18881 8316
rect 18849 8286 18851 8314
rect 18851 8286 18879 8314
rect 18879 8286 18881 8314
rect 18849 8284 18881 8286
rect 18849 8154 18881 8156
rect 18849 8126 18851 8154
rect 18851 8126 18879 8154
rect 18879 8126 18881 8154
rect 18849 8124 18881 8126
rect 18849 7994 18881 7996
rect 18849 7966 18851 7994
rect 18851 7966 18879 7994
rect 18879 7966 18881 7994
rect 18849 7964 18881 7966
rect 18849 7834 18881 7836
rect 18849 7806 18851 7834
rect 18851 7806 18879 7834
rect 18879 7806 18881 7834
rect 18849 7804 18881 7806
rect 18849 7674 18881 7676
rect 18849 7646 18851 7674
rect 18851 7646 18879 7674
rect 18879 7646 18881 7674
rect 18849 7644 18881 7646
rect 18849 7514 18881 7516
rect 18849 7486 18851 7514
rect 18851 7486 18879 7514
rect 18879 7486 18881 7514
rect 18849 7484 18881 7486
rect 18849 7354 18881 7356
rect 18849 7326 18851 7354
rect 18851 7326 18879 7354
rect 18879 7326 18881 7354
rect 18849 7324 18881 7326
rect 18849 7194 18881 7196
rect 18849 7166 18851 7194
rect 18851 7166 18879 7194
rect 18879 7166 18881 7194
rect 18849 7164 18881 7166
rect 18849 7034 18881 7036
rect 18849 7006 18851 7034
rect 18851 7006 18879 7034
rect 18879 7006 18881 7034
rect 18849 7004 18881 7006
rect 21304 9379 21336 9381
rect 21304 9351 21306 9379
rect 21306 9351 21334 9379
rect 21334 9351 21336 9379
rect 21304 9349 21336 9351
rect 21464 9379 21496 9381
rect 21464 9351 21466 9379
rect 21466 9351 21494 9379
rect 21494 9351 21496 9379
rect 21464 9349 21496 9351
rect 21624 9379 21656 9381
rect 21624 9351 21626 9379
rect 21626 9351 21654 9379
rect 21654 9351 21656 9379
rect 21624 9349 21656 9351
rect 21784 9379 21816 9381
rect 21784 9351 21786 9379
rect 21786 9351 21814 9379
rect 21814 9351 21816 9379
rect 21784 9349 21816 9351
rect 21944 9379 21976 9381
rect 21944 9351 21946 9379
rect 21946 9351 21974 9379
rect 21974 9351 21976 9379
rect 21944 9349 21976 9351
rect 22104 9379 22136 9381
rect 22104 9351 22106 9379
rect 22106 9351 22134 9379
rect 22134 9351 22136 9379
rect 22104 9349 22136 9351
rect 22264 9379 22296 9381
rect 22264 9351 22266 9379
rect 22266 9351 22294 9379
rect 22294 9351 22296 9379
rect 22264 9349 22296 9351
rect 22424 9379 22456 9381
rect 22424 9351 22426 9379
rect 22426 9351 22454 9379
rect 22454 9351 22456 9379
rect 22424 9349 22456 9351
rect 22584 9379 22616 9381
rect 22584 9351 22586 9379
rect 22586 9351 22614 9379
rect 22614 9351 22616 9379
rect 22584 9349 22616 9351
rect 22744 9379 22776 9381
rect 22744 9351 22746 9379
rect 22746 9351 22774 9379
rect 22774 9351 22776 9379
rect 22744 9349 22776 9351
rect 22904 9379 22936 9381
rect 22904 9351 22906 9379
rect 22906 9351 22934 9379
rect 22934 9351 22936 9379
rect 22904 9349 22936 9351
rect 23064 9379 23096 9381
rect 23064 9351 23066 9379
rect 23066 9351 23094 9379
rect 23094 9351 23096 9379
rect 23064 9349 23096 9351
rect 23224 9379 23256 9381
rect 23224 9351 23226 9379
rect 23226 9351 23254 9379
rect 23254 9351 23256 9379
rect 23224 9349 23256 9351
rect 23384 9379 23416 9381
rect 23384 9351 23386 9379
rect 23386 9351 23414 9379
rect 23414 9351 23416 9379
rect 23384 9349 23416 9351
rect 23544 9379 23576 9381
rect 23544 9351 23546 9379
rect 23546 9351 23574 9379
rect 23574 9351 23576 9379
rect 23544 9349 23576 9351
rect 23704 9379 23736 9381
rect 23704 9351 23706 9379
rect 23706 9351 23734 9379
rect 23734 9351 23736 9379
rect 23704 9349 23736 9351
rect 23864 9379 23896 9381
rect 23864 9351 23866 9379
rect 23866 9351 23894 9379
rect 23894 9351 23896 9379
rect 23864 9349 23896 9351
rect 24024 9379 24056 9381
rect 24024 9351 24026 9379
rect 24026 9351 24054 9379
rect 24054 9351 24056 9379
rect 24024 9349 24056 9351
rect 24184 9379 24216 9381
rect 24184 9351 24186 9379
rect 24186 9351 24214 9379
rect 24214 9351 24216 9379
rect 24184 9349 24216 9351
rect 24344 9379 24376 9381
rect 24344 9351 24346 9379
rect 24346 9351 24374 9379
rect 24374 9351 24376 9379
rect 24344 9349 24376 9351
rect 24504 9379 24536 9381
rect 24504 9351 24506 9379
rect 24506 9351 24534 9379
rect 24534 9351 24536 9379
rect 24504 9349 24536 9351
rect 24664 9379 24696 9381
rect 24664 9351 24666 9379
rect 24666 9351 24694 9379
rect 24694 9351 24696 9379
rect 24664 9349 24696 9351
rect 21116 9274 21148 9276
rect 21116 9246 21118 9274
rect 21118 9246 21146 9274
rect 21146 9246 21148 9274
rect 21116 9244 21148 9246
rect 24849 9274 24881 9276
rect 24849 9246 24851 9274
rect 24851 9246 24879 9274
rect 24879 9246 24881 9274
rect 24849 9244 24881 9246
rect 21116 9114 21148 9116
rect 21116 9086 21118 9114
rect 21118 9086 21146 9114
rect 21146 9086 21148 9114
rect 21116 9084 21148 9086
rect 21116 8954 21148 8956
rect 21116 8926 21118 8954
rect 21118 8926 21146 8954
rect 21146 8926 21148 8954
rect 21116 8924 21148 8926
rect 21116 8794 21148 8796
rect 21116 8766 21118 8794
rect 21118 8766 21146 8794
rect 21146 8766 21148 8794
rect 21116 8764 21148 8766
rect 21116 8634 21148 8636
rect 21116 8606 21118 8634
rect 21118 8606 21146 8634
rect 21146 8606 21148 8634
rect 21116 8604 21148 8606
rect 21116 8474 21148 8476
rect 21116 8446 21118 8474
rect 21118 8446 21146 8474
rect 21146 8446 21148 8474
rect 21116 8444 21148 8446
rect 21116 8314 21148 8316
rect 21116 8286 21118 8314
rect 21118 8286 21146 8314
rect 21146 8286 21148 8314
rect 21116 8284 21148 8286
rect 21116 8154 21148 8156
rect 21116 8126 21118 8154
rect 21118 8126 21146 8154
rect 21146 8126 21148 8154
rect 21116 8124 21148 8126
rect 21116 7994 21148 7996
rect 21116 7966 21118 7994
rect 21118 7966 21146 7994
rect 21146 7966 21148 7994
rect 21116 7964 21148 7966
rect 21116 7834 21148 7836
rect 21116 7806 21118 7834
rect 21118 7806 21146 7834
rect 21146 7806 21148 7834
rect 21116 7804 21148 7806
rect 21116 7674 21148 7676
rect 21116 7646 21118 7674
rect 21118 7646 21146 7674
rect 21146 7646 21148 7674
rect 21116 7644 21148 7646
rect 21116 7514 21148 7516
rect 21116 7486 21118 7514
rect 21118 7486 21146 7514
rect 21146 7486 21148 7514
rect 21116 7484 21148 7486
rect 21116 7354 21148 7356
rect 21116 7326 21118 7354
rect 21118 7326 21146 7354
rect 21146 7326 21148 7354
rect 21116 7324 21148 7326
rect 21116 7194 21148 7196
rect 21116 7166 21118 7194
rect 21118 7166 21146 7194
rect 21146 7166 21148 7194
rect 21116 7164 21148 7166
rect 21116 7034 21148 7036
rect 21116 7006 21118 7034
rect 21118 7006 21146 7034
rect 21146 7006 21148 7034
rect 21116 7004 21148 7006
rect 18849 6874 18881 6876
rect 18849 6846 18851 6874
rect 18851 6846 18879 6874
rect 18879 6846 18881 6874
rect 18849 6844 18881 6846
rect 18849 6714 18881 6716
rect 18849 6686 18851 6714
rect 18851 6686 18879 6714
rect 18879 6686 18881 6714
rect 18849 6684 18881 6686
rect 18849 6554 18881 6556
rect 18849 6526 18851 6554
rect 18851 6526 18879 6554
rect 18879 6526 18881 6554
rect 18849 6524 18881 6526
rect 18849 6394 18881 6396
rect 18849 6366 18851 6394
rect 18851 6366 18879 6394
rect 18879 6366 18881 6394
rect 18849 6364 18881 6366
rect 18849 6234 18881 6236
rect 18849 6206 18851 6234
rect 18851 6206 18879 6234
rect 18879 6206 18881 6234
rect 18849 6204 18881 6206
rect 18849 6074 18881 6076
rect 18849 6046 18851 6074
rect 18851 6046 18879 6074
rect 18879 6046 18881 6074
rect 18849 6044 18881 6046
rect 18849 5914 18881 5916
rect 18849 5886 18851 5914
rect 18851 5886 18879 5914
rect 18879 5886 18881 5914
rect 18849 5884 18881 5886
rect 15116 5754 15148 5756
rect 15116 5726 15118 5754
rect 15118 5726 15146 5754
rect 15146 5726 15148 5754
rect 15116 5724 15148 5726
rect 18849 5754 18881 5756
rect 18849 5726 18851 5754
rect 18851 5726 18879 5754
rect 18879 5726 18881 5754
rect 18849 5724 18881 5726
rect 15304 5651 15336 5653
rect 15304 5623 15306 5651
rect 15306 5623 15334 5651
rect 15334 5623 15336 5651
rect 15304 5621 15336 5623
rect 15464 5651 15496 5653
rect 15464 5623 15466 5651
rect 15466 5623 15494 5651
rect 15494 5623 15496 5651
rect 15464 5621 15496 5623
rect 15624 5651 15656 5653
rect 15624 5623 15626 5651
rect 15626 5623 15654 5651
rect 15654 5623 15656 5651
rect 15624 5621 15656 5623
rect 15784 5651 15816 5653
rect 15784 5623 15786 5651
rect 15786 5623 15814 5651
rect 15814 5623 15816 5651
rect 15784 5621 15816 5623
rect 15944 5651 15976 5653
rect 15944 5623 15946 5651
rect 15946 5623 15974 5651
rect 15974 5623 15976 5651
rect 15944 5621 15976 5623
rect 16104 5651 16136 5653
rect 16104 5623 16106 5651
rect 16106 5623 16134 5651
rect 16134 5623 16136 5651
rect 16104 5621 16136 5623
rect 16264 5651 16296 5653
rect 16264 5623 16266 5651
rect 16266 5623 16294 5651
rect 16294 5623 16296 5651
rect 16264 5621 16296 5623
rect 16424 5651 16456 5653
rect 16424 5623 16426 5651
rect 16426 5623 16454 5651
rect 16454 5623 16456 5651
rect 16424 5621 16456 5623
rect 16584 5651 16616 5653
rect 16584 5623 16586 5651
rect 16586 5623 16614 5651
rect 16614 5623 16616 5651
rect 16584 5621 16616 5623
rect 16744 5651 16776 5653
rect 16744 5623 16746 5651
rect 16746 5623 16774 5651
rect 16774 5623 16776 5651
rect 16744 5621 16776 5623
rect 16904 5651 16936 5653
rect 16904 5623 16906 5651
rect 16906 5623 16934 5651
rect 16934 5623 16936 5651
rect 16904 5621 16936 5623
rect 17064 5651 17096 5653
rect 17064 5623 17066 5651
rect 17066 5623 17094 5651
rect 17094 5623 17096 5651
rect 17064 5621 17096 5623
rect 17224 5651 17256 5653
rect 17224 5623 17226 5651
rect 17226 5623 17254 5651
rect 17254 5623 17256 5651
rect 17224 5621 17256 5623
rect 17384 5651 17416 5653
rect 17384 5623 17386 5651
rect 17386 5623 17414 5651
rect 17414 5623 17416 5651
rect 17384 5621 17416 5623
rect 17544 5651 17576 5653
rect 17544 5623 17546 5651
rect 17546 5623 17574 5651
rect 17574 5623 17576 5651
rect 17544 5621 17576 5623
rect 17704 5651 17736 5653
rect 17704 5623 17706 5651
rect 17706 5623 17734 5651
rect 17734 5623 17736 5651
rect 17704 5621 17736 5623
rect 17864 5651 17896 5653
rect 17864 5623 17866 5651
rect 17866 5623 17894 5651
rect 17894 5623 17896 5651
rect 17864 5621 17896 5623
rect 18024 5651 18056 5653
rect 18024 5623 18026 5651
rect 18026 5623 18054 5651
rect 18054 5623 18056 5651
rect 18024 5621 18056 5623
rect 18184 5651 18216 5653
rect 18184 5623 18186 5651
rect 18186 5623 18214 5651
rect 18214 5623 18216 5651
rect 18184 5621 18216 5623
rect 18344 5651 18376 5653
rect 18344 5623 18346 5651
rect 18346 5623 18374 5651
rect 18374 5623 18376 5651
rect 18344 5621 18376 5623
rect 18504 5651 18536 5653
rect 18504 5623 18506 5651
rect 18506 5623 18534 5651
rect 18534 5623 18536 5651
rect 18504 5621 18536 5623
rect 18664 5651 18696 5653
rect 18664 5623 18666 5651
rect 18666 5623 18694 5651
rect 18694 5623 18696 5651
rect 18664 5621 18696 5623
rect 3304 3379 3336 3381
rect 3304 3351 3306 3379
rect 3306 3351 3334 3379
rect 3334 3351 3336 3379
rect 3304 3349 3336 3351
rect 3464 3379 3496 3381
rect 3464 3351 3466 3379
rect 3466 3351 3494 3379
rect 3494 3351 3496 3379
rect 3464 3349 3496 3351
rect 3624 3379 3656 3381
rect 3624 3351 3626 3379
rect 3626 3351 3654 3379
rect 3654 3351 3656 3379
rect 3624 3349 3656 3351
rect 3784 3379 3816 3381
rect 3784 3351 3786 3379
rect 3786 3351 3814 3379
rect 3814 3351 3816 3379
rect 3784 3349 3816 3351
rect 3944 3379 3976 3381
rect 3944 3351 3946 3379
rect 3946 3351 3974 3379
rect 3974 3351 3976 3379
rect 3944 3349 3976 3351
rect 4104 3379 4136 3381
rect 4104 3351 4106 3379
rect 4106 3351 4134 3379
rect 4134 3351 4136 3379
rect 4104 3349 4136 3351
rect 4264 3379 4296 3381
rect 4264 3351 4266 3379
rect 4266 3351 4294 3379
rect 4294 3351 4296 3379
rect 4264 3349 4296 3351
rect 4424 3379 4456 3381
rect 4424 3351 4426 3379
rect 4426 3351 4454 3379
rect 4454 3351 4456 3379
rect 4424 3349 4456 3351
rect 4584 3379 4616 3381
rect 4584 3351 4586 3379
rect 4586 3351 4614 3379
rect 4614 3351 4616 3379
rect 4584 3349 4616 3351
rect 4744 3379 4776 3381
rect 4744 3351 4746 3379
rect 4746 3351 4774 3379
rect 4774 3351 4776 3379
rect 4744 3349 4776 3351
rect 4904 3379 4936 3381
rect 4904 3351 4906 3379
rect 4906 3351 4934 3379
rect 4934 3351 4936 3379
rect 4904 3349 4936 3351
rect 5064 3379 5096 3381
rect 5064 3351 5066 3379
rect 5066 3351 5094 3379
rect 5094 3351 5096 3379
rect 5064 3349 5096 3351
rect 5224 3379 5256 3381
rect 5224 3351 5226 3379
rect 5226 3351 5254 3379
rect 5254 3351 5256 3379
rect 5224 3349 5256 3351
rect 5384 3379 5416 3381
rect 5384 3351 5386 3379
rect 5386 3351 5414 3379
rect 5414 3351 5416 3379
rect 5384 3349 5416 3351
rect 5544 3379 5576 3381
rect 5544 3351 5546 3379
rect 5546 3351 5574 3379
rect 5574 3351 5576 3379
rect 5544 3349 5576 3351
rect 5704 3379 5736 3381
rect 5704 3351 5706 3379
rect 5706 3351 5734 3379
rect 5734 3351 5736 3379
rect 5704 3349 5736 3351
rect 5864 3379 5896 3381
rect 5864 3351 5866 3379
rect 5866 3351 5894 3379
rect 5894 3351 5896 3379
rect 5864 3349 5896 3351
rect 6024 3379 6056 3381
rect 6024 3351 6026 3379
rect 6026 3351 6054 3379
rect 6054 3351 6056 3379
rect 6024 3349 6056 3351
rect 6184 3379 6216 3381
rect 6184 3351 6186 3379
rect 6186 3351 6214 3379
rect 6214 3351 6216 3379
rect 6184 3349 6216 3351
rect 6344 3379 6376 3381
rect 6344 3351 6346 3379
rect 6346 3351 6374 3379
rect 6374 3351 6376 3379
rect 6344 3349 6376 3351
rect 6504 3379 6536 3381
rect 6504 3351 6506 3379
rect 6506 3351 6534 3379
rect 6534 3351 6536 3379
rect 6504 3349 6536 3351
rect 6664 3379 6696 3381
rect 6664 3351 6666 3379
rect 6666 3351 6694 3379
rect 6694 3351 6696 3379
rect 6664 3349 6696 3351
rect 3116 3274 3148 3276
rect 3116 3246 3118 3274
rect 3118 3246 3146 3274
rect 3146 3246 3148 3274
rect 3116 3244 3148 3246
rect 6849 3274 6881 3276
rect 6849 3246 6851 3274
rect 6851 3246 6879 3274
rect 6879 3246 6881 3274
rect 6849 3244 6881 3246
rect 3116 3114 3148 3116
rect 3116 3086 3118 3114
rect 3118 3086 3146 3114
rect 3146 3086 3148 3114
rect 3116 3084 3148 3086
rect 3116 2954 3148 2956
rect 3116 2926 3118 2954
rect 3118 2926 3146 2954
rect 3146 2926 3148 2954
rect 3116 2924 3148 2926
rect 3116 2794 3148 2796
rect 3116 2766 3118 2794
rect 3118 2766 3146 2794
rect 3146 2766 3148 2794
rect 3116 2764 3148 2766
rect 3116 2634 3148 2636
rect 3116 2606 3118 2634
rect 3118 2606 3146 2634
rect 3146 2606 3148 2634
rect 3116 2604 3148 2606
rect 3116 2474 3148 2476
rect 3116 2446 3118 2474
rect 3118 2446 3146 2474
rect 3146 2446 3148 2474
rect 3116 2444 3148 2446
rect 3116 2314 3148 2316
rect 3116 2286 3118 2314
rect 3118 2286 3146 2314
rect 3146 2286 3148 2314
rect 3116 2284 3148 2286
rect 3116 2154 3148 2156
rect 3116 2126 3118 2154
rect 3118 2126 3146 2154
rect 3146 2126 3148 2154
rect 3116 2124 3148 2126
rect 3116 1994 3148 1996
rect 3116 1966 3118 1994
rect 3118 1966 3146 1994
rect 3146 1966 3148 1994
rect 3116 1964 3148 1966
rect 3116 1834 3148 1836
rect 3116 1806 3118 1834
rect 3118 1806 3146 1834
rect 3146 1806 3148 1834
rect 3116 1804 3148 1806
rect 3116 1674 3148 1676
rect 3116 1646 3118 1674
rect 3118 1646 3146 1674
rect 3146 1646 3148 1674
rect 3116 1644 3148 1646
rect 3116 1514 3148 1516
rect 3116 1486 3118 1514
rect 3118 1486 3146 1514
rect 3146 1486 3148 1514
rect 3116 1484 3148 1486
rect 3116 1354 3148 1356
rect 3116 1326 3118 1354
rect 3118 1326 3146 1354
rect 3146 1326 3148 1354
rect 3116 1324 3148 1326
rect 3116 1194 3148 1196
rect 3116 1166 3118 1194
rect 3118 1166 3146 1194
rect 3146 1166 3148 1194
rect 3116 1164 3148 1166
rect 3116 1034 3148 1036
rect 3116 1006 3118 1034
rect 3118 1006 3146 1034
rect 3146 1006 3148 1034
rect 3116 1004 3148 1006
rect 3116 874 3148 876
rect 3116 846 3118 874
rect 3118 846 3146 874
rect 3146 846 3148 874
rect 3116 844 3148 846
rect 3116 714 3148 716
rect 3116 686 3118 714
rect 3118 686 3146 714
rect 3146 686 3148 714
rect 3116 684 3148 686
rect 3116 554 3148 556
rect 3116 526 3118 554
rect 3118 526 3146 554
rect 3146 526 3148 554
rect 3116 524 3148 526
rect 3116 394 3148 396
rect 3116 366 3118 394
rect 3118 366 3146 394
rect 3146 366 3148 394
rect 3116 364 3148 366
rect 3116 234 3148 236
rect 3116 206 3118 234
rect 3118 206 3146 234
rect 3146 206 3148 234
rect 3116 204 3148 206
rect 3116 74 3148 76
rect 3116 46 3118 74
rect 3118 46 3146 74
rect 3146 46 3148 74
rect 3116 44 3148 46
rect 3116 -86 3148 -84
rect 3116 -114 3118 -86
rect 3118 -114 3146 -86
rect 3146 -114 3148 -86
rect 3116 -116 3148 -114
rect 6849 3114 6881 3116
rect 6849 3086 6851 3114
rect 6851 3086 6879 3114
rect 6879 3086 6881 3114
rect 6849 3084 6881 3086
rect 6849 2954 6881 2956
rect 6849 2926 6851 2954
rect 6851 2926 6879 2954
rect 6879 2926 6881 2954
rect 6849 2924 6881 2926
rect 6849 2794 6881 2796
rect 6849 2766 6851 2794
rect 6851 2766 6879 2794
rect 6879 2766 6881 2794
rect 6849 2764 6881 2766
rect 6849 2634 6881 2636
rect 6849 2606 6851 2634
rect 6851 2606 6879 2634
rect 6879 2606 6881 2634
rect 6849 2604 6881 2606
rect 6849 2474 6881 2476
rect 6849 2446 6851 2474
rect 6851 2446 6879 2474
rect 6879 2446 6881 2474
rect 6849 2444 6881 2446
rect 6849 2314 6881 2316
rect 6849 2286 6851 2314
rect 6851 2286 6879 2314
rect 6879 2286 6881 2314
rect 6849 2284 6881 2286
rect 6849 2154 6881 2156
rect 6849 2126 6851 2154
rect 6851 2126 6879 2154
rect 6879 2126 6881 2154
rect 6849 2124 6881 2126
rect 6849 1994 6881 1996
rect 6849 1966 6851 1994
rect 6851 1966 6879 1994
rect 6879 1966 6881 1994
rect 6849 1964 6881 1966
rect 6849 1834 6881 1836
rect 6849 1806 6851 1834
rect 6851 1806 6879 1834
rect 6879 1806 6881 1834
rect 6849 1804 6881 1806
rect 6849 1674 6881 1676
rect 6849 1646 6851 1674
rect 6851 1646 6879 1674
rect 6879 1646 6881 1674
rect 6849 1644 6881 1646
rect 6849 1514 6881 1516
rect 6849 1486 6851 1514
rect 6851 1486 6879 1514
rect 6879 1486 6881 1514
rect 6849 1484 6881 1486
rect 6849 1354 6881 1356
rect 6849 1326 6851 1354
rect 6851 1326 6879 1354
rect 6879 1326 6881 1354
rect 6849 1324 6881 1326
rect 6849 1194 6881 1196
rect 6849 1166 6851 1194
rect 6851 1166 6879 1194
rect 6879 1166 6881 1194
rect 6849 1164 6881 1166
rect 6849 1034 6881 1036
rect 6849 1006 6851 1034
rect 6851 1006 6879 1034
rect 6879 1006 6881 1034
rect 6849 1004 6881 1006
rect 6849 874 6881 876
rect 6849 846 6851 874
rect 6851 846 6879 874
rect 6879 846 6881 874
rect 6849 844 6881 846
rect 6849 714 6881 716
rect 6849 686 6851 714
rect 6851 686 6879 714
rect 6879 686 6881 714
rect 6849 684 6881 686
rect 6849 554 6881 556
rect 6849 526 6851 554
rect 6851 526 6879 554
rect 6879 526 6881 554
rect 6849 524 6881 526
rect 6849 394 6881 396
rect 6849 366 6851 394
rect 6851 366 6879 394
rect 6879 366 6881 394
rect 6849 364 6881 366
rect 6849 234 6881 236
rect 6849 206 6851 234
rect 6851 206 6879 234
rect 6879 206 6881 234
rect 6849 204 6881 206
rect 6849 74 6881 76
rect 6849 46 6851 74
rect 6851 46 6879 74
rect 6879 46 6881 74
rect 6849 44 6881 46
rect 6849 -86 6881 -84
rect 6849 -114 6851 -86
rect 6851 -114 6879 -86
rect 6879 -114 6881 -86
rect 6849 -116 6881 -114
rect 3116 -246 3148 -244
rect 3116 -274 3118 -246
rect 3118 -274 3146 -246
rect 3146 -274 3148 -246
rect 3116 -276 3148 -274
rect 6849 -246 6881 -244
rect 6849 -274 6851 -246
rect 6851 -274 6879 -246
rect 6879 -274 6881 -246
rect 6849 -276 6881 -274
rect 3304 -349 3336 -347
rect 3304 -377 3306 -349
rect 3306 -377 3334 -349
rect 3334 -377 3336 -349
rect 3304 -379 3336 -377
rect 3464 -349 3496 -347
rect 3464 -377 3466 -349
rect 3466 -377 3494 -349
rect 3494 -377 3496 -349
rect 3464 -379 3496 -377
rect 3624 -349 3656 -347
rect 3624 -377 3626 -349
rect 3626 -377 3654 -349
rect 3654 -377 3656 -349
rect 3624 -379 3656 -377
rect 3784 -349 3816 -347
rect 3784 -377 3786 -349
rect 3786 -377 3814 -349
rect 3814 -377 3816 -349
rect 3784 -379 3816 -377
rect 3944 -349 3976 -347
rect 3944 -377 3946 -349
rect 3946 -377 3974 -349
rect 3974 -377 3976 -349
rect 3944 -379 3976 -377
rect 4104 -349 4136 -347
rect 4104 -377 4106 -349
rect 4106 -377 4134 -349
rect 4134 -377 4136 -349
rect 4104 -379 4136 -377
rect 4264 -349 4296 -347
rect 4264 -377 4266 -349
rect 4266 -377 4294 -349
rect 4294 -377 4296 -349
rect 4264 -379 4296 -377
rect 4424 -349 4456 -347
rect 4424 -377 4426 -349
rect 4426 -377 4454 -349
rect 4454 -377 4456 -349
rect 4424 -379 4456 -377
rect 4584 -349 4616 -347
rect 4584 -377 4586 -349
rect 4586 -377 4614 -349
rect 4614 -377 4616 -349
rect 4584 -379 4616 -377
rect 4744 -349 4776 -347
rect 4744 -377 4746 -349
rect 4746 -377 4774 -349
rect 4774 -377 4776 -349
rect 4744 -379 4776 -377
rect 4904 -349 4936 -347
rect 4904 -377 4906 -349
rect 4906 -377 4934 -349
rect 4934 -377 4936 -349
rect 4904 -379 4936 -377
rect 5064 -349 5096 -347
rect 5064 -377 5066 -349
rect 5066 -377 5094 -349
rect 5094 -377 5096 -349
rect 5064 -379 5096 -377
rect 5224 -349 5256 -347
rect 5224 -377 5226 -349
rect 5226 -377 5254 -349
rect 5254 -377 5256 -349
rect 5224 -379 5256 -377
rect 5384 -349 5416 -347
rect 5384 -377 5386 -349
rect 5386 -377 5414 -349
rect 5414 -377 5416 -349
rect 5384 -379 5416 -377
rect 5544 -349 5576 -347
rect 5544 -377 5546 -349
rect 5546 -377 5574 -349
rect 5574 -377 5576 -349
rect 5544 -379 5576 -377
rect 5704 -349 5736 -347
rect 5704 -377 5706 -349
rect 5706 -377 5734 -349
rect 5734 -377 5736 -349
rect 5704 -379 5736 -377
rect 5864 -349 5896 -347
rect 5864 -377 5866 -349
rect 5866 -377 5894 -349
rect 5894 -377 5896 -349
rect 5864 -379 5896 -377
rect 6024 -349 6056 -347
rect 6024 -377 6026 -349
rect 6026 -377 6054 -349
rect 6054 -377 6056 -349
rect 6024 -379 6056 -377
rect 6184 -349 6216 -347
rect 6184 -377 6186 -349
rect 6186 -377 6214 -349
rect 6214 -377 6216 -349
rect 6184 -379 6216 -377
rect 6344 -349 6376 -347
rect 6344 -377 6346 -349
rect 6346 -377 6374 -349
rect 6374 -377 6376 -349
rect 6344 -379 6376 -377
rect 6504 -349 6536 -347
rect 6504 -377 6506 -349
rect 6506 -377 6534 -349
rect 6534 -377 6536 -349
rect 6504 -379 6536 -377
rect 6664 -349 6696 -347
rect 6664 -377 6666 -349
rect 6666 -377 6694 -349
rect 6694 -377 6696 -349
rect 6664 -379 6696 -377
rect 9304 3379 9336 3381
rect 9304 3351 9306 3379
rect 9306 3351 9334 3379
rect 9334 3351 9336 3379
rect 9304 3349 9336 3351
rect 9464 3379 9496 3381
rect 9464 3351 9466 3379
rect 9466 3351 9494 3379
rect 9494 3351 9496 3379
rect 9464 3349 9496 3351
rect 9624 3379 9656 3381
rect 9624 3351 9626 3379
rect 9626 3351 9654 3379
rect 9654 3351 9656 3379
rect 9624 3349 9656 3351
rect 9784 3379 9816 3381
rect 9784 3351 9786 3379
rect 9786 3351 9814 3379
rect 9814 3351 9816 3379
rect 9784 3349 9816 3351
rect 9944 3379 9976 3381
rect 9944 3351 9946 3379
rect 9946 3351 9974 3379
rect 9974 3351 9976 3379
rect 9944 3349 9976 3351
rect 10104 3379 10136 3381
rect 10104 3351 10106 3379
rect 10106 3351 10134 3379
rect 10134 3351 10136 3379
rect 10104 3349 10136 3351
rect 10264 3379 10296 3381
rect 10264 3351 10266 3379
rect 10266 3351 10294 3379
rect 10294 3351 10296 3379
rect 10264 3349 10296 3351
rect 10424 3379 10456 3381
rect 10424 3351 10426 3379
rect 10426 3351 10454 3379
rect 10454 3351 10456 3379
rect 10424 3349 10456 3351
rect 10584 3379 10616 3381
rect 10584 3351 10586 3379
rect 10586 3351 10614 3379
rect 10614 3351 10616 3379
rect 10584 3349 10616 3351
rect 10744 3379 10776 3381
rect 10744 3351 10746 3379
rect 10746 3351 10774 3379
rect 10774 3351 10776 3379
rect 10744 3349 10776 3351
rect 10904 3379 10936 3381
rect 10904 3351 10906 3379
rect 10906 3351 10934 3379
rect 10934 3351 10936 3379
rect 10904 3349 10936 3351
rect 11064 3379 11096 3381
rect 11064 3351 11066 3379
rect 11066 3351 11094 3379
rect 11094 3351 11096 3379
rect 11064 3349 11096 3351
rect 11224 3379 11256 3381
rect 11224 3351 11226 3379
rect 11226 3351 11254 3379
rect 11254 3351 11256 3379
rect 11224 3349 11256 3351
rect 11384 3379 11416 3381
rect 11384 3351 11386 3379
rect 11386 3351 11414 3379
rect 11414 3351 11416 3379
rect 11384 3349 11416 3351
rect 11544 3379 11576 3381
rect 11544 3351 11546 3379
rect 11546 3351 11574 3379
rect 11574 3351 11576 3379
rect 11544 3349 11576 3351
rect 11704 3379 11736 3381
rect 11704 3351 11706 3379
rect 11706 3351 11734 3379
rect 11734 3351 11736 3379
rect 11704 3349 11736 3351
rect 11864 3379 11896 3381
rect 11864 3351 11866 3379
rect 11866 3351 11894 3379
rect 11894 3351 11896 3379
rect 11864 3349 11896 3351
rect 12024 3379 12056 3381
rect 12024 3351 12026 3379
rect 12026 3351 12054 3379
rect 12054 3351 12056 3379
rect 12024 3349 12056 3351
rect 12184 3379 12216 3381
rect 12184 3351 12186 3379
rect 12186 3351 12214 3379
rect 12214 3351 12216 3379
rect 12184 3349 12216 3351
rect 12344 3379 12376 3381
rect 12344 3351 12346 3379
rect 12346 3351 12374 3379
rect 12374 3351 12376 3379
rect 12344 3349 12376 3351
rect 12504 3379 12536 3381
rect 12504 3351 12506 3379
rect 12506 3351 12534 3379
rect 12534 3351 12536 3379
rect 12504 3349 12536 3351
rect 12664 3379 12696 3381
rect 12664 3351 12666 3379
rect 12666 3351 12694 3379
rect 12694 3351 12696 3379
rect 12664 3349 12696 3351
rect 9116 3274 9148 3276
rect 9116 3246 9118 3274
rect 9118 3246 9146 3274
rect 9146 3246 9148 3274
rect 9116 3244 9148 3246
rect 12849 3274 12881 3276
rect 12849 3246 12851 3274
rect 12851 3246 12879 3274
rect 12879 3246 12881 3274
rect 12849 3244 12881 3246
rect 9116 3114 9148 3116
rect 9116 3086 9118 3114
rect 9118 3086 9146 3114
rect 9146 3086 9148 3114
rect 9116 3084 9148 3086
rect 9116 2954 9148 2956
rect 9116 2926 9118 2954
rect 9118 2926 9146 2954
rect 9146 2926 9148 2954
rect 9116 2924 9148 2926
rect 9116 2794 9148 2796
rect 9116 2766 9118 2794
rect 9118 2766 9146 2794
rect 9146 2766 9148 2794
rect 9116 2764 9148 2766
rect 9116 2634 9148 2636
rect 9116 2606 9118 2634
rect 9118 2606 9146 2634
rect 9146 2606 9148 2634
rect 9116 2604 9148 2606
rect 9116 2474 9148 2476
rect 9116 2446 9118 2474
rect 9118 2446 9146 2474
rect 9146 2446 9148 2474
rect 9116 2444 9148 2446
rect 9116 2314 9148 2316
rect 9116 2286 9118 2314
rect 9118 2286 9146 2314
rect 9146 2286 9148 2314
rect 9116 2284 9148 2286
rect 9116 2154 9148 2156
rect 9116 2126 9118 2154
rect 9118 2126 9146 2154
rect 9146 2126 9148 2154
rect 9116 2124 9148 2126
rect 9116 1994 9148 1996
rect 9116 1966 9118 1994
rect 9118 1966 9146 1994
rect 9146 1966 9148 1994
rect 9116 1964 9148 1966
rect 9116 1834 9148 1836
rect 9116 1806 9118 1834
rect 9118 1806 9146 1834
rect 9146 1806 9148 1834
rect 9116 1804 9148 1806
rect 9116 1674 9148 1676
rect 9116 1646 9118 1674
rect 9118 1646 9146 1674
rect 9146 1646 9148 1674
rect 9116 1644 9148 1646
rect 9116 1514 9148 1516
rect 9116 1486 9118 1514
rect 9118 1486 9146 1514
rect 9146 1486 9148 1514
rect 9116 1484 9148 1486
rect 9116 1354 9148 1356
rect 9116 1326 9118 1354
rect 9118 1326 9146 1354
rect 9146 1326 9148 1354
rect 9116 1324 9148 1326
rect 9116 1194 9148 1196
rect 9116 1166 9118 1194
rect 9118 1166 9146 1194
rect 9146 1166 9148 1194
rect 9116 1164 9148 1166
rect 9116 1034 9148 1036
rect 9116 1006 9118 1034
rect 9118 1006 9146 1034
rect 9146 1006 9148 1034
rect 9116 1004 9148 1006
rect 9116 874 9148 876
rect 9116 846 9118 874
rect 9118 846 9146 874
rect 9146 846 9148 874
rect 9116 844 9148 846
rect 9116 714 9148 716
rect 9116 686 9118 714
rect 9118 686 9146 714
rect 9146 686 9148 714
rect 9116 684 9148 686
rect 9116 554 9148 556
rect 9116 526 9118 554
rect 9118 526 9146 554
rect 9146 526 9148 554
rect 9116 524 9148 526
rect 9116 394 9148 396
rect 9116 366 9118 394
rect 9118 366 9146 394
rect 9146 366 9148 394
rect 9116 364 9148 366
rect 9116 234 9148 236
rect 9116 206 9118 234
rect 9118 206 9146 234
rect 9146 206 9148 234
rect 9116 204 9148 206
rect 9116 74 9148 76
rect 9116 46 9118 74
rect 9118 46 9146 74
rect 9146 46 9148 74
rect 9116 44 9148 46
rect 9116 -86 9148 -84
rect 9116 -114 9118 -86
rect 9118 -114 9146 -86
rect 9146 -114 9148 -86
rect 9116 -116 9148 -114
rect 12849 3114 12881 3116
rect 12849 3086 12851 3114
rect 12851 3086 12879 3114
rect 12879 3086 12881 3114
rect 12849 3084 12881 3086
rect 12849 2954 12881 2956
rect 12849 2926 12851 2954
rect 12851 2926 12879 2954
rect 12879 2926 12881 2954
rect 12849 2924 12881 2926
rect 12849 2794 12881 2796
rect 12849 2766 12851 2794
rect 12851 2766 12879 2794
rect 12879 2766 12881 2794
rect 12849 2764 12881 2766
rect 12849 2634 12881 2636
rect 12849 2606 12851 2634
rect 12851 2606 12879 2634
rect 12879 2606 12881 2634
rect 12849 2604 12881 2606
rect 12849 2474 12881 2476
rect 12849 2446 12851 2474
rect 12851 2446 12879 2474
rect 12879 2446 12881 2474
rect 12849 2444 12881 2446
rect 12849 2314 12881 2316
rect 12849 2286 12851 2314
rect 12851 2286 12879 2314
rect 12879 2286 12881 2314
rect 12849 2284 12881 2286
rect 12849 2154 12881 2156
rect 12849 2126 12851 2154
rect 12851 2126 12879 2154
rect 12879 2126 12881 2154
rect 12849 2124 12881 2126
rect 12849 1994 12881 1996
rect 12849 1966 12851 1994
rect 12851 1966 12879 1994
rect 12879 1966 12881 1994
rect 12849 1964 12881 1966
rect 12849 1834 12881 1836
rect 12849 1806 12851 1834
rect 12851 1806 12879 1834
rect 12879 1806 12881 1834
rect 12849 1804 12881 1806
rect 15304 3379 15336 3381
rect 15304 3351 15306 3379
rect 15306 3351 15334 3379
rect 15334 3351 15336 3379
rect 15304 3349 15336 3351
rect 15464 3379 15496 3381
rect 15464 3351 15466 3379
rect 15466 3351 15494 3379
rect 15494 3351 15496 3379
rect 15464 3349 15496 3351
rect 15624 3379 15656 3381
rect 15624 3351 15626 3379
rect 15626 3351 15654 3379
rect 15654 3351 15656 3379
rect 15624 3349 15656 3351
rect 15784 3379 15816 3381
rect 15784 3351 15786 3379
rect 15786 3351 15814 3379
rect 15814 3351 15816 3379
rect 15784 3349 15816 3351
rect 15944 3379 15976 3381
rect 15944 3351 15946 3379
rect 15946 3351 15974 3379
rect 15974 3351 15976 3379
rect 15944 3349 15976 3351
rect 16104 3379 16136 3381
rect 16104 3351 16106 3379
rect 16106 3351 16134 3379
rect 16134 3351 16136 3379
rect 16104 3349 16136 3351
rect 16264 3379 16296 3381
rect 16264 3351 16266 3379
rect 16266 3351 16294 3379
rect 16294 3351 16296 3379
rect 16264 3349 16296 3351
rect 16424 3379 16456 3381
rect 16424 3351 16426 3379
rect 16426 3351 16454 3379
rect 16454 3351 16456 3379
rect 16424 3349 16456 3351
rect 16584 3379 16616 3381
rect 16584 3351 16586 3379
rect 16586 3351 16614 3379
rect 16614 3351 16616 3379
rect 16584 3349 16616 3351
rect 16744 3379 16776 3381
rect 16744 3351 16746 3379
rect 16746 3351 16774 3379
rect 16774 3351 16776 3379
rect 16744 3349 16776 3351
rect 16904 3379 16936 3381
rect 16904 3351 16906 3379
rect 16906 3351 16934 3379
rect 16934 3351 16936 3379
rect 16904 3349 16936 3351
rect 17064 3379 17096 3381
rect 17064 3351 17066 3379
rect 17066 3351 17094 3379
rect 17094 3351 17096 3379
rect 17064 3349 17096 3351
rect 17224 3379 17256 3381
rect 17224 3351 17226 3379
rect 17226 3351 17254 3379
rect 17254 3351 17256 3379
rect 17224 3349 17256 3351
rect 17384 3379 17416 3381
rect 17384 3351 17386 3379
rect 17386 3351 17414 3379
rect 17414 3351 17416 3379
rect 17384 3349 17416 3351
rect 17544 3379 17576 3381
rect 17544 3351 17546 3379
rect 17546 3351 17574 3379
rect 17574 3351 17576 3379
rect 17544 3349 17576 3351
rect 17704 3379 17736 3381
rect 17704 3351 17706 3379
rect 17706 3351 17734 3379
rect 17734 3351 17736 3379
rect 17704 3349 17736 3351
rect 17864 3379 17896 3381
rect 17864 3351 17866 3379
rect 17866 3351 17894 3379
rect 17894 3351 17896 3379
rect 17864 3349 17896 3351
rect 18024 3379 18056 3381
rect 18024 3351 18026 3379
rect 18026 3351 18054 3379
rect 18054 3351 18056 3379
rect 18024 3349 18056 3351
rect 18184 3379 18216 3381
rect 18184 3351 18186 3379
rect 18186 3351 18214 3379
rect 18214 3351 18216 3379
rect 18184 3349 18216 3351
rect 18344 3379 18376 3381
rect 18344 3351 18346 3379
rect 18346 3351 18374 3379
rect 18374 3351 18376 3379
rect 18344 3349 18376 3351
rect 18504 3379 18536 3381
rect 18504 3351 18506 3379
rect 18506 3351 18534 3379
rect 18534 3351 18536 3379
rect 18504 3349 18536 3351
rect 18664 3379 18696 3381
rect 18664 3351 18666 3379
rect 18666 3351 18694 3379
rect 18694 3351 18696 3379
rect 18664 3349 18696 3351
rect 15116 3274 15148 3276
rect 15116 3246 15118 3274
rect 15118 3246 15146 3274
rect 15146 3246 15148 3274
rect 15116 3244 15148 3246
rect 18849 3274 18881 3276
rect 18849 3246 18851 3274
rect 18851 3246 18879 3274
rect 18879 3246 18881 3274
rect 18849 3244 18881 3246
rect 15116 3114 15148 3116
rect 15116 3086 15118 3114
rect 15118 3086 15146 3114
rect 15146 3086 15148 3114
rect 15116 3084 15148 3086
rect 15116 2954 15148 2956
rect 15116 2926 15118 2954
rect 15118 2926 15146 2954
rect 15146 2926 15148 2954
rect 15116 2924 15148 2926
rect 15116 2794 15148 2796
rect 15116 2766 15118 2794
rect 15118 2766 15146 2794
rect 15146 2766 15148 2794
rect 15116 2764 15148 2766
rect 15116 2634 15148 2636
rect 15116 2606 15118 2634
rect 15118 2606 15146 2634
rect 15146 2606 15148 2634
rect 15116 2604 15148 2606
rect 15116 2474 15148 2476
rect 15116 2446 15118 2474
rect 15118 2446 15146 2474
rect 15146 2446 15148 2474
rect 15116 2444 15148 2446
rect 15116 2314 15148 2316
rect 15116 2286 15118 2314
rect 15118 2286 15146 2314
rect 15146 2286 15148 2314
rect 15116 2284 15148 2286
rect 15116 2154 15148 2156
rect 15116 2126 15118 2154
rect 15118 2126 15146 2154
rect 15146 2126 15148 2154
rect 15116 2124 15148 2126
rect 15116 1994 15148 1996
rect 15116 1966 15118 1994
rect 15118 1966 15146 1994
rect 15146 1966 15148 1994
rect 15116 1964 15148 1966
rect 12849 1674 12881 1676
rect 12849 1646 12851 1674
rect 12851 1646 12879 1674
rect 12879 1646 12881 1674
rect 12849 1644 12881 1646
rect 12849 1514 12881 1516
rect 12849 1486 12851 1514
rect 12851 1486 12879 1514
rect 12879 1486 12881 1514
rect 12849 1484 12881 1486
rect 12849 1354 12881 1356
rect 12849 1326 12851 1354
rect 12851 1326 12879 1354
rect 12879 1326 12881 1354
rect 12849 1324 12881 1326
rect 12849 1194 12881 1196
rect 12849 1166 12851 1194
rect 12851 1166 12879 1194
rect 12879 1166 12881 1194
rect 12849 1164 12881 1166
rect 12849 1034 12881 1036
rect 12849 1006 12851 1034
rect 12851 1006 12879 1034
rect 12879 1006 12881 1034
rect 12849 1004 12881 1006
rect 12849 874 12881 876
rect 12849 846 12851 874
rect 12851 846 12879 874
rect 12879 846 12881 874
rect 12849 844 12881 846
rect 12849 714 12881 716
rect 12849 686 12851 714
rect 12851 686 12879 714
rect 12879 686 12881 714
rect 12849 684 12881 686
rect 12849 554 12881 556
rect 12849 526 12851 554
rect 12851 526 12879 554
rect 12879 526 12881 554
rect 12849 524 12881 526
rect 12849 394 12881 396
rect 12849 366 12851 394
rect 12851 366 12879 394
rect 12879 366 12881 394
rect 12849 364 12881 366
rect 12849 234 12881 236
rect 12849 206 12851 234
rect 12851 206 12879 234
rect 12879 206 12881 234
rect 12849 204 12881 206
rect 12849 74 12881 76
rect 12849 46 12851 74
rect 12851 46 12879 74
rect 12879 46 12881 74
rect 12849 44 12881 46
rect 12849 -86 12881 -84
rect 12849 -114 12851 -86
rect 12851 -114 12879 -86
rect 12879 -114 12881 -86
rect 12849 -116 12881 -114
rect 9116 -246 9148 -244
rect 9116 -274 9118 -246
rect 9118 -274 9146 -246
rect 9146 -274 9148 -246
rect 9116 -276 9148 -274
rect 12849 -246 12881 -244
rect 12849 -274 12851 -246
rect 12851 -274 12879 -246
rect 12879 -274 12881 -246
rect 12849 -276 12881 -274
rect 9304 -349 9336 -347
rect 9304 -377 9306 -349
rect 9306 -377 9334 -349
rect 9334 -377 9336 -349
rect 9304 -379 9336 -377
rect 9464 -349 9496 -347
rect 9464 -377 9466 -349
rect 9466 -377 9494 -349
rect 9494 -377 9496 -349
rect 9464 -379 9496 -377
rect 9624 -349 9656 -347
rect 9624 -377 9626 -349
rect 9626 -377 9654 -349
rect 9654 -377 9656 -349
rect 9624 -379 9656 -377
rect 9784 -349 9816 -347
rect 9784 -377 9786 -349
rect 9786 -377 9814 -349
rect 9814 -377 9816 -349
rect 9784 -379 9816 -377
rect 9944 -349 9976 -347
rect 9944 -377 9946 -349
rect 9946 -377 9974 -349
rect 9974 -377 9976 -349
rect 9944 -379 9976 -377
rect 10104 -349 10136 -347
rect 10104 -377 10106 -349
rect 10106 -377 10134 -349
rect 10134 -377 10136 -349
rect 10104 -379 10136 -377
rect 10264 -349 10296 -347
rect 10264 -377 10266 -349
rect 10266 -377 10294 -349
rect 10294 -377 10296 -349
rect 10264 -379 10296 -377
rect 10424 -349 10456 -347
rect 10424 -377 10426 -349
rect 10426 -377 10454 -349
rect 10454 -377 10456 -349
rect 10424 -379 10456 -377
rect 10584 -349 10616 -347
rect 10584 -377 10586 -349
rect 10586 -377 10614 -349
rect 10614 -377 10616 -349
rect 10584 -379 10616 -377
rect 10744 -349 10776 -347
rect 10744 -377 10746 -349
rect 10746 -377 10774 -349
rect 10774 -377 10776 -349
rect 10744 -379 10776 -377
rect 10904 -349 10936 -347
rect 10904 -377 10906 -349
rect 10906 -377 10934 -349
rect 10934 -377 10936 -349
rect 10904 -379 10936 -377
rect 11064 -349 11096 -347
rect 11064 -377 11066 -349
rect 11066 -377 11094 -349
rect 11094 -377 11096 -349
rect 11064 -379 11096 -377
rect 11224 -349 11256 -347
rect 11224 -377 11226 -349
rect 11226 -377 11254 -349
rect 11254 -377 11256 -349
rect 11224 -379 11256 -377
rect 11384 -349 11416 -347
rect 11384 -377 11386 -349
rect 11386 -377 11414 -349
rect 11414 -377 11416 -349
rect 11384 -379 11416 -377
rect 11544 -349 11576 -347
rect 11544 -377 11546 -349
rect 11546 -377 11574 -349
rect 11574 -377 11576 -349
rect 11544 -379 11576 -377
rect 11704 -349 11736 -347
rect 11704 -377 11706 -349
rect 11706 -377 11734 -349
rect 11734 -377 11736 -349
rect 11704 -379 11736 -377
rect 11864 -349 11896 -347
rect 11864 -377 11866 -349
rect 11866 -377 11894 -349
rect 11894 -377 11896 -349
rect 11864 -379 11896 -377
rect 12024 -349 12056 -347
rect 12024 -377 12026 -349
rect 12026 -377 12054 -349
rect 12054 -377 12056 -349
rect 12024 -379 12056 -377
rect 12184 -349 12216 -347
rect 12184 -377 12186 -349
rect 12186 -377 12214 -349
rect 12214 -377 12216 -349
rect 12184 -379 12216 -377
rect 12344 -349 12376 -347
rect 12344 -377 12346 -349
rect 12346 -377 12374 -349
rect 12374 -377 12376 -349
rect 12344 -379 12376 -377
rect 12504 -349 12536 -347
rect 12504 -377 12506 -349
rect 12506 -377 12534 -349
rect 12534 -377 12536 -349
rect 12504 -379 12536 -377
rect 12664 -349 12696 -347
rect 12664 -377 12666 -349
rect 12666 -377 12694 -349
rect 12694 -377 12696 -349
rect 12664 -379 12696 -377
rect 15116 1834 15148 1836
rect 15116 1806 15118 1834
rect 15118 1806 15146 1834
rect 15146 1806 15148 1834
rect 15116 1804 15148 1806
rect 15116 1674 15148 1676
rect 15116 1646 15118 1674
rect 15118 1646 15146 1674
rect 15146 1646 15148 1674
rect 15116 1644 15148 1646
rect 15116 1514 15148 1516
rect 15116 1486 15118 1514
rect 15118 1486 15146 1514
rect 15146 1486 15148 1514
rect 15116 1484 15148 1486
rect 15116 1354 15148 1356
rect 15116 1326 15118 1354
rect 15118 1326 15146 1354
rect 15146 1326 15148 1354
rect 15116 1324 15148 1326
rect 15116 1194 15148 1196
rect 15116 1166 15118 1194
rect 15118 1166 15146 1194
rect 15146 1166 15148 1194
rect 15116 1164 15148 1166
rect 15116 1034 15148 1036
rect 15116 1006 15118 1034
rect 15118 1006 15146 1034
rect 15146 1006 15148 1034
rect 15116 1004 15148 1006
rect 15116 874 15148 876
rect 15116 846 15118 874
rect 15118 846 15146 874
rect 15146 846 15148 874
rect 15116 844 15148 846
rect 15116 714 15148 716
rect 15116 686 15118 714
rect 15118 686 15146 714
rect 15146 686 15148 714
rect 15116 684 15148 686
rect 15116 554 15148 556
rect 15116 526 15118 554
rect 15118 526 15146 554
rect 15146 526 15148 554
rect 15116 524 15148 526
rect 15116 394 15148 396
rect 15116 366 15118 394
rect 15118 366 15146 394
rect 15146 366 15148 394
rect 15116 364 15148 366
rect 15116 234 15148 236
rect 15116 206 15118 234
rect 15118 206 15146 234
rect 15146 206 15148 234
rect 15116 204 15148 206
rect 15116 74 15148 76
rect 15116 46 15118 74
rect 15118 46 15146 74
rect 15146 46 15148 74
rect 15116 44 15148 46
rect 15116 -86 15148 -84
rect 15116 -114 15118 -86
rect 15118 -114 15146 -86
rect 15146 -114 15148 -86
rect 15116 -116 15148 -114
rect 18849 3114 18881 3116
rect 18849 3086 18851 3114
rect 18851 3086 18879 3114
rect 18879 3086 18881 3114
rect 18849 3084 18881 3086
rect 18849 2954 18881 2956
rect 18849 2926 18851 2954
rect 18851 2926 18879 2954
rect 18879 2926 18881 2954
rect 18849 2924 18881 2926
rect 18849 2794 18881 2796
rect 18849 2766 18851 2794
rect 18851 2766 18879 2794
rect 18879 2766 18881 2794
rect 18849 2764 18881 2766
rect 18849 2634 18881 2636
rect 18849 2606 18851 2634
rect 18851 2606 18879 2634
rect 18879 2606 18881 2634
rect 18849 2604 18881 2606
rect 18849 2474 18881 2476
rect 18849 2446 18851 2474
rect 18851 2446 18879 2474
rect 18879 2446 18881 2474
rect 18849 2444 18881 2446
rect 18849 2314 18881 2316
rect 18849 2286 18851 2314
rect 18851 2286 18879 2314
rect 18879 2286 18881 2314
rect 18849 2284 18881 2286
rect 18849 2154 18881 2156
rect 18849 2126 18851 2154
rect 18851 2126 18879 2154
rect 18879 2126 18881 2154
rect 18849 2124 18881 2126
rect 18849 1994 18881 1996
rect 18849 1966 18851 1994
rect 18851 1966 18879 1994
rect 18879 1966 18881 1994
rect 18849 1964 18881 1966
rect 18849 1834 18881 1836
rect 18849 1806 18851 1834
rect 18851 1806 18879 1834
rect 18879 1806 18881 1834
rect 18849 1804 18881 1806
rect 18849 1674 18881 1676
rect 18849 1646 18851 1674
rect 18851 1646 18879 1674
rect 18879 1646 18881 1674
rect 18849 1644 18881 1646
rect 18849 1514 18881 1516
rect 18849 1486 18851 1514
rect 18851 1486 18879 1514
rect 18879 1486 18881 1514
rect 18849 1484 18881 1486
rect 18849 1354 18881 1356
rect 18849 1326 18851 1354
rect 18851 1326 18879 1354
rect 18879 1326 18881 1354
rect 18849 1324 18881 1326
rect 18849 1194 18881 1196
rect 18849 1166 18851 1194
rect 18851 1166 18879 1194
rect 18879 1166 18881 1194
rect 18849 1164 18881 1166
rect 18849 1034 18881 1036
rect 18849 1006 18851 1034
rect 18851 1006 18879 1034
rect 18879 1006 18881 1034
rect 18849 1004 18881 1006
rect 18849 874 18881 876
rect 18849 846 18851 874
rect 18851 846 18879 874
rect 18879 846 18881 874
rect 18849 844 18881 846
rect 18849 714 18881 716
rect 18849 686 18851 714
rect 18851 686 18879 714
rect 18879 686 18881 714
rect 18849 684 18881 686
rect 18849 554 18881 556
rect 18849 526 18851 554
rect 18851 526 18879 554
rect 18879 526 18881 554
rect 18849 524 18881 526
rect 18849 394 18881 396
rect 18849 366 18851 394
rect 18851 366 18879 394
rect 18879 366 18881 394
rect 18849 364 18881 366
rect 18849 234 18881 236
rect 18849 206 18851 234
rect 18851 206 18879 234
rect 18879 206 18881 234
rect 18849 204 18881 206
rect 18849 74 18881 76
rect 18849 46 18851 74
rect 18851 46 18879 74
rect 18879 46 18881 74
rect 18849 44 18881 46
rect 18849 -86 18881 -84
rect 18849 -114 18851 -86
rect 18851 -114 18879 -86
rect 18879 -114 18881 -86
rect 18849 -116 18881 -114
rect 15116 -246 15148 -244
rect 15116 -274 15118 -246
rect 15118 -274 15146 -246
rect 15146 -274 15148 -246
rect 15116 -276 15148 -274
rect 18849 -246 18881 -244
rect 18849 -274 18851 -246
rect 18851 -274 18879 -246
rect 18879 -274 18881 -246
rect 18849 -276 18881 -274
rect 15304 -349 15336 -347
rect 15304 -377 15306 -349
rect 15306 -377 15334 -349
rect 15334 -377 15336 -349
rect 15304 -379 15336 -377
rect 15464 -349 15496 -347
rect 15464 -377 15466 -349
rect 15466 -377 15494 -349
rect 15494 -377 15496 -349
rect 15464 -379 15496 -377
rect 15624 -349 15656 -347
rect 15624 -377 15626 -349
rect 15626 -377 15654 -349
rect 15654 -377 15656 -349
rect 15624 -379 15656 -377
rect 15784 -349 15816 -347
rect 15784 -377 15786 -349
rect 15786 -377 15814 -349
rect 15814 -377 15816 -349
rect 15784 -379 15816 -377
rect 15944 -349 15976 -347
rect 15944 -377 15946 -349
rect 15946 -377 15974 -349
rect 15974 -377 15976 -349
rect 15944 -379 15976 -377
rect 16104 -349 16136 -347
rect 16104 -377 16106 -349
rect 16106 -377 16134 -349
rect 16134 -377 16136 -349
rect 16104 -379 16136 -377
rect 16264 -349 16296 -347
rect 16264 -377 16266 -349
rect 16266 -377 16294 -349
rect 16294 -377 16296 -349
rect 16264 -379 16296 -377
rect 16424 -349 16456 -347
rect 16424 -377 16426 -349
rect 16426 -377 16454 -349
rect 16454 -377 16456 -349
rect 16424 -379 16456 -377
rect 16584 -349 16616 -347
rect 16584 -377 16586 -349
rect 16586 -377 16614 -349
rect 16614 -377 16616 -349
rect 16584 -379 16616 -377
rect 16744 -349 16776 -347
rect 16744 -377 16746 -349
rect 16746 -377 16774 -349
rect 16774 -377 16776 -349
rect 16744 -379 16776 -377
rect 16904 -349 16936 -347
rect 16904 -377 16906 -349
rect 16906 -377 16934 -349
rect 16934 -377 16936 -349
rect 16904 -379 16936 -377
rect 17064 -349 17096 -347
rect 17064 -377 17066 -349
rect 17066 -377 17094 -349
rect 17094 -377 17096 -349
rect 17064 -379 17096 -377
rect 17224 -349 17256 -347
rect 17224 -377 17226 -349
rect 17226 -377 17254 -349
rect 17254 -377 17256 -349
rect 17224 -379 17256 -377
rect 17384 -349 17416 -347
rect 17384 -377 17386 -349
rect 17386 -377 17414 -349
rect 17414 -377 17416 -349
rect 17384 -379 17416 -377
rect 17544 -349 17576 -347
rect 17544 -377 17546 -349
rect 17546 -377 17574 -349
rect 17574 -377 17576 -349
rect 17544 -379 17576 -377
rect 17704 -349 17736 -347
rect 17704 -377 17706 -349
rect 17706 -377 17734 -349
rect 17734 -377 17736 -349
rect 17704 -379 17736 -377
rect 17864 -349 17896 -347
rect 17864 -377 17866 -349
rect 17866 -377 17894 -349
rect 17894 -377 17896 -349
rect 17864 -379 17896 -377
rect 18024 -349 18056 -347
rect 18024 -377 18026 -349
rect 18026 -377 18054 -349
rect 18054 -377 18056 -349
rect 18024 -379 18056 -377
rect 18184 -349 18216 -347
rect 18184 -377 18186 -349
rect 18186 -377 18214 -349
rect 18214 -377 18216 -349
rect 18184 -379 18216 -377
rect 18344 -349 18376 -347
rect 18344 -377 18346 -349
rect 18346 -377 18374 -349
rect 18374 -377 18376 -349
rect 18344 -379 18376 -377
rect 18504 -349 18536 -347
rect 18504 -377 18506 -349
rect 18506 -377 18534 -349
rect 18534 -377 18536 -349
rect 18504 -379 18536 -377
rect 18664 -349 18696 -347
rect 18664 -377 18666 -349
rect 18666 -377 18694 -349
rect 18694 -377 18696 -349
rect 18664 -379 18696 -377
rect 21116 6874 21148 6876
rect 21116 6846 21118 6874
rect 21118 6846 21146 6874
rect 21146 6846 21148 6874
rect 21116 6844 21148 6846
rect 21116 6714 21148 6716
rect 21116 6686 21118 6714
rect 21118 6686 21146 6714
rect 21146 6686 21148 6714
rect 21116 6684 21148 6686
rect 21116 6554 21148 6556
rect 21116 6526 21118 6554
rect 21118 6526 21146 6554
rect 21146 6526 21148 6554
rect 21116 6524 21148 6526
rect 21116 6394 21148 6396
rect 21116 6366 21118 6394
rect 21118 6366 21146 6394
rect 21146 6366 21148 6394
rect 21116 6364 21148 6366
rect 21116 6234 21148 6236
rect 21116 6206 21118 6234
rect 21118 6206 21146 6234
rect 21146 6206 21148 6234
rect 21116 6204 21148 6206
rect 21116 6074 21148 6076
rect 21116 6046 21118 6074
rect 21118 6046 21146 6074
rect 21146 6046 21148 6074
rect 21116 6044 21148 6046
rect 21116 5914 21148 5916
rect 21116 5886 21118 5914
rect 21118 5886 21146 5914
rect 21146 5886 21148 5914
rect 21116 5884 21148 5886
rect 24849 9114 24881 9116
rect 24849 9086 24851 9114
rect 24851 9086 24879 9114
rect 24879 9086 24881 9114
rect 24849 9084 24881 9086
rect 24849 8954 24881 8956
rect 24849 8926 24851 8954
rect 24851 8926 24879 8954
rect 24879 8926 24881 8954
rect 24849 8924 24881 8926
rect 24849 8794 24881 8796
rect 24849 8766 24851 8794
rect 24851 8766 24879 8794
rect 24879 8766 24881 8794
rect 24849 8764 24881 8766
rect 24849 8634 24881 8636
rect 24849 8606 24851 8634
rect 24851 8606 24879 8634
rect 24879 8606 24881 8634
rect 24849 8604 24881 8606
rect 24849 8474 24881 8476
rect 24849 8446 24851 8474
rect 24851 8446 24879 8474
rect 24879 8446 24881 8474
rect 24849 8444 24881 8446
rect 24849 8314 24881 8316
rect 24849 8286 24851 8314
rect 24851 8286 24879 8314
rect 24879 8286 24881 8314
rect 24849 8284 24881 8286
rect 24849 8154 24881 8156
rect 24849 8126 24851 8154
rect 24851 8126 24879 8154
rect 24879 8126 24881 8154
rect 24849 8124 24881 8126
rect 24849 7994 24881 7996
rect 24849 7966 24851 7994
rect 24851 7966 24879 7994
rect 24879 7966 24881 7994
rect 24849 7964 24881 7966
rect 24849 7834 24881 7836
rect 24849 7806 24851 7834
rect 24851 7806 24879 7834
rect 24879 7806 24881 7834
rect 24849 7804 24881 7806
rect 24849 7674 24881 7676
rect 24849 7646 24851 7674
rect 24851 7646 24879 7674
rect 24879 7646 24881 7674
rect 24849 7644 24881 7646
rect 24849 7514 24881 7516
rect 24849 7486 24851 7514
rect 24851 7486 24879 7514
rect 24879 7486 24881 7514
rect 24849 7484 24881 7486
rect 24849 7354 24881 7356
rect 24849 7326 24851 7354
rect 24851 7326 24879 7354
rect 24879 7326 24881 7354
rect 24849 7324 24881 7326
rect 24849 7194 24881 7196
rect 24849 7166 24851 7194
rect 24851 7166 24879 7194
rect 24879 7166 24881 7194
rect 24849 7164 24881 7166
rect 24849 7034 24881 7036
rect 24849 7006 24851 7034
rect 24851 7006 24879 7034
rect 24879 7006 24881 7034
rect 24849 7004 24881 7006
rect 24849 6874 24881 6876
rect 24849 6846 24851 6874
rect 24851 6846 24879 6874
rect 24879 6846 24881 6874
rect 24849 6844 24881 6846
rect 24849 6714 24881 6716
rect 24849 6686 24851 6714
rect 24851 6686 24879 6714
rect 24879 6686 24881 6714
rect 24849 6684 24881 6686
rect 24849 6554 24881 6556
rect 24849 6526 24851 6554
rect 24851 6526 24879 6554
rect 24879 6526 24881 6554
rect 24849 6524 24881 6526
rect 24849 6394 24881 6396
rect 24849 6366 24851 6394
rect 24851 6366 24879 6394
rect 24879 6366 24881 6394
rect 24849 6364 24881 6366
rect 24849 6234 24881 6236
rect 24849 6206 24851 6234
rect 24851 6206 24879 6234
rect 24879 6206 24881 6234
rect 24849 6204 24881 6206
rect 24849 6074 24881 6076
rect 24849 6046 24851 6074
rect 24851 6046 24879 6074
rect 24879 6046 24881 6074
rect 24849 6044 24881 6046
rect 24849 5914 24881 5916
rect 24849 5886 24851 5914
rect 24851 5886 24879 5914
rect 24879 5886 24881 5914
rect 24849 5884 24881 5886
rect 21116 5754 21148 5756
rect 21116 5726 21118 5754
rect 21118 5726 21146 5754
rect 21146 5726 21148 5754
rect 21116 5724 21148 5726
rect 24849 5754 24881 5756
rect 24849 5726 24851 5754
rect 24851 5726 24879 5754
rect 24879 5726 24881 5754
rect 24849 5724 24881 5726
rect 21304 5651 21336 5653
rect 21304 5623 21306 5651
rect 21306 5623 21334 5651
rect 21334 5623 21336 5651
rect 21304 5621 21336 5623
rect 21464 5651 21496 5653
rect 21464 5623 21466 5651
rect 21466 5623 21494 5651
rect 21494 5623 21496 5651
rect 21464 5621 21496 5623
rect 21624 5651 21656 5653
rect 21624 5623 21626 5651
rect 21626 5623 21654 5651
rect 21654 5623 21656 5651
rect 21624 5621 21656 5623
rect 21784 5651 21816 5653
rect 21784 5623 21786 5651
rect 21786 5623 21814 5651
rect 21814 5623 21816 5651
rect 21784 5621 21816 5623
rect 21944 5651 21976 5653
rect 21944 5623 21946 5651
rect 21946 5623 21974 5651
rect 21974 5623 21976 5651
rect 21944 5621 21976 5623
rect 22104 5651 22136 5653
rect 22104 5623 22106 5651
rect 22106 5623 22134 5651
rect 22134 5623 22136 5651
rect 22104 5621 22136 5623
rect 22264 5651 22296 5653
rect 22264 5623 22266 5651
rect 22266 5623 22294 5651
rect 22294 5623 22296 5651
rect 22264 5621 22296 5623
rect 22424 5651 22456 5653
rect 22424 5623 22426 5651
rect 22426 5623 22454 5651
rect 22454 5623 22456 5651
rect 22424 5621 22456 5623
rect 22584 5651 22616 5653
rect 22584 5623 22586 5651
rect 22586 5623 22614 5651
rect 22614 5623 22616 5651
rect 22584 5621 22616 5623
rect 22744 5651 22776 5653
rect 22744 5623 22746 5651
rect 22746 5623 22774 5651
rect 22774 5623 22776 5651
rect 22744 5621 22776 5623
rect 22904 5651 22936 5653
rect 22904 5623 22906 5651
rect 22906 5623 22934 5651
rect 22934 5623 22936 5651
rect 22904 5621 22936 5623
rect 23064 5651 23096 5653
rect 23064 5623 23066 5651
rect 23066 5623 23094 5651
rect 23094 5623 23096 5651
rect 23064 5621 23096 5623
rect 23224 5651 23256 5653
rect 23224 5623 23226 5651
rect 23226 5623 23254 5651
rect 23254 5623 23256 5651
rect 23224 5621 23256 5623
rect 23384 5651 23416 5653
rect 23384 5623 23386 5651
rect 23386 5623 23414 5651
rect 23414 5623 23416 5651
rect 23384 5621 23416 5623
rect 23544 5651 23576 5653
rect 23544 5623 23546 5651
rect 23546 5623 23574 5651
rect 23574 5623 23576 5651
rect 23544 5621 23576 5623
rect 23704 5651 23736 5653
rect 23704 5623 23706 5651
rect 23706 5623 23734 5651
rect 23734 5623 23736 5651
rect 23704 5621 23736 5623
rect 23864 5651 23896 5653
rect 23864 5623 23866 5651
rect 23866 5623 23894 5651
rect 23894 5623 23896 5651
rect 23864 5621 23896 5623
rect 24024 5651 24056 5653
rect 24024 5623 24026 5651
rect 24026 5623 24054 5651
rect 24054 5623 24056 5651
rect 24024 5621 24056 5623
rect 24184 5651 24216 5653
rect 24184 5623 24186 5651
rect 24186 5623 24214 5651
rect 24214 5623 24216 5651
rect 24184 5621 24216 5623
rect 24344 5651 24376 5653
rect 24344 5623 24346 5651
rect 24346 5623 24374 5651
rect 24374 5623 24376 5651
rect 24344 5621 24376 5623
rect 24504 5651 24536 5653
rect 24504 5623 24506 5651
rect 24506 5623 24534 5651
rect 24534 5623 24536 5651
rect 24504 5621 24536 5623
rect 24664 5651 24696 5653
rect 24664 5623 24666 5651
rect 24666 5623 24694 5651
rect 24694 5623 24696 5651
rect 24664 5621 24696 5623
rect 21304 3379 21336 3381
rect 21304 3351 21306 3379
rect 21306 3351 21334 3379
rect 21334 3351 21336 3379
rect 21304 3349 21336 3351
rect 21464 3379 21496 3381
rect 21464 3351 21466 3379
rect 21466 3351 21494 3379
rect 21494 3351 21496 3379
rect 21464 3349 21496 3351
rect 21624 3379 21656 3381
rect 21624 3351 21626 3379
rect 21626 3351 21654 3379
rect 21654 3351 21656 3379
rect 21624 3349 21656 3351
rect 21784 3379 21816 3381
rect 21784 3351 21786 3379
rect 21786 3351 21814 3379
rect 21814 3351 21816 3379
rect 21784 3349 21816 3351
rect 21944 3379 21976 3381
rect 21944 3351 21946 3379
rect 21946 3351 21974 3379
rect 21974 3351 21976 3379
rect 21944 3349 21976 3351
rect 22104 3379 22136 3381
rect 22104 3351 22106 3379
rect 22106 3351 22134 3379
rect 22134 3351 22136 3379
rect 22104 3349 22136 3351
rect 22264 3379 22296 3381
rect 22264 3351 22266 3379
rect 22266 3351 22294 3379
rect 22294 3351 22296 3379
rect 22264 3349 22296 3351
rect 22424 3379 22456 3381
rect 22424 3351 22426 3379
rect 22426 3351 22454 3379
rect 22454 3351 22456 3379
rect 22424 3349 22456 3351
rect 22584 3379 22616 3381
rect 22584 3351 22586 3379
rect 22586 3351 22614 3379
rect 22614 3351 22616 3379
rect 22584 3349 22616 3351
rect 22744 3379 22776 3381
rect 22744 3351 22746 3379
rect 22746 3351 22774 3379
rect 22774 3351 22776 3379
rect 22744 3349 22776 3351
rect 22904 3379 22936 3381
rect 22904 3351 22906 3379
rect 22906 3351 22934 3379
rect 22934 3351 22936 3379
rect 22904 3349 22936 3351
rect 23064 3379 23096 3381
rect 23064 3351 23066 3379
rect 23066 3351 23094 3379
rect 23094 3351 23096 3379
rect 23064 3349 23096 3351
rect 23224 3379 23256 3381
rect 23224 3351 23226 3379
rect 23226 3351 23254 3379
rect 23254 3351 23256 3379
rect 23224 3349 23256 3351
rect 23384 3379 23416 3381
rect 23384 3351 23386 3379
rect 23386 3351 23414 3379
rect 23414 3351 23416 3379
rect 23384 3349 23416 3351
rect 23544 3379 23576 3381
rect 23544 3351 23546 3379
rect 23546 3351 23574 3379
rect 23574 3351 23576 3379
rect 23544 3349 23576 3351
rect 23704 3379 23736 3381
rect 23704 3351 23706 3379
rect 23706 3351 23734 3379
rect 23734 3351 23736 3379
rect 23704 3349 23736 3351
rect 23864 3379 23896 3381
rect 23864 3351 23866 3379
rect 23866 3351 23894 3379
rect 23894 3351 23896 3379
rect 23864 3349 23896 3351
rect 24024 3379 24056 3381
rect 24024 3351 24026 3379
rect 24026 3351 24054 3379
rect 24054 3351 24056 3379
rect 24024 3349 24056 3351
rect 24184 3379 24216 3381
rect 24184 3351 24186 3379
rect 24186 3351 24214 3379
rect 24214 3351 24216 3379
rect 24184 3349 24216 3351
rect 24344 3379 24376 3381
rect 24344 3351 24346 3379
rect 24346 3351 24374 3379
rect 24374 3351 24376 3379
rect 24344 3349 24376 3351
rect 24504 3379 24536 3381
rect 24504 3351 24506 3379
rect 24506 3351 24534 3379
rect 24534 3351 24536 3379
rect 24504 3349 24536 3351
rect 24664 3379 24696 3381
rect 24664 3351 24666 3379
rect 24666 3351 24694 3379
rect 24694 3351 24696 3379
rect 24664 3349 24696 3351
rect 21116 3274 21148 3276
rect 21116 3246 21118 3274
rect 21118 3246 21146 3274
rect 21146 3246 21148 3274
rect 21116 3244 21148 3246
rect 24849 3274 24881 3276
rect 24849 3246 24851 3274
rect 24851 3246 24879 3274
rect 24879 3246 24881 3274
rect 24849 3244 24881 3246
rect 21116 3114 21148 3116
rect 21116 3086 21118 3114
rect 21118 3086 21146 3114
rect 21146 3086 21148 3114
rect 21116 3084 21148 3086
rect 21116 2954 21148 2956
rect 21116 2926 21118 2954
rect 21118 2926 21146 2954
rect 21146 2926 21148 2954
rect 21116 2924 21148 2926
rect 21116 2794 21148 2796
rect 21116 2766 21118 2794
rect 21118 2766 21146 2794
rect 21146 2766 21148 2794
rect 21116 2764 21148 2766
rect 21116 2634 21148 2636
rect 21116 2606 21118 2634
rect 21118 2606 21146 2634
rect 21146 2606 21148 2634
rect 21116 2604 21148 2606
rect 21116 2474 21148 2476
rect 21116 2446 21118 2474
rect 21118 2446 21146 2474
rect 21146 2446 21148 2474
rect 21116 2444 21148 2446
rect 21116 2314 21148 2316
rect 21116 2286 21118 2314
rect 21118 2286 21146 2314
rect 21146 2286 21148 2314
rect 21116 2284 21148 2286
rect 21116 2154 21148 2156
rect 21116 2126 21118 2154
rect 21118 2126 21146 2154
rect 21146 2126 21148 2154
rect 21116 2124 21148 2126
rect 21116 1994 21148 1996
rect 21116 1966 21118 1994
rect 21118 1966 21146 1994
rect 21146 1966 21148 1994
rect 21116 1964 21148 1966
rect 21116 1834 21148 1836
rect 21116 1806 21118 1834
rect 21118 1806 21146 1834
rect 21146 1806 21148 1834
rect 21116 1804 21148 1806
rect 21116 1674 21148 1676
rect 21116 1646 21118 1674
rect 21118 1646 21146 1674
rect 21146 1646 21148 1674
rect 21116 1644 21148 1646
rect 21116 1514 21148 1516
rect 21116 1486 21118 1514
rect 21118 1486 21146 1514
rect 21146 1486 21148 1514
rect 21116 1484 21148 1486
rect 21116 1354 21148 1356
rect 21116 1326 21118 1354
rect 21118 1326 21146 1354
rect 21146 1326 21148 1354
rect 21116 1324 21148 1326
rect 21116 1194 21148 1196
rect 21116 1166 21118 1194
rect 21118 1166 21146 1194
rect 21146 1166 21148 1194
rect 21116 1164 21148 1166
rect 21116 1034 21148 1036
rect 21116 1006 21118 1034
rect 21118 1006 21146 1034
rect 21146 1006 21148 1034
rect 21116 1004 21148 1006
rect 21116 874 21148 876
rect 21116 846 21118 874
rect 21118 846 21146 874
rect 21146 846 21148 874
rect 21116 844 21148 846
rect 21116 714 21148 716
rect 21116 686 21118 714
rect 21118 686 21146 714
rect 21146 686 21148 714
rect 21116 684 21148 686
rect 21116 554 21148 556
rect 21116 526 21118 554
rect 21118 526 21146 554
rect 21146 526 21148 554
rect 21116 524 21148 526
rect 21116 394 21148 396
rect 21116 366 21118 394
rect 21118 366 21146 394
rect 21146 366 21148 394
rect 21116 364 21148 366
rect 21116 234 21148 236
rect 21116 206 21118 234
rect 21118 206 21146 234
rect 21146 206 21148 234
rect 21116 204 21148 206
rect 21116 74 21148 76
rect 21116 46 21118 74
rect 21118 46 21146 74
rect 21146 46 21148 74
rect 21116 44 21148 46
rect 21116 -86 21148 -84
rect 21116 -114 21118 -86
rect 21118 -114 21146 -86
rect 21146 -114 21148 -86
rect 21116 -116 21148 -114
rect 24849 3114 24881 3116
rect 24849 3086 24851 3114
rect 24851 3086 24879 3114
rect 24879 3086 24881 3114
rect 24849 3084 24881 3086
rect 24849 2954 24881 2956
rect 24849 2926 24851 2954
rect 24851 2926 24879 2954
rect 24879 2926 24881 2954
rect 24849 2924 24881 2926
rect 24849 2794 24881 2796
rect 24849 2766 24851 2794
rect 24851 2766 24879 2794
rect 24879 2766 24881 2794
rect 24849 2764 24881 2766
rect 24849 2634 24881 2636
rect 24849 2606 24851 2634
rect 24851 2606 24879 2634
rect 24879 2606 24881 2634
rect 24849 2604 24881 2606
rect 24849 2474 24881 2476
rect 24849 2446 24851 2474
rect 24851 2446 24879 2474
rect 24879 2446 24881 2474
rect 24849 2444 24881 2446
rect 24849 2314 24881 2316
rect 24849 2286 24851 2314
rect 24851 2286 24879 2314
rect 24879 2286 24881 2314
rect 24849 2284 24881 2286
rect 24849 2154 24881 2156
rect 24849 2126 24851 2154
rect 24851 2126 24879 2154
rect 24879 2126 24881 2154
rect 24849 2124 24881 2126
rect 24849 1994 24881 1996
rect 24849 1966 24851 1994
rect 24851 1966 24879 1994
rect 24879 1966 24881 1994
rect 24849 1964 24881 1966
rect 24849 1834 24881 1836
rect 24849 1806 24851 1834
rect 24851 1806 24879 1834
rect 24879 1806 24881 1834
rect 24849 1804 24881 1806
rect 24849 1674 24881 1676
rect 24849 1646 24851 1674
rect 24851 1646 24879 1674
rect 24879 1646 24881 1674
rect 24849 1644 24881 1646
rect 24849 1514 24881 1516
rect 24849 1486 24851 1514
rect 24851 1486 24879 1514
rect 24879 1486 24881 1514
rect 24849 1484 24881 1486
rect 24849 1354 24881 1356
rect 24849 1326 24851 1354
rect 24851 1326 24879 1354
rect 24879 1326 24881 1354
rect 24849 1324 24881 1326
rect 24849 1194 24881 1196
rect 24849 1166 24851 1194
rect 24851 1166 24879 1194
rect 24879 1166 24881 1194
rect 24849 1164 24881 1166
rect 24849 1034 24881 1036
rect 24849 1006 24851 1034
rect 24851 1006 24879 1034
rect 24879 1006 24881 1034
rect 24849 1004 24881 1006
rect 24849 874 24881 876
rect 24849 846 24851 874
rect 24851 846 24879 874
rect 24879 846 24881 874
rect 24849 844 24881 846
rect 24849 714 24881 716
rect 24849 686 24851 714
rect 24851 686 24879 714
rect 24879 686 24881 714
rect 24849 684 24881 686
rect 24849 554 24881 556
rect 24849 526 24851 554
rect 24851 526 24879 554
rect 24879 526 24881 554
rect 24849 524 24881 526
rect 24849 394 24881 396
rect 24849 366 24851 394
rect 24851 366 24879 394
rect 24879 366 24881 394
rect 24849 364 24881 366
rect 24849 234 24881 236
rect 24849 206 24851 234
rect 24851 206 24879 234
rect 24879 206 24881 234
rect 24849 204 24881 206
rect 24849 74 24881 76
rect 24849 46 24851 74
rect 24851 46 24879 74
rect 24879 46 24881 74
rect 24849 44 24881 46
rect 24849 -86 24881 -84
rect 24849 -114 24851 -86
rect 24851 -114 24879 -86
rect 24879 -114 24881 -86
rect 24849 -116 24881 -114
rect 21116 -246 21148 -244
rect 21116 -274 21118 -246
rect 21118 -274 21146 -246
rect 21146 -274 21148 -246
rect 21116 -276 21148 -274
rect 24849 -246 24881 -244
rect 24849 -274 24851 -246
rect 24851 -274 24879 -246
rect 24879 -274 24881 -246
rect 24849 -276 24881 -274
rect 21304 -349 21336 -347
rect 21304 -377 21306 -349
rect 21306 -377 21334 -349
rect 21334 -377 21336 -349
rect 21304 -379 21336 -377
rect 21464 -349 21496 -347
rect 21464 -377 21466 -349
rect 21466 -377 21494 -349
rect 21494 -377 21496 -349
rect 21464 -379 21496 -377
rect 21624 -349 21656 -347
rect 21624 -377 21626 -349
rect 21626 -377 21654 -349
rect 21654 -377 21656 -349
rect 21624 -379 21656 -377
rect 21784 -349 21816 -347
rect 21784 -377 21786 -349
rect 21786 -377 21814 -349
rect 21814 -377 21816 -349
rect 21784 -379 21816 -377
rect 21944 -349 21976 -347
rect 21944 -377 21946 -349
rect 21946 -377 21974 -349
rect 21974 -377 21976 -349
rect 21944 -379 21976 -377
rect 22104 -349 22136 -347
rect 22104 -377 22106 -349
rect 22106 -377 22134 -349
rect 22134 -377 22136 -349
rect 22104 -379 22136 -377
rect 22264 -349 22296 -347
rect 22264 -377 22266 -349
rect 22266 -377 22294 -349
rect 22294 -377 22296 -349
rect 22264 -379 22296 -377
rect 22424 -349 22456 -347
rect 22424 -377 22426 -349
rect 22426 -377 22454 -349
rect 22454 -377 22456 -349
rect 22424 -379 22456 -377
rect 22584 -349 22616 -347
rect 22584 -377 22586 -349
rect 22586 -377 22614 -349
rect 22614 -377 22616 -349
rect 22584 -379 22616 -377
rect 22744 -349 22776 -347
rect 22744 -377 22746 -349
rect 22746 -377 22774 -349
rect 22774 -377 22776 -349
rect 22744 -379 22776 -377
rect 22904 -349 22936 -347
rect 22904 -377 22906 -349
rect 22906 -377 22934 -349
rect 22934 -377 22936 -349
rect 22904 -379 22936 -377
rect 23064 -349 23096 -347
rect 23064 -377 23066 -349
rect 23066 -377 23094 -349
rect 23094 -377 23096 -349
rect 23064 -379 23096 -377
rect 23224 -349 23256 -347
rect 23224 -377 23226 -349
rect 23226 -377 23254 -349
rect 23254 -377 23256 -349
rect 23224 -379 23256 -377
rect 23384 -349 23416 -347
rect 23384 -377 23386 -349
rect 23386 -377 23414 -349
rect 23414 -377 23416 -349
rect 23384 -379 23416 -377
rect 23544 -349 23576 -347
rect 23544 -377 23546 -349
rect 23546 -377 23574 -349
rect 23574 -377 23576 -349
rect 23544 -379 23576 -377
rect 23704 -349 23736 -347
rect 23704 -377 23706 -349
rect 23706 -377 23734 -349
rect 23734 -377 23736 -349
rect 23704 -379 23736 -377
rect 23864 -349 23896 -347
rect 23864 -377 23866 -349
rect 23866 -377 23894 -349
rect 23894 -377 23896 -349
rect 23864 -379 23896 -377
rect 24024 -349 24056 -347
rect 24024 -377 24026 -349
rect 24026 -377 24054 -349
rect 24054 -377 24056 -349
rect 24024 -379 24056 -377
rect 24184 -349 24216 -347
rect 24184 -377 24186 -349
rect 24186 -377 24214 -349
rect 24214 -377 24216 -349
rect 24184 -379 24216 -377
rect 24344 -349 24376 -347
rect 24344 -377 24346 -349
rect 24346 -377 24374 -349
rect 24374 -377 24376 -349
rect 24344 -379 24376 -377
rect 24504 -349 24536 -347
rect 24504 -377 24506 -349
rect 24506 -377 24534 -349
rect 24534 -377 24536 -349
rect 24504 -379 24536 -377
rect 24664 -349 24696 -347
rect 24664 -377 24666 -349
rect 24666 -377 24694 -349
rect 24694 -377 24696 -349
rect 24664 -379 24696 -377
rect 3304 -5623 3336 -5621
rect 3304 -5651 3306 -5623
rect 3306 -5651 3334 -5623
rect 3334 -5651 3336 -5623
rect 3304 -5653 3336 -5651
rect 3464 -5623 3496 -5621
rect 3464 -5651 3466 -5623
rect 3466 -5651 3494 -5623
rect 3494 -5651 3496 -5623
rect 3464 -5653 3496 -5651
rect 3624 -5623 3656 -5621
rect 3624 -5651 3626 -5623
rect 3626 -5651 3654 -5623
rect 3654 -5651 3656 -5623
rect 3624 -5653 3656 -5651
rect 3784 -5623 3816 -5621
rect 3784 -5651 3786 -5623
rect 3786 -5651 3814 -5623
rect 3814 -5651 3816 -5623
rect 3784 -5653 3816 -5651
rect 3944 -5623 3976 -5621
rect 3944 -5651 3946 -5623
rect 3946 -5651 3974 -5623
rect 3974 -5651 3976 -5623
rect 3944 -5653 3976 -5651
rect 4104 -5623 4136 -5621
rect 4104 -5651 4106 -5623
rect 4106 -5651 4134 -5623
rect 4134 -5651 4136 -5623
rect 4104 -5653 4136 -5651
rect 4264 -5623 4296 -5621
rect 4264 -5651 4266 -5623
rect 4266 -5651 4294 -5623
rect 4294 -5651 4296 -5623
rect 4264 -5653 4296 -5651
rect 4424 -5623 4456 -5621
rect 4424 -5651 4426 -5623
rect 4426 -5651 4454 -5623
rect 4454 -5651 4456 -5623
rect 4424 -5653 4456 -5651
rect 4584 -5623 4616 -5621
rect 4584 -5651 4586 -5623
rect 4586 -5651 4614 -5623
rect 4614 -5651 4616 -5623
rect 4584 -5653 4616 -5651
rect 4744 -5623 4776 -5621
rect 4744 -5651 4746 -5623
rect 4746 -5651 4774 -5623
rect 4774 -5651 4776 -5623
rect 4744 -5653 4776 -5651
rect 4904 -5623 4936 -5621
rect 4904 -5651 4906 -5623
rect 4906 -5651 4934 -5623
rect 4934 -5651 4936 -5623
rect 4904 -5653 4936 -5651
rect 5064 -5623 5096 -5621
rect 5064 -5651 5066 -5623
rect 5066 -5651 5094 -5623
rect 5094 -5651 5096 -5623
rect 5064 -5653 5096 -5651
rect 5224 -5623 5256 -5621
rect 5224 -5651 5226 -5623
rect 5226 -5651 5254 -5623
rect 5254 -5651 5256 -5623
rect 5224 -5653 5256 -5651
rect 5384 -5623 5416 -5621
rect 5384 -5651 5386 -5623
rect 5386 -5651 5414 -5623
rect 5414 -5651 5416 -5623
rect 5384 -5653 5416 -5651
rect 5544 -5623 5576 -5621
rect 5544 -5651 5546 -5623
rect 5546 -5651 5574 -5623
rect 5574 -5651 5576 -5623
rect 5544 -5653 5576 -5651
rect 5704 -5623 5736 -5621
rect 5704 -5651 5706 -5623
rect 5706 -5651 5734 -5623
rect 5734 -5651 5736 -5623
rect 5704 -5653 5736 -5651
rect 5864 -5623 5896 -5621
rect 5864 -5651 5866 -5623
rect 5866 -5651 5894 -5623
rect 5894 -5651 5896 -5623
rect 5864 -5653 5896 -5651
rect 6024 -5623 6056 -5621
rect 6024 -5651 6026 -5623
rect 6026 -5651 6054 -5623
rect 6054 -5651 6056 -5623
rect 6024 -5653 6056 -5651
rect 6184 -5623 6216 -5621
rect 6184 -5651 6186 -5623
rect 6186 -5651 6214 -5623
rect 6214 -5651 6216 -5623
rect 6184 -5653 6216 -5651
rect 6344 -5623 6376 -5621
rect 6344 -5651 6346 -5623
rect 6346 -5651 6374 -5623
rect 6374 -5651 6376 -5623
rect 6344 -5653 6376 -5651
rect 6504 -5623 6536 -5621
rect 6504 -5651 6506 -5623
rect 6506 -5651 6534 -5623
rect 6534 -5651 6536 -5623
rect 6504 -5653 6536 -5651
rect 6664 -5623 6696 -5621
rect 6664 -5651 6666 -5623
rect 6666 -5651 6694 -5623
rect 6694 -5651 6696 -5623
rect 6664 -5653 6696 -5651
rect 3119 -5726 3151 -5724
rect 3119 -5754 3121 -5726
rect 3121 -5754 3149 -5726
rect 3149 -5754 3151 -5726
rect 3119 -5756 3151 -5754
rect 6852 -5726 6884 -5724
rect 6852 -5754 6854 -5726
rect 6854 -5754 6882 -5726
rect 6882 -5754 6884 -5726
rect 6852 -5756 6884 -5754
rect 3119 -5886 3151 -5884
rect 3119 -5914 3121 -5886
rect 3121 -5914 3149 -5886
rect 3149 -5914 3151 -5886
rect 3119 -5916 3151 -5914
rect 3119 -6046 3151 -6044
rect 3119 -6074 3121 -6046
rect 3121 -6074 3149 -6046
rect 3149 -6074 3151 -6046
rect 3119 -6076 3151 -6074
rect 3119 -6206 3151 -6204
rect 3119 -6234 3121 -6206
rect 3121 -6234 3149 -6206
rect 3149 -6234 3151 -6206
rect 3119 -6236 3151 -6234
rect 3119 -6366 3151 -6364
rect 3119 -6394 3121 -6366
rect 3121 -6394 3149 -6366
rect 3149 -6394 3151 -6366
rect 3119 -6396 3151 -6394
rect 3119 -6526 3151 -6524
rect 3119 -6554 3121 -6526
rect 3121 -6554 3149 -6526
rect 3149 -6554 3151 -6526
rect 3119 -6556 3151 -6554
rect 3119 -6686 3151 -6684
rect 3119 -6714 3121 -6686
rect 3121 -6714 3149 -6686
rect 3149 -6714 3151 -6686
rect 3119 -6716 3151 -6714
rect 3119 -6846 3151 -6844
rect 3119 -6874 3121 -6846
rect 3121 -6874 3149 -6846
rect 3149 -6874 3151 -6846
rect 3119 -6876 3151 -6874
rect 3119 -7006 3151 -7004
rect 3119 -7034 3121 -7006
rect 3121 -7034 3149 -7006
rect 3149 -7034 3151 -7006
rect 3119 -7036 3151 -7034
rect 3119 -7166 3151 -7164
rect 3119 -7194 3121 -7166
rect 3121 -7194 3149 -7166
rect 3149 -7194 3151 -7166
rect 3119 -7196 3151 -7194
rect 3119 -7326 3151 -7324
rect 3119 -7354 3121 -7326
rect 3121 -7354 3149 -7326
rect 3149 -7354 3151 -7326
rect 3119 -7356 3151 -7354
rect 3119 -7486 3151 -7484
rect 3119 -7514 3121 -7486
rect 3121 -7514 3149 -7486
rect 3149 -7514 3151 -7486
rect 3119 -7516 3151 -7514
rect 3119 -7646 3151 -7644
rect 3119 -7674 3121 -7646
rect 3121 -7674 3149 -7646
rect 3149 -7674 3151 -7646
rect 3119 -7676 3151 -7674
rect 3119 -7806 3151 -7804
rect 3119 -7834 3121 -7806
rect 3121 -7834 3149 -7806
rect 3149 -7834 3151 -7806
rect 3119 -7836 3151 -7834
rect 3119 -7966 3151 -7964
rect 3119 -7994 3121 -7966
rect 3121 -7994 3149 -7966
rect 3149 -7994 3151 -7966
rect 3119 -7996 3151 -7994
rect 3119 -8126 3151 -8124
rect 3119 -8154 3121 -8126
rect 3121 -8154 3149 -8126
rect 3149 -8154 3151 -8126
rect 3119 -8156 3151 -8154
rect 3119 -8286 3151 -8284
rect 3119 -8314 3121 -8286
rect 3121 -8314 3149 -8286
rect 3149 -8314 3151 -8286
rect 3119 -8316 3151 -8314
rect 3119 -8446 3151 -8444
rect 3119 -8474 3121 -8446
rect 3121 -8474 3149 -8446
rect 3149 -8474 3151 -8446
rect 3119 -8476 3151 -8474
rect 3119 -8606 3151 -8604
rect 3119 -8634 3121 -8606
rect 3121 -8634 3149 -8606
rect 3149 -8634 3151 -8606
rect 3119 -8636 3151 -8634
rect 3119 -8766 3151 -8764
rect 3119 -8794 3121 -8766
rect 3121 -8794 3149 -8766
rect 3149 -8794 3151 -8766
rect 3119 -8796 3151 -8794
rect 3119 -8926 3151 -8924
rect 3119 -8954 3121 -8926
rect 3121 -8954 3149 -8926
rect 3149 -8954 3151 -8926
rect 3119 -8956 3151 -8954
rect 3119 -9086 3151 -9084
rect 3119 -9114 3121 -9086
rect 3121 -9114 3149 -9086
rect 3149 -9114 3151 -9086
rect 3119 -9116 3151 -9114
rect 6852 -5886 6884 -5884
rect 6852 -5914 6854 -5886
rect 6854 -5914 6882 -5886
rect 6882 -5914 6884 -5886
rect 6852 -5916 6884 -5914
rect 6852 -6046 6884 -6044
rect 6852 -6074 6854 -6046
rect 6854 -6074 6882 -6046
rect 6882 -6074 6884 -6046
rect 6852 -6076 6884 -6074
rect 6852 -6206 6884 -6204
rect 6852 -6234 6854 -6206
rect 6854 -6234 6882 -6206
rect 6882 -6234 6884 -6206
rect 6852 -6236 6884 -6234
rect 6852 -6366 6884 -6364
rect 6852 -6394 6854 -6366
rect 6854 -6394 6882 -6366
rect 6882 -6394 6884 -6366
rect 6852 -6396 6884 -6394
rect 6852 -6526 6884 -6524
rect 6852 -6554 6854 -6526
rect 6854 -6554 6882 -6526
rect 6882 -6554 6884 -6526
rect 6852 -6556 6884 -6554
rect 6852 -6686 6884 -6684
rect 6852 -6714 6854 -6686
rect 6854 -6714 6882 -6686
rect 6882 -6714 6884 -6686
rect 6852 -6716 6884 -6714
rect 6852 -6846 6884 -6844
rect 6852 -6874 6854 -6846
rect 6854 -6874 6882 -6846
rect 6882 -6874 6884 -6846
rect 6852 -6876 6884 -6874
rect 6852 -7006 6884 -7004
rect 6852 -7034 6854 -7006
rect 6854 -7034 6882 -7006
rect 6882 -7034 6884 -7006
rect 6852 -7036 6884 -7034
rect 6852 -7166 6884 -7164
rect 6852 -7194 6854 -7166
rect 6854 -7194 6882 -7166
rect 6882 -7194 6884 -7166
rect 6852 -7196 6884 -7194
rect 6852 -7326 6884 -7324
rect 6852 -7354 6854 -7326
rect 6854 -7354 6882 -7326
rect 6882 -7354 6884 -7326
rect 6852 -7356 6884 -7354
rect 6852 -7486 6884 -7484
rect 6852 -7514 6854 -7486
rect 6854 -7514 6882 -7486
rect 6882 -7514 6884 -7486
rect 6852 -7516 6884 -7514
rect 6852 -7646 6884 -7644
rect 6852 -7674 6854 -7646
rect 6854 -7674 6882 -7646
rect 6882 -7674 6884 -7646
rect 6852 -7676 6884 -7674
rect 6852 -7806 6884 -7804
rect 6852 -7834 6854 -7806
rect 6854 -7834 6882 -7806
rect 6882 -7834 6884 -7806
rect 6852 -7836 6884 -7834
rect 6852 -7966 6884 -7964
rect 6852 -7994 6854 -7966
rect 6854 -7994 6882 -7966
rect 6882 -7994 6884 -7966
rect 6852 -7996 6884 -7994
rect 6852 -8126 6884 -8124
rect 6852 -8154 6854 -8126
rect 6854 -8154 6882 -8126
rect 6882 -8154 6884 -8126
rect 6852 -8156 6884 -8154
rect 6852 -8286 6884 -8284
rect 6852 -8314 6854 -8286
rect 6854 -8314 6882 -8286
rect 6882 -8314 6884 -8286
rect 6852 -8316 6884 -8314
rect 6852 -8446 6884 -8444
rect 6852 -8474 6854 -8446
rect 6854 -8474 6882 -8446
rect 6882 -8474 6884 -8446
rect 6852 -8476 6884 -8474
rect 6852 -8606 6884 -8604
rect 6852 -8634 6854 -8606
rect 6854 -8634 6882 -8606
rect 6882 -8634 6884 -8606
rect 6852 -8636 6884 -8634
rect 6852 -8766 6884 -8764
rect 6852 -8794 6854 -8766
rect 6854 -8794 6882 -8766
rect 6882 -8794 6884 -8766
rect 6852 -8796 6884 -8794
rect 6852 -8926 6884 -8924
rect 6852 -8954 6854 -8926
rect 6854 -8954 6882 -8926
rect 6882 -8954 6884 -8926
rect 6852 -8956 6884 -8954
rect 6852 -9086 6884 -9084
rect 6852 -9114 6854 -9086
rect 6854 -9114 6882 -9086
rect 6882 -9114 6884 -9086
rect 6852 -9116 6884 -9114
rect 3119 -9246 3151 -9244
rect 3119 -9274 3121 -9246
rect 3121 -9274 3149 -9246
rect 3149 -9274 3151 -9246
rect 3119 -9276 3151 -9274
rect 6852 -9246 6884 -9244
rect 6852 -9274 6854 -9246
rect 6854 -9274 6882 -9246
rect 6882 -9274 6884 -9246
rect 6852 -9276 6884 -9274
rect 3304 -9351 3336 -9349
rect 3304 -9379 3306 -9351
rect 3306 -9379 3334 -9351
rect 3334 -9379 3336 -9351
rect 3304 -9381 3336 -9379
rect 3464 -9351 3496 -9349
rect 3464 -9379 3466 -9351
rect 3466 -9379 3494 -9351
rect 3494 -9379 3496 -9351
rect 3464 -9381 3496 -9379
rect 3624 -9351 3656 -9349
rect 3624 -9379 3626 -9351
rect 3626 -9379 3654 -9351
rect 3654 -9379 3656 -9351
rect 3624 -9381 3656 -9379
rect 3784 -9351 3816 -9349
rect 3784 -9379 3786 -9351
rect 3786 -9379 3814 -9351
rect 3814 -9379 3816 -9351
rect 3784 -9381 3816 -9379
rect 3944 -9351 3976 -9349
rect 3944 -9379 3946 -9351
rect 3946 -9379 3974 -9351
rect 3974 -9379 3976 -9351
rect 3944 -9381 3976 -9379
rect 4104 -9351 4136 -9349
rect 4104 -9379 4106 -9351
rect 4106 -9379 4134 -9351
rect 4134 -9379 4136 -9351
rect 4104 -9381 4136 -9379
rect 4264 -9351 4296 -9349
rect 4264 -9379 4266 -9351
rect 4266 -9379 4294 -9351
rect 4294 -9379 4296 -9351
rect 4264 -9381 4296 -9379
rect 4424 -9351 4456 -9349
rect 4424 -9379 4426 -9351
rect 4426 -9379 4454 -9351
rect 4454 -9379 4456 -9351
rect 4424 -9381 4456 -9379
rect 4584 -9351 4616 -9349
rect 4584 -9379 4586 -9351
rect 4586 -9379 4614 -9351
rect 4614 -9379 4616 -9351
rect 4584 -9381 4616 -9379
rect 4744 -9351 4776 -9349
rect 4744 -9379 4746 -9351
rect 4746 -9379 4774 -9351
rect 4774 -9379 4776 -9351
rect 4744 -9381 4776 -9379
rect 4904 -9351 4936 -9349
rect 4904 -9379 4906 -9351
rect 4906 -9379 4934 -9351
rect 4934 -9379 4936 -9351
rect 4904 -9381 4936 -9379
rect 5064 -9351 5096 -9349
rect 5064 -9379 5066 -9351
rect 5066 -9379 5094 -9351
rect 5094 -9379 5096 -9351
rect 5064 -9381 5096 -9379
rect 5224 -9351 5256 -9349
rect 5224 -9379 5226 -9351
rect 5226 -9379 5254 -9351
rect 5254 -9379 5256 -9351
rect 5224 -9381 5256 -9379
rect 5384 -9351 5416 -9349
rect 5384 -9379 5386 -9351
rect 5386 -9379 5414 -9351
rect 5414 -9379 5416 -9351
rect 5384 -9381 5416 -9379
rect 5544 -9351 5576 -9349
rect 5544 -9379 5546 -9351
rect 5546 -9379 5574 -9351
rect 5574 -9379 5576 -9351
rect 5544 -9381 5576 -9379
rect 5704 -9351 5736 -9349
rect 5704 -9379 5706 -9351
rect 5706 -9379 5734 -9351
rect 5734 -9379 5736 -9351
rect 5704 -9381 5736 -9379
rect 5864 -9351 5896 -9349
rect 5864 -9379 5866 -9351
rect 5866 -9379 5894 -9351
rect 5894 -9379 5896 -9351
rect 5864 -9381 5896 -9379
rect 6024 -9351 6056 -9349
rect 6024 -9379 6026 -9351
rect 6026 -9379 6054 -9351
rect 6054 -9379 6056 -9351
rect 6024 -9381 6056 -9379
rect 6184 -9351 6216 -9349
rect 6184 -9379 6186 -9351
rect 6186 -9379 6214 -9351
rect 6214 -9379 6216 -9351
rect 6184 -9381 6216 -9379
rect 6344 -9351 6376 -9349
rect 6344 -9379 6346 -9351
rect 6346 -9379 6374 -9351
rect 6374 -9379 6376 -9351
rect 6344 -9381 6376 -9379
rect 6504 -9351 6536 -9349
rect 6504 -9379 6506 -9351
rect 6506 -9379 6534 -9351
rect 6534 -9379 6536 -9351
rect 6504 -9381 6536 -9379
rect 6664 -9351 6696 -9349
rect 6664 -9379 6666 -9351
rect 6666 -9379 6694 -9351
rect 6694 -9379 6696 -9351
rect 6664 -9381 6696 -9379
rect 3304 -11623 3336 -11621
rect 3304 -11651 3306 -11623
rect 3306 -11651 3334 -11623
rect 3334 -11651 3336 -11623
rect 3304 -11653 3336 -11651
rect 3464 -11623 3496 -11621
rect 3464 -11651 3466 -11623
rect 3466 -11651 3494 -11623
rect 3494 -11651 3496 -11623
rect 3464 -11653 3496 -11651
rect 3624 -11623 3656 -11621
rect 3624 -11651 3626 -11623
rect 3626 -11651 3654 -11623
rect 3654 -11651 3656 -11623
rect 3624 -11653 3656 -11651
rect 3784 -11623 3816 -11621
rect 3784 -11651 3786 -11623
rect 3786 -11651 3814 -11623
rect 3814 -11651 3816 -11623
rect 3784 -11653 3816 -11651
rect 3944 -11623 3976 -11621
rect 3944 -11651 3946 -11623
rect 3946 -11651 3974 -11623
rect 3974 -11651 3976 -11623
rect 3944 -11653 3976 -11651
rect 4104 -11623 4136 -11621
rect 4104 -11651 4106 -11623
rect 4106 -11651 4134 -11623
rect 4134 -11651 4136 -11623
rect 4104 -11653 4136 -11651
rect 4264 -11623 4296 -11621
rect 4264 -11651 4266 -11623
rect 4266 -11651 4294 -11623
rect 4294 -11651 4296 -11623
rect 4264 -11653 4296 -11651
rect 4424 -11623 4456 -11621
rect 4424 -11651 4426 -11623
rect 4426 -11651 4454 -11623
rect 4454 -11651 4456 -11623
rect 4424 -11653 4456 -11651
rect 4584 -11623 4616 -11621
rect 4584 -11651 4586 -11623
rect 4586 -11651 4614 -11623
rect 4614 -11651 4616 -11623
rect 4584 -11653 4616 -11651
rect 4744 -11623 4776 -11621
rect 4744 -11651 4746 -11623
rect 4746 -11651 4774 -11623
rect 4774 -11651 4776 -11623
rect 4744 -11653 4776 -11651
rect 4904 -11623 4936 -11621
rect 4904 -11651 4906 -11623
rect 4906 -11651 4934 -11623
rect 4934 -11651 4936 -11623
rect 4904 -11653 4936 -11651
rect 5064 -11623 5096 -11621
rect 5064 -11651 5066 -11623
rect 5066 -11651 5094 -11623
rect 5094 -11651 5096 -11623
rect 5064 -11653 5096 -11651
rect 5224 -11623 5256 -11621
rect 5224 -11651 5226 -11623
rect 5226 -11651 5254 -11623
rect 5254 -11651 5256 -11623
rect 5224 -11653 5256 -11651
rect 5384 -11623 5416 -11621
rect 5384 -11651 5386 -11623
rect 5386 -11651 5414 -11623
rect 5414 -11651 5416 -11623
rect 5384 -11653 5416 -11651
rect 5544 -11623 5576 -11621
rect 5544 -11651 5546 -11623
rect 5546 -11651 5574 -11623
rect 5574 -11651 5576 -11623
rect 5544 -11653 5576 -11651
rect 5704 -11623 5736 -11621
rect 5704 -11651 5706 -11623
rect 5706 -11651 5734 -11623
rect 5734 -11651 5736 -11623
rect 5704 -11653 5736 -11651
rect 5864 -11623 5896 -11621
rect 5864 -11651 5866 -11623
rect 5866 -11651 5894 -11623
rect 5894 -11651 5896 -11623
rect 5864 -11653 5896 -11651
rect 6024 -11623 6056 -11621
rect 6024 -11651 6026 -11623
rect 6026 -11651 6054 -11623
rect 6054 -11651 6056 -11623
rect 6024 -11653 6056 -11651
rect 6184 -11623 6216 -11621
rect 6184 -11651 6186 -11623
rect 6186 -11651 6214 -11623
rect 6214 -11651 6216 -11623
rect 6184 -11653 6216 -11651
rect 6344 -11623 6376 -11621
rect 6344 -11651 6346 -11623
rect 6346 -11651 6374 -11623
rect 6374 -11651 6376 -11623
rect 6344 -11653 6376 -11651
rect 6504 -11623 6536 -11621
rect 6504 -11651 6506 -11623
rect 6506 -11651 6534 -11623
rect 6534 -11651 6536 -11623
rect 6504 -11653 6536 -11651
rect 6664 -11623 6696 -11621
rect 6664 -11651 6666 -11623
rect 6666 -11651 6694 -11623
rect 6694 -11651 6696 -11623
rect 6664 -11653 6696 -11651
rect 3119 -11726 3151 -11724
rect 3119 -11754 3121 -11726
rect 3121 -11754 3149 -11726
rect 3149 -11754 3151 -11726
rect 3119 -11756 3151 -11754
rect 6852 -11726 6884 -11724
rect 6852 -11754 6854 -11726
rect 6854 -11754 6882 -11726
rect 6882 -11754 6884 -11726
rect 6852 -11756 6884 -11754
rect 3119 -11886 3151 -11884
rect 3119 -11914 3121 -11886
rect 3121 -11914 3149 -11886
rect 3149 -11914 3151 -11886
rect 3119 -11916 3151 -11914
rect 3119 -12046 3151 -12044
rect 3119 -12074 3121 -12046
rect 3121 -12074 3149 -12046
rect 3149 -12074 3151 -12046
rect 3119 -12076 3151 -12074
rect 3119 -12206 3151 -12204
rect 3119 -12234 3121 -12206
rect 3121 -12234 3149 -12206
rect 3149 -12234 3151 -12206
rect 3119 -12236 3151 -12234
rect 3119 -12366 3151 -12364
rect 3119 -12394 3121 -12366
rect 3121 -12394 3149 -12366
rect 3149 -12394 3151 -12366
rect 3119 -12396 3151 -12394
rect 3119 -12526 3151 -12524
rect 3119 -12554 3121 -12526
rect 3121 -12554 3149 -12526
rect 3149 -12554 3151 -12526
rect 3119 -12556 3151 -12554
rect 3119 -12686 3151 -12684
rect 3119 -12714 3121 -12686
rect 3121 -12714 3149 -12686
rect 3149 -12714 3151 -12686
rect 3119 -12716 3151 -12714
rect 3119 -12846 3151 -12844
rect 3119 -12874 3121 -12846
rect 3121 -12874 3149 -12846
rect 3149 -12874 3151 -12846
rect 3119 -12876 3151 -12874
rect 3119 -13006 3151 -13004
rect 3119 -13034 3121 -13006
rect 3121 -13034 3149 -13006
rect 3149 -13034 3151 -13006
rect 3119 -13036 3151 -13034
rect 3119 -13166 3151 -13164
rect 3119 -13194 3121 -13166
rect 3121 -13194 3149 -13166
rect 3149 -13194 3151 -13166
rect 3119 -13196 3151 -13194
rect 3119 -13326 3151 -13324
rect 3119 -13354 3121 -13326
rect 3121 -13354 3149 -13326
rect 3149 -13354 3151 -13326
rect 3119 -13356 3151 -13354
rect 3119 -13486 3151 -13484
rect 3119 -13514 3121 -13486
rect 3121 -13514 3149 -13486
rect 3149 -13514 3151 -13486
rect 3119 -13516 3151 -13514
rect 3119 -13646 3151 -13644
rect 3119 -13674 3121 -13646
rect 3121 -13674 3149 -13646
rect 3149 -13674 3151 -13646
rect 3119 -13676 3151 -13674
rect 3119 -13806 3151 -13804
rect 3119 -13834 3121 -13806
rect 3121 -13834 3149 -13806
rect 3149 -13834 3151 -13806
rect 3119 -13836 3151 -13834
rect 3119 -13966 3151 -13964
rect 3119 -13994 3121 -13966
rect 3121 -13994 3149 -13966
rect 3149 -13994 3151 -13966
rect 3119 -13996 3151 -13994
rect 3119 -14126 3151 -14124
rect 3119 -14154 3121 -14126
rect 3121 -14154 3149 -14126
rect 3149 -14154 3151 -14126
rect 3119 -14156 3151 -14154
rect 3119 -14286 3151 -14284
rect 3119 -14314 3121 -14286
rect 3121 -14314 3149 -14286
rect 3149 -14314 3151 -14286
rect 3119 -14316 3151 -14314
rect 3119 -14446 3151 -14444
rect 3119 -14474 3121 -14446
rect 3121 -14474 3149 -14446
rect 3149 -14474 3151 -14446
rect 3119 -14476 3151 -14474
rect 3119 -14606 3151 -14604
rect 3119 -14634 3121 -14606
rect 3121 -14634 3149 -14606
rect 3149 -14634 3151 -14606
rect 3119 -14636 3151 -14634
rect 3119 -14766 3151 -14764
rect 3119 -14794 3121 -14766
rect 3121 -14794 3149 -14766
rect 3149 -14794 3151 -14766
rect 3119 -14796 3151 -14794
rect 3119 -14926 3151 -14924
rect 3119 -14954 3121 -14926
rect 3121 -14954 3149 -14926
rect 3149 -14954 3151 -14926
rect 3119 -14956 3151 -14954
rect 3119 -15086 3151 -15084
rect 3119 -15114 3121 -15086
rect 3121 -15114 3149 -15086
rect 3149 -15114 3151 -15086
rect 3119 -15116 3151 -15114
rect 6852 -11886 6884 -11884
rect 6852 -11914 6854 -11886
rect 6854 -11914 6882 -11886
rect 6882 -11914 6884 -11886
rect 6852 -11916 6884 -11914
rect 6852 -12046 6884 -12044
rect 6852 -12074 6854 -12046
rect 6854 -12074 6882 -12046
rect 6882 -12074 6884 -12046
rect 6852 -12076 6884 -12074
rect 6852 -12206 6884 -12204
rect 6852 -12234 6854 -12206
rect 6854 -12234 6882 -12206
rect 6882 -12234 6884 -12206
rect 6852 -12236 6884 -12234
rect 6852 -12366 6884 -12364
rect 6852 -12394 6854 -12366
rect 6854 -12394 6882 -12366
rect 6882 -12394 6884 -12366
rect 6852 -12396 6884 -12394
rect 6852 -12526 6884 -12524
rect 6852 -12554 6854 -12526
rect 6854 -12554 6882 -12526
rect 6882 -12554 6884 -12526
rect 6852 -12556 6884 -12554
rect 6852 -12686 6884 -12684
rect 6852 -12714 6854 -12686
rect 6854 -12714 6882 -12686
rect 6882 -12714 6884 -12686
rect 6852 -12716 6884 -12714
rect 6852 -12846 6884 -12844
rect 6852 -12874 6854 -12846
rect 6854 -12874 6882 -12846
rect 6882 -12874 6884 -12846
rect 6852 -12876 6884 -12874
rect 9304 -5623 9336 -5621
rect 9304 -5651 9306 -5623
rect 9306 -5651 9334 -5623
rect 9334 -5651 9336 -5623
rect 9304 -5653 9336 -5651
rect 9464 -5623 9496 -5621
rect 9464 -5651 9466 -5623
rect 9466 -5651 9494 -5623
rect 9494 -5651 9496 -5623
rect 9464 -5653 9496 -5651
rect 9624 -5623 9656 -5621
rect 9624 -5651 9626 -5623
rect 9626 -5651 9654 -5623
rect 9654 -5651 9656 -5623
rect 9624 -5653 9656 -5651
rect 9784 -5623 9816 -5621
rect 9784 -5651 9786 -5623
rect 9786 -5651 9814 -5623
rect 9814 -5651 9816 -5623
rect 9784 -5653 9816 -5651
rect 9944 -5623 9976 -5621
rect 9944 -5651 9946 -5623
rect 9946 -5651 9974 -5623
rect 9974 -5651 9976 -5623
rect 9944 -5653 9976 -5651
rect 10104 -5623 10136 -5621
rect 10104 -5651 10106 -5623
rect 10106 -5651 10134 -5623
rect 10134 -5651 10136 -5623
rect 10104 -5653 10136 -5651
rect 10264 -5623 10296 -5621
rect 10264 -5651 10266 -5623
rect 10266 -5651 10294 -5623
rect 10294 -5651 10296 -5623
rect 10264 -5653 10296 -5651
rect 10424 -5623 10456 -5621
rect 10424 -5651 10426 -5623
rect 10426 -5651 10454 -5623
rect 10454 -5651 10456 -5623
rect 10424 -5653 10456 -5651
rect 10584 -5623 10616 -5621
rect 10584 -5651 10586 -5623
rect 10586 -5651 10614 -5623
rect 10614 -5651 10616 -5623
rect 10584 -5653 10616 -5651
rect 10744 -5623 10776 -5621
rect 10744 -5651 10746 -5623
rect 10746 -5651 10774 -5623
rect 10774 -5651 10776 -5623
rect 10744 -5653 10776 -5651
rect 10904 -5623 10936 -5621
rect 10904 -5651 10906 -5623
rect 10906 -5651 10934 -5623
rect 10934 -5651 10936 -5623
rect 10904 -5653 10936 -5651
rect 11064 -5623 11096 -5621
rect 11064 -5651 11066 -5623
rect 11066 -5651 11094 -5623
rect 11094 -5651 11096 -5623
rect 11064 -5653 11096 -5651
rect 11224 -5623 11256 -5621
rect 11224 -5651 11226 -5623
rect 11226 -5651 11254 -5623
rect 11254 -5651 11256 -5623
rect 11224 -5653 11256 -5651
rect 11384 -5623 11416 -5621
rect 11384 -5651 11386 -5623
rect 11386 -5651 11414 -5623
rect 11414 -5651 11416 -5623
rect 11384 -5653 11416 -5651
rect 11544 -5623 11576 -5621
rect 11544 -5651 11546 -5623
rect 11546 -5651 11574 -5623
rect 11574 -5651 11576 -5623
rect 11544 -5653 11576 -5651
rect 11704 -5623 11736 -5621
rect 11704 -5651 11706 -5623
rect 11706 -5651 11734 -5623
rect 11734 -5651 11736 -5623
rect 11704 -5653 11736 -5651
rect 11864 -5623 11896 -5621
rect 11864 -5651 11866 -5623
rect 11866 -5651 11894 -5623
rect 11894 -5651 11896 -5623
rect 11864 -5653 11896 -5651
rect 12024 -5623 12056 -5621
rect 12024 -5651 12026 -5623
rect 12026 -5651 12054 -5623
rect 12054 -5651 12056 -5623
rect 12024 -5653 12056 -5651
rect 12184 -5623 12216 -5621
rect 12184 -5651 12186 -5623
rect 12186 -5651 12214 -5623
rect 12214 -5651 12216 -5623
rect 12184 -5653 12216 -5651
rect 12344 -5623 12376 -5621
rect 12344 -5651 12346 -5623
rect 12346 -5651 12374 -5623
rect 12374 -5651 12376 -5623
rect 12344 -5653 12376 -5651
rect 12504 -5623 12536 -5621
rect 12504 -5651 12506 -5623
rect 12506 -5651 12534 -5623
rect 12534 -5651 12536 -5623
rect 12504 -5653 12536 -5651
rect 12664 -5623 12696 -5621
rect 12664 -5651 12666 -5623
rect 12666 -5651 12694 -5623
rect 12694 -5651 12696 -5623
rect 12664 -5653 12696 -5651
rect 9119 -5726 9151 -5724
rect 9119 -5754 9121 -5726
rect 9121 -5754 9149 -5726
rect 9149 -5754 9151 -5726
rect 9119 -5756 9151 -5754
rect 12852 -5726 12884 -5724
rect 12852 -5754 12854 -5726
rect 12854 -5754 12882 -5726
rect 12882 -5754 12884 -5726
rect 12852 -5756 12884 -5754
rect 9119 -5886 9151 -5884
rect 9119 -5914 9121 -5886
rect 9121 -5914 9149 -5886
rect 9149 -5914 9151 -5886
rect 9119 -5916 9151 -5914
rect 9119 -6046 9151 -6044
rect 9119 -6074 9121 -6046
rect 9121 -6074 9149 -6046
rect 9149 -6074 9151 -6046
rect 9119 -6076 9151 -6074
rect 9119 -6206 9151 -6204
rect 9119 -6234 9121 -6206
rect 9121 -6234 9149 -6206
rect 9149 -6234 9151 -6206
rect 9119 -6236 9151 -6234
rect 9119 -6366 9151 -6364
rect 9119 -6394 9121 -6366
rect 9121 -6394 9149 -6366
rect 9149 -6394 9151 -6366
rect 9119 -6396 9151 -6394
rect 9119 -6526 9151 -6524
rect 9119 -6554 9121 -6526
rect 9121 -6554 9149 -6526
rect 9149 -6554 9151 -6526
rect 9119 -6556 9151 -6554
rect 9119 -6686 9151 -6684
rect 9119 -6714 9121 -6686
rect 9121 -6714 9149 -6686
rect 9149 -6714 9151 -6686
rect 9119 -6716 9151 -6714
rect 9119 -6846 9151 -6844
rect 9119 -6874 9121 -6846
rect 9121 -6874 9149 -6846
rect 9149 -6874 9151 -6846
rect 9119 -6876 9151 -6874
rect 9119 -7006 9151 -7004
rect 9119 -7034 9121 -7006
rect 9121 -7034 9149 -7006
rect 9149 -7034 9151 -7006
rect 9119 -7036 9151 -7034
rect 9119 -7166 9151 -7164
rect 9119 -7194 9121 -7166
rect 9121 -7194 9149 -7166
rect 9149 -7194 9151 -7166
rect 9119 -7196 9151 -7194
rect 9119 -7326 9151 -7324
rect 9119 -7354 9121 -7326
rect 9121 -7354 9149 -7326
rect 9149 -7354 9151 -7326
rect 9119 -7356 9151 -7354
rect 9119 -7486 9151 -7484
rect 9119 -7514 9121 -7486
rect 9121 -7514 9149 -7486
rect 9149 -7514 9151 -7486
rect 9119 -7516 9151 -7514
rect 9119 -7646 9151 -7644
rect 9119 -7674 9121 -7646
rect 9121 -7674 9149 -7646
rect 9149 -7674 9151 -7646
rect 9119 -7676 9151 -7674
rect 9119 -7806 9151 -7804
rect 9119 -7834 9121 -7806
rect 9121 -7834 9149 -7806
rect 9149 -7834 9151 -7806
rect 9119 -7836 9151 -7834
rect 9119 -7966 9151 -7964
rect 9119 -7994 9121 -7966
rect 9121 -7994 9149 -7966
rect 9149 -7994 9151 -7966
rect 9119 -7996 9151 -7994
rect 9119 -8126 9151 -8124
rect 9119 -8154 9121 -8126
rect 9121 -8154 9149 -8126
rect 9149 -8154 9151 -8126
rect 9119 -8156 9151 -8154
rect 9119 -8286 9151 -8284
rect 9119 -8314 9121 -8286
rect 9121 -8314 9149 -8286
rect 9149 -8314 9151 -8286
rect 9119 -8316 9151 -8314
rect 9119 -8446 9151 -8444
rect 9119 -8474 9121 -8446
rect 9121 -8474 9149 -8446
rect 9149 -8474 9151 -8446
rect 9119 -8476 9151 -8474
rect 9119 -8606 9151 -8604
rect 9119 -8634 9121 -8606
rect 9121 -8634 9149 -8606
rect 9149 -8634 9151 -8606
rect 9119 -8636 9151 -8634
rect 9119 -8766 9151 -8764
rect 9119 -8794 9121 -8766
rect 9121 -8794 9149 -8766
rect 9149 -8794 9151 -8766
rect 9119 -8796 9151 -8794
rect 9119 -8926 9151 -8924
rect 9119 -8954 9121 -8926
rect 9121 -8954 9149 -8926
rect 9149 -8954 9151 -8926
rect 9119 -8956 9151 -8954
rect 9119 -9086 9151 -9084
rect 9119 -9114 9121 -9086
rect 9121 -9114 9149 -9086
rect 9149 -9114 9151 -9086
rect 9119 -9116 9151 -9114
rect 12852 -5886 12884 -5884
rect 12852 -5914 12854 -5886
rect 12854 -5914 12882 -5886
rect 12882 -5914 12884 -5886
rect 12852 -5916 12884 -5914
rect 12852 -6046 12884 -6044
rect 12852 -6074 12854 -6046
rect 12854 -6074 12882 -6046
rect 12882 -6074 12884 -6046
rect 12852 -6076 12884 -6074
rect 12852 -6206 12884 -6204
rect 12852 -6234 12854 -6206
rect 12854 -6234 12882 -6206
rect 12882 -6234 12884 -6206
rect 12852 -6236 12884 -6234
rect 12852 -6366 12884 -6364
rect 12852 -6394 12854 -6366
rect 12854 -6394 12882 -6366
rect 12882 -6394 12884 -6366
rect 12852 -6396 12884 -6394
rect 12852 -6526 12884 -6524
rect 12852 -6554 12854 -6526
rect 12854 -6554 12882 -6526
rect 12882 -6554 12884 -6526
rect 12852 -6556 12884 -6554
rect 12852 -6686 12884 -6684
rect 12852 -6714 12854 -6686
rect 12854 -6714 12882 -6686
rect 12882 -6714 12884 -6686
rect 12852 -6716 12884 -6714
rect 12852 -6846 12884 -6844
rect 12852 -6874 12854 -6846
rect 12854 -6874 12882 -6846
rect 12882 -6874 12884 -6846
rect 12852 -6876 12884 -6874
rect 12852 -7006 12884 -7004
rect 12852 -7034 12854 -7006
rect 12854 -7034 12882 -7006
rect 12882 -7034 12884 -7006
rect 12852 -7036 12884 -7034
rect 12852 -7166 12884 -7164
rect 12852 -7194 12854 -7166
rect 12854 -7194 12882 -7166
rect 12882 -7194 12884 -7166
rect 12852 -7196 12884 -7194
rect 12852 -7326 12884 -7324
rect 12852 -7354 12854 -7326
rect 12854 -7354 12882 -7326
rect 12882 -7354 12884 -7326
rect 12852 -7356 12884 -7354
rect 12852 -7486 12884 -7484
rect 12852 -7514 12854 -7486
rect 12854 -7514 12882 -7486
rect 12882 -7514 12884 -7486
rect 12852 -7516 12884 -7514
rect 12852 -7646 12884 -7644
rect 12852 -7674 12854 -7646
rect 12854 -7674 12882 -7646
rect 12882 -7674 12884 -7646
rect 12852 -7676 12884 -7674
rect 12852 -7806 12884 -7804
rect 12852 -7834 12854 -7806
rect 12854 -7834 12882 -7806
rect 12882 -7834 12884 -7806
rect 12852 -7836 12884 -7834
rect 15304 -5623 15336 -5621
rect 15304 -5651 15306 -5623
rect 15306 -5651 15334 -5623
rect 15334 -5651 15336 -5623
rect 15304 -5653 15336 -5651
rect 15464 -5623 15496 -5621
rect 15464 -5651 15466 -5623
rect 15466 -5651 15494 -5623
rect 15494 -5651 15496 -5623
rect 15464 -5653 15496 -5651
rect 15624 -5623 15656 -5621
rect 15624 -5651 15626 -5623
rect 15626 -5651 15654 -5623
rect 15654 -5651 15656 -5623
rect 15624 -5653 15656 -5651
rect 15784 -5623 15816 -5621
rect 15784 -5651 15786 -5623
rect 15786 -5651 15814 -5623
rect 15814 -5651 15816 -5623
rect 15784 -5653 15816 -5651
rect 15944 -5623 15976 -5621
rect 15944 -5651 15946 -5623
rect 15946 -5651 15974 -5623
rect 15974 -5651 15976 -5623
rect 15944 -5653 15976 -5651
rect 16104 -5623 16136 -5621
rect 16104 -5651 16106 -5623
rect 16106 -5651 16134 -5623
rect 16134 -5651 16136 -5623
rect 16104 -5653 16136 -5651
rect 16264 -5623 16296 -5621
rect 16264 -5651 16266 -5623
rect 16266 -5651 16294 -5623
rect 16294 -5651 16296 -5623
rect 16264 -5653 16296 -5651
rect 16424 -5623 16456 -5621
rect 16424 -5651 16426 -5623
rect 16426 -5651 16454 -5623
rect 16454 -5651 16456 -5623
rect 16424 -5653 16456 -5651
rect 16584 -5623 16616 -5621
rect 16584 -5651 16586 -5623
rect 16586 -5651 16614 -5623
rect 16614 -5651 16616 -5623
rect 16584 -5653 16616 -5651
rect 16744 -5623 16776 -5621
rect 16744 -5651 16746 -5623
rect 16746 -5651 16774 -5623
rect 16774 -5651 16776 -5623
rect 16744 -5653 16776 -5651
rect 16904 -5623 16936 -5621
rect 16904 -5651 16906 -5623
rect 16906 -5651 16934 -5623
rect 16934 -5651 16936 -5623
rect 16904 -5653 16936 -5651
rect 17064 -5623 17096 -5621
rect 17064 -5651 17066 -5623
rect 17066 -5651 17094 -5623
rect 17094 -5651 17096 -5623
rect 17064 -5653 17096 -5651
rect 17224 -5623 17256 -5621
rect 17224 -5651 17226 -5623
rect 17226 -5651 17254 -5623
rect 17254 -5651 17256 -5623
rect 17224 -5653 17256 -5651
rect 17384 -5623 17416 -5621
rect 17384 -5651 17386 -5623
rect 17386 -5651 17414 -5623
rect 17414 -5651 17416 -5623
rect 17384 -5653 17416 -5651
rect 17544 -5623 17576 -5621
rect 17544 -5651 17546 -5623
rect 17546 -5651 17574 -5623
rect 17574 -5651 17576 -5623
rect 17544 -5653 17576 -5651
rect 17704 -5623 17736 -5621
rect 17704 -5651 17706 -5623
rect 17706 -5651 17734 -5623
rect 17734 -5651 17736 -5623
rect 17704 -5653 17736 -5651
rect 17864 -5623 17896 -5621
rect 17864 -5651 17866 -5623
rect 17866 -5651 17894 -5623
rect 17894 -5651 17896 -5623
rect 17864 -5653 17896 -5651
rect 18024 -5623 18056 -5621
rect 18024 -5651 18026 -5623
rect 18026 -5651 18054 -5623
rect 18054 -5651 18056 -5623
rect 18024 -5653 18056 -5651
rect 18184 -5623 18216 -5621
rect 18184 -5651 18186 -5623
rect 18186 -5651 18214 -5623
rect 18214 -5651 18216 -5623
rect 18184 -5653 18216 -5651
rect 18344 -5623 18376 -5621
rect 18344 -5651 18346 -5623
rect 18346 -5651 18374 -5623
rect 18374 -5651 18376 -5623
rect 18344 -5653 18376 -5651
rect 18504 -5623 18536 -5621
rect 18504 -5651 18506 -5623
rect 18506 -5651 18534 -5623
rect 18534 -5651 18536 -5623
rect 18504 -5653 18536 -5651
rect 18664 -5623 18696 -5621
rect 18664 -5651 18666 -5623
rect 18666 -5651 18694 -5623
rect 18694 -5651 18696 -5623
rect 18664 -5653 18696 -5651
rect 15119 -5726 15151 -5724
rect 15119 -5754 15121 -5726
rect 15121 -5754 15149 -5726
rect 15149 -5754 15151 -5726
rect 15119 -5756 15151 -5754
rect 18852 -5726 18884 -5724
rect 18852 -5754 18854 -5726
rect 18854 -5754 18882 -5726
rect 18882 -5754 18884 -5726
rect 18852 -5756 18884 -5754
rect 15119 -5886 15151 -5884
rect 15119 -5914 15121 -5886
rect 15121 -5914 15149 -5886
rect 15149 -5914 15151 -5886
rect 15119 -5916 15151 -5914
rect 15119 -6046 15151 -6044
rect 15119 -6074 15121 -6046
rect 15121 -6074 15149 -6046
rect 15149 -6074 15151 -6046
rect 15119 -6076 15151 -6074
rect 15119 -6206 15151 -6204
rect 15119 -6234 15121 -6206
rect 15121 -6234 15149 -6206
rect 15149 -6234 15151 -6206
rect 15119 -6236 15151 -6234
rect 15119 -6366 15151 -6364
rect 15119 -6394 15121 -6366
rect 15121 -6394 15149 -6366
rect 15149 -6394 15151 -6366
rect 15119 -6396 15151 -6394
rect 15119 -6526 15151 -6524
rect 15119 -6554 15121 -6526
rect 15121 -6554 15149 -6526
rect 15149 -6554 15151 -6526
rect 15119 -6556 15151 -6554
rect 15119 -6686 15151 -6684
rect 15119 -6714 15121 -6686
rect 15121 -6714 15149 -6686
rect 15149 -6714 15151 -6686
rect 15119 -6716 15151 -6714
rect 15119 -6846 15151 -6844
rect 15119 -6874 15121 -6846
rect 15121 -6874 15149 -6846
rect 15149 -6874 15151 -6846
rect 15119 -6876 15151 -6874
rect 15119 -7006 15151 -7004
rect 15119 -7034 15121 -7006
rect 15121 -7034 15149 -7006
rect 15149 -7034 15151 -7006
rect 15119 -7036 15151 -7034
rect 15119 -7166 15151 -7164
rect 15119 -7194 15121 -7166
rect 15121 -7194 15149 -7166
rect 15149 -7194 15151 -7166
rect 15119 -7196 15151 -7194
rect 15119 -7326 15151 -7324
rect 15119 -7354 15121 -7326
rect 15121 -7354 15149 -7326
rect 15149 -7354 15151 -7326
rect 15119 -7356 15151 -7354
rect 15119 -7486 15151 -7484
rect 15119 -7514 15121 -7486
rect 15121 -7514 15149 -7486
rect 15149 -7514 15151 -7486
rect 15119 -7516 15151 -7514
rect 15119 -7646 15151 -7644
rect 15119 -7674 15121 -7646
rect 15121 -7674 15149 -7646
rect 15149 -7674 15151 -7646
rect 15119 -7676 15151 -7674
rect 12852 -7966 12884 -7964
rect 12852 -7994 12854 -7966
rect 12854 -7994 12882 -7966
rect 12882 -7994 12884 -7966
rect 12852 -7996 12884 -7994
rect 12852 -8126 12884 -8124
rect 12852 -8154 12854 -8126
rect 12854 -8154 12882 -8126
rect 12882 -8154 12884 -8126
rect 12852 -8156 12884 -8154
rect 12852 -8286 12884 -8284
rect 12852 -8314 12854 -8286
rect 12854 -8314 12882 -8286
rect 12882 -8314 12884 -8286
rect 12852 -8316 12884 -8314
rect 12852 -8446 12884 -8444
rect 12852 -8474 12854 -8446
rect 12854 -8474 12882 -8446
rect 12882 -8474 12884 -8446
rect 12852 -8476 12884 -8474
rect 12852 -8606 12884 -8604
rect 12852 -8634 12854 -8606
rect 12854 -8634 12882 -8606
rect 12882 -8634 12884 -8606
rect 12852 -8636 12884 -8634
rect 12852 -8766 12884 -8764
rect 12852 -8794 12854 -8766
rect 12854 -8794 12882 -8766
rect 12882 -8794 12884 -8766
rect 12852 -8796 12884 -8794
rect 12852 -8926 12884 -8924
rect 12852 -8954 12854 -8926
rect 12854 -8954 12882 -8926
rect 12882 -8954 12884 -8926
rect 12852 -8956 12884 -8954
rect 12852 -9086 12884 -9084
rect 12852 -9114 12854 -9086
rect 12854 -9114 12882 -9086
rect 12882 -9114 12884 -9086
rect 12852 -9116 12884 -9114
rect 9119 -9246 9151 -9244
rect 9119 -9274 9121 -9246
rect 9121 -9274 9149 -9246
rect 9149 -9274 9151 -9246
rect 9119 -9276 9151 -9274
rect 12852 -9246 12884 -9244
rect 12852 -9274 12854 -9246
rect 12854 -9274 12882 -9246
rect 12882 -9274 12884 -9246
rect 12852 -9276 12884 -9274
rect 9304 -9351 9336 -9349
rect 9304 -9379 9306 -9351
rect 9306 -9379 9334 -9351
rect 9334 -9379 9336 -9351
rect 9304 -9381 9336 -9379
rect 9464 -9351 9496 -9349
rect 9464 -9379 9466 -9351
rect 9466 -9379 9494 -9351
rect 9494 -9379 9496 -9351
rect 9464 -9381 9496 -9379
rect 9624 -9351 9656 -9349
rect 9624 -9379 9626 -9351
rect 9626 -9379 9654 -9351
rect 9654 -9379 9656 -9351
rect 9624 -9381 9656 -9379
rect 9784 -9351 9816 -9349
rect 9784 -9379 9786 -9351
rect 9786 -9379 9814 -9351
rect 9814 -9379 9816 -9351
rect 9784 -9381 9816 -9379
rect 9944 -9351 9976 -9349
rect 9944 -9379 9946 -9351
rect 9946 -9379 9974 -9351
rect 9974 -9379 9976 -9351
rect 9944 -9381 9976 -9379
rect 10104 -9351 10136 -9349
rect 10104 -9379 10106 -9351
rect 10106 -9379 10134 -9351
rect 10134 -9379 10136 -9351
rect 10104 -9381 10136 -9379
rect 10264 -9351 10296 -9349
rect 10264 -9379 10266 -9351
rect 10266 -9379 10294 -9351
rect 10294 -9379 10296 -9351
rect 10264 -9381 10296 -9379
rect 10424 -9351 10456 -9349
rect 10424 -9379 10426 -9351
rect 10426 -9379 10454 -9351
rect 10454 -9379 10456 -9351
rect 10424 -9381 10456 -9379
rect 10584 -9351 10616 -9349
rect 10584 -9379 10586 -9351
rect 10586 -9379 10614 -9351
rect 10614 -9379 10616 -9351
rect 10584 -9381 10616 -9379
rect 10744 -9351 10776 -9349
rect 10744 -9379 10746 -9351
rect 10746 -9379 10774 -9351
rect 10774 -9379 10776 -9351
rect 10744 -9381 10776 -9379
rect 10904 -9351 10936 -9349
rect 10904 -9379 10906 -9351
rect 10906 -9379 10934 -9351
rect 10934 -9379 10936 -9351
rect 10904 -9381 10936 -9379
rect 11064 -9351 11096 -9349
rect 11064 -9379 11066 -9351
rect 11066 -9379 11094 -9351
rect 11094 -9379 11096 -9351
rect 11064 -9381 11096 -9379
rect 11224 -9351 11256 -9349
rect 11224 -9379 11226 -9351
rect 11226 -9379 11254 -9351
rect 11254 -9379 11256 -9351
rect 11224 -9381 11256 -9379
rect 11384 -9351 11416 -9349
rect 11384 -9379 11386 -9351
rect 11386 -9379 11414 -9351
rect 11414 -9379 11416 -9351
rect 11384 -9381 11416 -9379
rect 11544 -9351 11576 -9349
rect 11544 -9379 11546 -9351
rect 11546 -9379 11574 -9351
rect 11574 -9379 11576 -9351
rect 11544 -9381 11576 -9379
rect 11704 -9351 11736 -9349
rect 11704 -9379 11706 -9351
rect 11706 -9379 11734 -9351
rect 11734 -9379 11736 -9351
rect 11704 -9381 11736 -9379
rect 11864 -9351 11896 -9349
rect 11864 -9379 11866 -9351
rect 11866 -9379 11894 -9351
rect 11894 -9379 11896 -9351
rect 11864 -9381 11896 -9379
rect 12024 -9351 12056 -9349
rect 12024 -9379 12026 -9351
rect 12026 -9379 12054 -9351
rect 12054 -9379 12056 -9351
rect 12024 -9381 12056 -9379
rect 12184 -9351 12216 -9349
rect 12184 -9379 12186 -9351
rect 12186 -9379 12214 -9351
rect 12214 -9379 12216 -9351
rect 12184 -9381 12216 -9379
rect 12344 -9351 12376 -9349
rect 12344 -9379 12346 -9351
rect 12346 -9379 12374 -9351
rect 12374 -9379 12376 -9351
rect 12344 -9381 12376 -9379
rect 12504 -9351 12536 -9349
rect 12504 -9379 12506 -9351
rect 12506 -9379 12534 -9351
rect 12534 -9379 12536 -9351
rect 12504 -9381 12536 -9379
rect 12664 -9351 12696 -9349
rect 12664 -9379 12666 -9351
rect 12666 -9379 12694 -9351
rect 12694 -9379 12696 -9351
rect 12664 -9381 12696 -9379
rect 15119 -7806 15151 -7804
rect 15119 -7834 15121 -7806
rect 15121 -7834 15149 -7806
rect 15149 -7834 15151 -7806
rect 15119 -7836 15151 -7834
rect 15119 -7966 15151 -7964
rect 15119 -7994 15121 -7966
rect 15121 -7994 15149 -7966
rect 15149 -7994 15151 -7966
rect 15119 -7996 15151 -7994
rect 15119 -8126 15151 -8124
rect 15119 -8154 15121 -8126
rect 15121 -8154 15149 -8126
rect 15149 -8154 15151 -8126
rect 15119 -8156 15151 -8154
rect 15119 -8286 15151 -8284
rect 15119 -8314 15121 -8286
rect 15121 -8314 15149 -8286
rect 15149 -8314 15151 -8286
rect 15119 -8316 15151 -8314
rect 15119 -8446 15151 -8444
rect 15119 -8474 15121 -8446
rect 15121 -8474 15149 -8446
rect 15149 -8474 15151 -8446
rect 15119 -8476 15151 -8474
rect 15119 -8606 15151 -8604
rect 15119 -8634 15121 -8606
rect 15121 -8634 15149 -8606
rect 15149 -8634 15151 -8606
rect 15119 -8636 15151 -8634
rect 15119 -8766 15151 -8764
rect 15119 -8794 15121 -8766
rect 15121 -8794 15149 -8766
rect 15149 -8794 15151 -8766
rect 15119 -8796 15151 -8794
rect 15119 -8926 15151 -8924
rect 15119 -8954 15121 -8926
rect 15121 -8954 15149 -8926
rect 15149 -8954 15151 -8926
rect 15119 -8956 15151 -8954
rect 15119 -9086 15151 -9084
rect 15119 -9114 15121 -9086
rect 15121 -9114 15149 -9086
rect 15149 -9114 15151 -9086
rect 15119 -9116 15151 -9114
rect 18852 -5886 18884 -5884
rect 18852 -5914 18854 -5886
rect 18854 -5914 18882 -5886
rect 18882 -5914 18884 -5886
rect 18852 -5916 18884 -5914
rect 18852 -6046 18884 -6044
rect 18852 -6074 18854 -6046
rect 18854 -6074 18882 -6046
rect 18882 -6074 18884 -6046
rect 18852 -6076 18884 -6074
rect 18852 -6206 18884 -6204
rect 18852 -6234 18854 -6206
rect 18854 -6234 18882 -6206
rect 18882 -6234 18884 -6206
rect 18852 -6236 18884 -6234
rect 18852 -6366 18884 -6364
rect 18852 -6394 18854 -6366
rect 18854 -6394 18882 -6366
rect 18882 -6394 18884 -6366
rect 18852 -6396 18884 -6394
rect 18852 -6526 18884 -6524
rect 18852 -6554 18854 -6526
rect 18854 -6554 18882 -6526
rect 18882 -6554 18884 -6526
rect 18852 -6556 18884 -6554
rect 18852 -6686 18884 -6684
rect 18852 -6714 18854 -6686
rect 18854 -6714 18882 -6686
rect 18882 -6714 18884 -6686
rect 18852 -6716 18884 -6714
rect 18852 -6846 18884 -6844
rect 18852 -6874 18854 -6846
rect 18854 -6874 18882 -6846
rect 18882 -6874 18884 -6846
rect 18852 -6876 18884 -6874
rect 18852 -7006 18884 -7004
rect 18852 -7034 18854 -7006
rect 18854 -7034 18882 -7006
rect 18882 -7034 18884 -7006
rect 18852 -7036 18884 -7034
rect 18852 -7166 18884 -7164
rect 18852 -7194 18854 -7166
rect 18854 -7194 18882 -7166
rect 18882 -7194 18884 -7166
rect 18852 -7196 18884 -7194
rect 18852 -7326 18884 -7324
rect 18852 -7354 18854 -7326
rect 18854 -7354 18882 -7326
rect 18882 -7354 18884 -7326
rect 18852 -7356 18884 -7354
rect 18852 -7486 18884 -7484
rect 18852 -7514 18854 -7486
rect 18854 -7514 18882 -7486
rect 18882 -7514 18884 -7486
rect 18852 -7516 18884 -7514
rect 18852 -7646 18884 -7644
rect 18852 -7674 18854 -7646
rect 18854 -7674 18882 -7646
rect 18882 -7674 18884 -7646
rect 18852 -7676 18884 -7674
rect 18852 -7806 18884 -7804
rect 18852 -7834 18854 -7806
rect 18854 -7834 18882 -7806
rect 18882 -7834 18884 -7806
rect 18852 -7836 18884 -7834
rect 18852 -7966 18884 -7964
rect 18852 -7994 18854 -7966
rect 18854 -7994 18882 -7966
rect 18882 -7994 18884 -7966
rect 18852 -7996 18884 -7994
rect 18852 -8126 18884 -8124
rect 18852 -8154 18854 -8126
rect 18854 -8154 18882 -8126
rect 18882 -8154 18884 -8126
rect 18852 -8156 18884 -8154
rect 18852 -8286 18884 -8284
rect 18852 -8314 18854 -8286
rect 18854 -8314 18882 -8286
rect 18882 -8314 18884 -8286
rect 18852 -8316 18884 -8314
rect 18852 -8446 18884 -8444
rect 18852 -8474 18854 -8446
rect 18854 -8474 18882 -8446
rect 18882 -8474 18884 -8446
rect 18852 -8476 18884 -8474
rect 18852 -8606 18884 -8604
rect 18852 -8634 18854 -8606
rect 18854 -8634 18882 -8606
rect 18882 -8634 18884 -8606
rect 18852 -8636 18884 -8634
rect 18852 -8766 18884 -8764
rect 18852 -8794 18854 -8766
rect 18854 -8794 18882 -8766
rect 18882 -8794 18884 -8766
rect 18852 -8796 18884 -8794
rect 18852 -8926 18884 -8924
rect 18852 -8954 18854 -8926
rect 18854 -8954 18882 -8926
rect 18882 -8954 18884 -8926
rect 18852 -8956 18884 -8954
rect 18852 -9086 18884 -9084
rect 18852 -9114 18854 -9086
rect 18854 -9114 18882 -9086
rect 18882 -9114 18884 -9086
rect 18852 -9116 18884 -9114
rect 15119 -9246 15151 -9244
rect 15119 -9274 15121 -9246
rect 15121 -9274 15149 -9246
rect 15149 -9274 15151 -9246
rect 15119 -9276 15151 -9274
rect 18852 -9246 18884 -9244
rect 18852 -9274 18854 -9246
rect 18854 -9274 18882 -9246
rect 18882 -9274 18884 -9246
rect 18852 -9276 18884 -9274
rect 15304 -9351 15336 -9349
rect 15304 -9379 15306 -9351
rect 15306 -9379 15334 -9351
rect 15334 -9379 15336 -9351
rect 15304 -9381 15336 -9379
rect 15464 -9351 15496 -9349
rect 15464 -9379 15466 -9351
rect 15466 -9379 15494 -9351
rect 15494 -9379 15496 -9351
rect 15464 -9381 15496 -9379
rect 15624 -9351 15656 -9349
rect 15624 -9379 15626 -9351
rect 15626 -9379 15654 -9351
rect 15654 -9379 15656 -9351
rect 15624 -9381 15656 -9379
rect 15784 -9351 15816 -9349
rect 15784 -9379 15786 -9351
rect 15786 -9379 15814 -9351
rect 15814 -9379 15816 -9351
rect 15784 -9381 15816 -9379
rect 15944 -9351 15976 -9349
rect 15944 -9379 15946 -9351
rect 15946 -9379 15974 -9351
rect 15974 -9379 15976 -9351
rect 15944 -9381 15976 -9379
rect 16104 -9351 16136 -9349
rect 16104 -9379 16106 -9351
rect 16106 -9379 16134 -9351
rect 16134 -9379 16136 -9351
rect 16104 -9381 16136 -9379
rect 16264 -9351 16296 -9349
rect 16264 -9379 16266 -9351
rect 16266 -9379 16294 -9351
rect 16294 -9379 16296 -9351
rect 16264 -9381 16296 -9379
rect 16424 -9351 16456 -9349
rect 16424 -9379 16426 -9351
rect 16426 -9379 16454 -9351
rect 16454 -9379 16456 -9351
rect 16424 -9381 16456 -9379
rect 16584 -9351 16616 -9349
rect 16584 -9379 16586 -9351
rect 16586 -9379 16614 -9351
rect 16614 -9379 16616 -9351
rect 16584 -9381 16616 -9379
rect 16744 -9351 16776 -9349
rect 16744 -9379 16746 -9351
rect 16746 -9379 16774 -9351
rect 16774 -9379 16776 -9351
rect 16744 -9381 16776 -9379
rect 16904 -9351 16936 -9349
rect 16904 -9379 16906 -9351
rect 16906 -9379 16934 -9351
rect 16934 -9379 16936 -9351
rect 16904 -9381 16936 -9379
rect 17064 -9351 17096 -9349
rect 17064 -9379 17066 -9351
rect 17066 -9379 17094 -9351
rect 17094 -9379 17096 -9351
rect 17064 -9381 17096 -9379
rect 17224 -9351 17256 -9349
rect 17224 -9379 17226 -9351
rect 17226 -9379 17254 -9351
rect 17254 -9379 17256 -9351
rect 17224 -9381 17256 -9379
rect 17384 -9351 17416 -9349
rect 17384 -9379 17386 -9351
rect 17386 -9379 17414 -9351
rect 17414 -9379 17416 -9351
rect 17384 -9381 17416 -9379
rect 17544 -9351 17576 -9349
rect 17544 -9379 17546 -9351
rect 17546 -9379 17574 -9351
rect 17574 -9379 17576 -9351
rect 17544 -9381 17576 -9379
rect 17704 -9351 17736 -9349
rect 17704 -9379 17706 -9351
rect 17706 -9379 17734 -9351
rect 17734 -9379 17736 -9351
rect 17704 -9381 17736 -9379
rect 17864 -9351 17896 -9349
rect 17864 -9379 17866 -9351
rect 17866 -9379 17894 -9351
rect 17894 -9379 17896 -9351
rect 17864 -9381 17896 -9379
rect 18024 -9351 18056 -9349
rect 18024 -9379 18026 -9351
rect 18026 -9379 18054 -9351
rect 18054 -9379 18056 -9351
rect 18024 -9381 18056 -9379
rect 18184 -9351 18216 -9349
rect 18184 -9379 18186 -9351
rect 18186 -9379 18214 -9351
rect 18214 -9379 18216 -9351
rect 18184 -9381 18216 -9379
rect 18344 -9351 18376 -9349
rect 18344 -9379 18346 -9351
rect 18346 -9379 18374 -9351
rect 18374 -9379 18376 -9351
rect 18344 -9381 18376 -9379
rect 18504 -9351 18536 -9349
rect 18504 -9379 18506 -9351
rect 18506 -9379 18534 -9351
rect 18534 -9379 18536 -9351
rect 18504 -9381 18536 -9379
rect 18664 -9351 18696 -9349
rect 18664 -9379 18666 -9351
rect 18666 -9379 18694 -9351
rect 18694 -9379 18696 -9351
rect 18664 -9381 18696 -9379
rect 21304 -5623 21336 -5621
rect 21304 -5651 21306 -5623
rect 21306 -5651 21334 -5623
rect 21334 -5651 21336 -5623
rect 21304 -5653 21336 -5651
rect 21464 -5623 21496 -5621
rect 21464 -5651 21466 -5623
rect 21466 -5651 21494 -5623
rect 21494 -5651 21496 -5623
rect 21464 -5653 21496 -5651
rect 21624 -5623 21656 -5621
rect 21624 -5651 21626 -5623
rect 21626 -5651 21654 -5623
rect 21654 -5651 21656 -5623
rect 21624 -5653 21656 -5651
rect 21784 -5623 21816 -5621
rect 21784 -5651 21786 -5623
rect 21786 -5651 21814 -5623
rect 21814 -5651 21816 -5623
rect 21784 -5653 21816 -5651
rect 21944 -5623 21976 -5621
rect 21944 -5651 21946 -5623
rect 21946 -5651 21974 -5623
rect 21974 -5651 21976 -5623
rect 21944 -5653 21976 -5651
rect 22104 -5623 22136 -5621
rect 22104 -5651 22106 -5623
rect 22106 -5651 22134 -5623
rect 22134 -5651 22136 -5623
rect 22104 -5653 22136 -5651
rect 22264 -5623 22296 -5621
rect 22264 -5651 22266 -5623
rect 22266 -5651 22294 -5623
rect 22294 -5651 22296 -5623
rect 22264 -5653 22296 -5651
rect 22424 -5623 22456 -5621
rect 22424 -5651 22426 -5623
rect 22426 -5651 22454 -5623
rect 22454 -5651 22456 -5623
rect 22424 -5653 22456 -5651
rect 22584 -5623 22616 -5621
rect 22584 -5651 22586 -5623
rect 22586 -5651 22614 -5623
rect 22614 -5651 22616 -5623
rect 22584 -5653 22616 -5651
rect 22744 -5623 22776 -5621
rect 22744 -5651 22746 -5623
rect 22746 -5651 22774 -5623
rect 22774 -5651 22776 -5623
rect 22744 -5653 22776 -5651
rect 22904 -5623 22936 -5621
rect 22904 -5651 22906 -5623
rect 22906 -5651 22934 -5623
rect 22934 -5651 22936 -5623
rect 22904 -5653 22936 -5651
rect 23064 -5623 23096 -5621
rect 23064 -5651 23066 -5623
rect 23066 -5651 23094 -5623
rect 23094 -5651 23096 -5623
rect 23064 -5653 23096 -5651
rect 23224 -5623 23256 -5621
rect 23224 -5651 23226 -5623
rect 23226 -5651 23254 -5623
rect 23254 -5651 23256 -5623
rect 23224 -5653 23256 -5651
rect 23384 -5623 23416 -5621
rect 23384 -5651 23386 -5623
rect 23386 -5651 23414 -5623
rect 23414 -5651 23416 -5623
rect 23384 -5653 23416 -5651
rect 23544 -5623 23576 -5621
rect 23544 -5651 23546 -5623
rect 23546 -5651 23574 -5623
rect 23574 -5651 23576 -5623
rect 23544 -5653 23576 -5651
rect 23704 -5623 23736 -5621
rect 23704 -5651 23706 -5623
rect 23706 -5651 23734 -5623
rect 23734 -5651 23736 -5623
rect 23704 -5653 23736 -5651
rect 23864 -5623 23896 -5621
rect 23864 -5651 23866 -5623
rect 23866 -5651 23894 -5623
rect 23894 -5651 23896 -5623
rect 23864 -5653 23896 -5651
rect 24024 -5623 24056 -5621
rect 24024 -5651 24026 -5623
rect 24026 -5651 24054 -5623
rect 24054 -5651 24056 -5623
rect 24024 -5653 24056 -5651
rect 24184 -5623 24216 -5621
rect 24184 -5651 24186 -5623
rect 24186 -5651 24214 -5623
rect 24214 -5651 24216 -5623
rect 24184 -5653 24216 -5651
rect 24344 -5623 24376 -5621
rect 24344 -5651 24346 -5623
rect 24346 -5651 24374 -5623
rect 24374 -5651 24376 -5623
rect 24344 -5653 24376 -5651
rect 24504 -5623 24536 -5621
rect 24504 -5651 24506 -5623
rect 24506 -5651 24534 -5623
rect 24534 -5651 24536 -5623
rect 24504 -5653 24536 -5651
rect 24664 -5623 24696 -5621
rect 24664 -5651 24666 -5623
rect 24666 -5651 24694 -5623
rect 24694 -5651 24696 -5623
rect 24664 -5653 24696 -5651
rect 21119 -5726 21151 -5724
rect 21119 -5754 21121 -5726
rect 21121 -5754 21149 -5726
rect 21149 -5754 21151 -5726
rect 21119 -5756 21151 -5754
rect 24852 -5726 24884 -5724
rect 24852 -5754 24854 -5726
rect 24854 -5754 24882 -5726
rect 24882 -5754 24884 -5726
rect 24852 -5756 24884 -5754
rect 21119 -5886 21151 -5884
rect 21119 -5914 21121 -5886
rect 21121 -5914 21149 -5886
rect 21149 -5914 21151 -5886
rect 21119 -5916 21151 -5914
rect 21119 -6046 21151 -6044
rect 21119 -6074 21121 -6046
rect 21121 -6074 21149 -6046
rect 21149 -6074 21151 -6046
rect 21119 -6076 21151 -6074
rect 21119 -6206 21151 -6204
rect 21119 -6234 21121 -6206
rect 21121 -6234 21149 -6206
rect 21149 -6234 21151 -6206
rect 21119 -6236 21151 -6234
rect 21119 -6366 21151 -6364
rect 21119 -6394 21121 -6366
rect 21121 -6394 21149 -6366
rect 21149 -6394 21151 -6366
rect 21119 -6396 21151 -6394
rect 21119 -6526 21151 -6524
rect 21119 -6554 21121 -6526
rect 21121 -6554 21149 -6526
rect 21149 -6554 21151 -6526
rect 21119 -6556 21151 -6554
rect 21119 -6686 21151 -6684
rect 21119 -6714 21121 -6686
rect 21121 -6714 21149 -6686
rect 21149 -6714 21151 -6686
rect 21119 -6716 21151 -6714
rect 21119 -6846 21151 -6844
rect 21119 -6874 21121 -6846
rect 21121 -6874 21149 -6846
rect 21149 -6874 21151 -6846
rect 21119 -6876 21151 -6874
rect 21119 -7006 21151 -7004
rect 21119 -7034 21121 -7006
rect 21121 -7034 21149 -7006
rect 21149 -7034 21151 -7006
rect 21119 -7036 21151 -7034
rect 21119 -7166 21151 -7164
rect 21119 -7194 21121 -7166
rect 21121 -7194 21149 -7166
rect 21149 -7194 21151 -7166
rect 21119 -7196 21151 -7194
rect 21119 -7326 21151 -7324
rect 21119 -7354 21121 -7326
rect 21121 -7354 21149 -7326
rect 21149 -7354 21151 -7326
rect 21119 -7356 21151 -7354
rect 21119 -7486 21151 -7484
rect 21119 -7514 21121 -7486
rect 21121 -7514 21149 -7486
rect 21149 -7514 21151 -7486
rect 21119 -7516 21151 -7514
rect 21119 -7646 21151 -7644
rect 21119 -7674 21121 -7646
rect 21121 -7674 21149 -7646
rect 21149 -7674 21151 -7646
rect 21119 -7676 21151 -7674
rect 21119 -7806 21151 -7804
rect 21119 -7834 21121 -7806
rect 21121 -7834 21149 -7806
rect 21149 -7834 21151 -7806
rect 21119 -7836 21151 -7834
rect 21119 -7966 21151 -7964
rect 21119 -7994 21121 -7966
rect 21121 -7994 21149 -7966
rect 21149 -7994 21151 -7966
rect 21119 -7996 21151 -7994
rect 21119 -8126 21151 -8124
rect 21119 -8154 21121 -8126
rect 21121 -8154 21149 -8126
rect 21149 -8154 21151 -8126
rect 21119 -8156 21151 -8154
rect 21119 -8286 21151 -8284
rect 21119 -8314 21121 -8286
rect 21121 -8314 21149 -8286
rect 21149 -8314 21151 -8286
rect 21119 -8316 21151 -8314
rect 21119 -8446 21151 -8444
rect 21119 -8474 21121 -8446
rect 21121 -8474 21149 -8446
rect 21149 -8474 21151 -8446
rect 21119 -8476 21151 -8474
rect 21119 -8606 21151 -8604
rect 21119 -8634 21121 -8606
rect 21121 -8634 21149 -8606
rect 21149 -8634 21151 -8606
rect 21119 -8636 21151 -8634
rect 21119 -8766 21151 -8764
rect 21119 -8794 21121 -8766
rect 21121 -8794 21149 -8766
rect 21149 -8794 21151 -8766
rect 21119 -8796 21151 -8794
rect 21119 -8926 21151 -8924
rect 21119 -8954 21121 -8926
rect 21121 -8954 21149 -8926
rect 21149 -8954 21151 -8926
rect 21119 -8956 21151 -8954
rect 21119 -9086 21151 -9084
rect 21119 -9114 21121 -9086
rect 21121 -9114 21149 -9086
rect 21149 -9114 21151 -9086
rect 21119 -9116 21151 -9114
rect 24852 -5886 24884 -5884
rect 24852 -5914 24854 -5886
rect 24854 -5914 24882 -5886
rect 24882 -5914 24884 -5886
rect 24852 -5916 24884 -5914
rect 24852 -6046 24884 -6044
rect 24852 -6074 24854 -6046
rect 24854 -6074 24882 -6046
rect 24882 -6074 24884 -6046
rect 24852 -6076 24884 -6074
rect 24852 -6206 24884 -6204
rect 24852 -6234 24854 -6206
rect 24854 -6234 24882 -6206
rect 24882 -6234 24884 -6206
rect 24852 -6236 24884 -6234
rect 24852 -6366 24884 -6364
rect 24852 -6394 24854 -6366
rect 24854 -6394 24882 -6366
rect 24882 -6394 24884 -6366
rect 24852 -6396 24884 -6394
rect 24852 -6526 24884 -6524
rect 24852 -6554 24854 -6526
rect 24854 -6554 24882 -6526
rect 24882 -6554 24884 -6526
rect 24852 -6556 24884 -6554
rect 24852 -6686 24884 -6684
rect 24852 -6714 24854 -6686
rect 24854 -6714 24882 -6686
rect 24882 -6714 24884 -6686
rect 24852 -6716 24884 -6714
rect 24852 -6846 24884 -6844
rect 24852 -6874 24854 -6846
rect 24854 -6874 24882 -6846
rect 24882 -6874 24884 -6846
rect 24852 -6876 24884 -6874
rect 24852 -7006 24884 -7004
rect 24852 -7034 24854 -7006
rect 24854 -7034 24882 -7006
rect 24882 -7034 24884 -7006
rect 24852 -7036 24884 -7034
rect 24852 -7166 24884 -7164
rect 24852 -7194 24854 -7166
rect 24854 -7194 24882 -7166
rect 24882 -7194 24884 -7166
rect 24852 -7196 24884 -7194
rect 24852 -7326 24884 -7324
rect 24852 -7354 24854 -7326
rect 24854 -7354 24882 -7326
rect 24882 -7354 24884 -7326
rect 24852 -7356 24884 -7354
rect 24852 -7486 24884 -7484
rect 24852 -7514 24854 -7486
rect 24854 -7514 24882 -7486
rect 24882 -7514 24884 -7486
rect 24852 -7516 24884 -7514
rect 24852 -7646 24884 -7644
rect 24852 -7674 24854 -7646
rect 24854 -7674 24882 -7646
rect 24882 -7674 24884 -7646
rect 24852 -7676 24884 -7674
rect 24852 -7806 24884 -7804
rect 24852 -7834 24854 -7806
rect 24854 -7834 24882 -7806
rect 24882 -7834 24884 -7806
rect 24852 -7836 24884 -7834
rect 24852 -7966 24884 -7964
rect 24852 -7994 24854 -7966
rect 24854 -7994 24882 -7966
rect 24882 -7994 24884 -7966
rect 24852 -7996 24884 -7994
rect 24852 -8126 24884 -8124
rect 24852 -8154 24854 -8126
rect 24854 -8154 24882 -8126
rect 24882 -8154 24884 -8126
rect 24852 -8156 24884 -8154
rect 24852 -8286 24884 -8284
rect 24852 -8314 24854 -8286
rect 24854 -8314 24882 -8286
rect 24882 -8314 24884 -8286
rect 24852 -8316 24884 -8314
rect 24852 -8446 24884 -8444
rect 24852 -8474 24854 -8446
rect 24854 -8474 24882 -8446
rect 24882 -8474 24884 -8446
rect 24852 -8476 24884 -8474
rect 24852 -8606 24884 -8604
rect 24852 -8634 24854 -8606
rect 24854 -8634 24882 -8606
rect 24882 -8634 24884 -8606
rect 24852 -8636 24884 -8634
rect 24852 -8766 24884 -8764
rect 24852 -8794 24854 -8766
rect 24854 -8794 24882 -8766
rect 24882 -8794 24884 -8766
rect 24852 -8796 24884 -8794
rect 24852 -8926 24884 -8924
rect 24852 -8954 24854 -8926
rect 24854 -8954 24882 -8926
rect 24882 -8954 24884 -8926
rect 24852 -8956 24884 -8954
rect 24852 -9086 24884 -9084
rect 24852 -9114 24854 -9086
rect 24854 -9114 24882 -9086
rect 24882 -9114 24884 -9086
rect 24852 -9116 24884 -9114
rect 21119 -9246 21151 -9244
rect 21119 -9274 21121 -9246
rect 21121 -9274 21149 -9246
rect 21149 -9274 21151 -9246
rect 21119 -9276 21151 -9274
rect 24852 -9246 24884 -9244
rect 24852 -9274 24854 -9246
rect 24854 -9274 24882 -9246
rect 24882 -9274 24884 -9246
rect 24852 -9276 24884 -9274
rect 21304 -9351 21336 -9349
rect 21304 -9379 21306 -9351
rect 21306 -9379 21334 -9351
rect 21334 -9379 21336 -9351
rect 21304 -9381 21336 -9379
rect 21464 -9351 21496 -9349
rect 21464 -9379 21466 -9351
rect 21466 -9379 21494 -9351
rect 21494 -9379 21496 -9351
rect 21464 -9381 21496 -9379
rect 21624 -9351 21656 -9349
rect 21624 -9379 21626 -9351
rect 21626 -9379 21654 -9351
rect 21654 -9379 21656 -9351
rect 21624 -9381 21656 -9379
rect 21784 -9351 21816 -9349
rect 21784 -9379 21786 -9351
rect 21786 -9379 21814 -9351
rect 21814 -9379 21816 -9351
rect 21784 -9381 21816 -9379
rect 21944 -9351 21976 -9349
rect 21944 -9379 21946 -9351
rect 21946 -9379 21974 -9351
rect 21974 -9379 21976 -9351
rect 21944 -9381 21976 -9379
rect 22104 -9351 22136 -9349
rect 22104 -9379 22106 -9351
rect 22106 -9379 22134 -9351
rect 22134 -9379 22136 -9351
rect 22104 -9381 22136 -9379
rect 22264 -9351 22296 -9349
rect 22264 -9379 22266 -9351
rect 22266 -9379 22294 -9351
rect 22294 -9379 22296 -9351
rect 22264 -9381 22296 -9379
rect 22424 -9351 22456 -9349
rect 22424 -9379 22426 -9351
rect 22426 -9379 22454 -9351
rect 22454 -9379 22456 -9351
rect 22424 -9381 22456 -9379
rect 22584 -9351 22616 -9349
rect 22584 -9379 22586 -9351
rect 22586 -9379 22614 -9351
rect 22614 -9379 22616 -9351
rect 22584 -9381 22616 -9379
rect 22744 -9351 22776 -9349
rect 22744 -9379 22746 -9351
rect 22746 -9379 22774 -9351
rect 22774 -9379 22776 -9351
rect 22744 -9381 22776 -9379
rect 22904 -9351 22936 -9349
rect 22904 -9379 22906 -9351
rect 22906 -9379 22934 -9351
rect 22934 -9379 22936 -9351
rect 22904 -9381 22936 -9379
rect 23064 -9351 23096 -9349
rect 23064 -9379 23066 -9351
rect 23066 -9379 23094 -9351
rect 23094 -9379 23096 -9351
rect 23064 -9381 23096 -9379
rect 23224 -9351 23256 -9349
rect 23224 -9379 23226 -9351
rect 23226 -9379 23254 -9351
rect 23254 -9379 23256 -9351
rect 23224 -9381 23256 -9379
rect 23384 -9351 23416 -9349
rect 23384 -9379 23386 -9351
rect 23386 -9379 23414 -9351
rect 23414 -9379 23416 -9351
rect 23384 -9381 23416 -9379
rect 23544 -9351 23576 -9349
rect 23544 -9379 23546 -9351
rect 23546 -9379 23574 -9351
rect 23574 -9379 23576 -9351
rect 23544 -9381 23576 -9379
rect 23704 -9351 23736 -9349
rect 23704 -9379 23706 -9351
rect 23706 -9379 23734 -9351
rect 23734 -9379 23736 -9351
rect 23704 -9381 23736 -9379
rect 23864 -9351 23896 -9349
rect 23864 -9379 23866 -9351
rect 23866 -9379 23894 -9351
rect 23894 -9379 23896 -9351
rect 23864 -9381 23896 -9379
rect 24024 -9351 24056 -9349
rect 24024 -9379 24026 -9351
rect 24026 -9379 24054 -9351
rect 24054 -9379 24056 -9351
rect 24024 -9381 24056 -9379
rect 24184 -9351 24216 -9349
rect 24184 -9379 24186 -9351
rect 24186 -9379 24214 -9351
rect 24214 -9379 24216 -9351
rect 24184 -9381 24216 -9379
rect 24344 -9351 24376 -9349
rect 24344 -9379 24346 -9351
rect 24346 -9379 24374 -9351
rect 24374 -9379 24376 -9351
rect 24344 -9381 24376 -9379
rect 24504 -9351 24536 -9349
rect 24504 -9379 24506 -9351
rect 24506 -9379 24534 -9351
rect 24534 -9379 24536 -9351
rect 24504 -9381 24536 -9379
rect 24664 -9351 24696 -9349
rect 24664 -9379 24666 -9351
rect 24666 -9379 24694 -9351
rect 24694 -9379 24696 -9351
rect 24664 -9381 24696 -9379
rect 9304 -11623 9336 -11621
rect 9304 -11651 9306 -11623
rect 9306 -11651 9334 -11623
rect 9334 -11651 9336 -11623
rect 9304 -11653 9336 -11651
rect 9464 -11623 9496 -11621
rect 9464 -11651 9466 -11623
rect 9466 -11651 9494 -11623
rect 9494 -11651 9496 -11623
rect 9464 -11653 9496 -11651
rect 9624 -11623 9656 -11621
rect 9624 -11651 9626 -11623
rect 9626 -11651 9654 -11623
rect 9654 -11651 9656 -11623
rect 9624 -11653 9656 -11651
rect 9784 -11623 9816 -11621
rect 9784 -11651 9786 -11623
rect 9786 -11651 9814 -11623
rect 9814 -11651 9816 -11623
rect 9784 -11653 9816 -11651
rect 9944 -11623 9976 -11621
rect 9944 -11651 9946 -11623
rect 9946 -11651 9974 -11623
rect 9974 -11651 9976 -11623
rect 9944 -11653 9976 -11651
rect 10104 -11623 10136 -11621
rect 10104 -11651 10106 -11623
rect 10106 -11651 10134 -11623
rect 10134 -11651 10136 -11623
rect 10104 -11653 10136 -11651
rect 10264 -11623 10296 -11621
rect 10264 -11651 10266 -11623
rect 10266 -11651 10294 -11623
rect 10294 -11651 10296 -11623
rect 10264 -11653 10296 -11651
rect 10424 -11623 10456 -11621
rect 10424 -11651 10426 -11623
rect 10426 -11651 10454 -11623
rect 10454 -11651 10456 -11623
rect 10424 -11653 10456 -11651
rect 10584 -11623 10616 -11621
rect 10584 -11651 10586 -11623
rect 10586 -11651 10614 -11623
rect 10614 -11651 10616 -11623
rect 10584 -11653 10616 -11651
rect 10744 -11623 10776 -11621
rect 10744 -11651 10746 -11623
rect 10746 -11651 10774 -11623
rect 10774 -11651 10776 -11623
rect 10744 -11653 10776 -11651
rect 10904 -11623 10936 -11621
rect 10904 -11651 10906 -11623
rect 10906 -11651 10934 -11623
rect 10934 -11651 10936 -11623
rect 10904 -11653 10936 -11651
rect 11064 -11623 11096 -11621
rect 11064 -11651 11066 -11623
rect 11066 -11651 11094 -11623
rect 11094 -11651 11096 -11623
rect 11064 -11653 11096 -11651
rect 11224 -11623 11256 -11621
rect 11224 -11651 11226 -11623
rect 11226 -11651 11254 -11623
rect 11254 -11651 11256 -11623
rect 11224 -11653 11256 -11651
rect 11384 -11623 11416 -11621
rect 11384 -11651 11386 -11623
rect 11386 -11651 11414 -11623
rect 11414 -11651 11416 -11623
rect 11384 -11653 11416 -11651
rect 11544 -11623 11576 -11621
rect 11544 -11651 11546 -11623
rect 11546 -11651 11574 -11623
rect 11574 -11651 11576 -11623
rect 11544 -11653 11576 -11651
rect 11704 -11623 11736 -11621
rect 11704 -11651 11706 -11623
rect 11706 -11651 11734 -11623
rect 11734 -11651 11736 -11623
rect 11704 -11653 11736 -11651
rect 11864 -11623 11896 -11621
rect 11864 -11651 11866 -11623
rect 11866 -11651 11894 -11623
rect 11894 -11651 11896 -11623
rect 11864 -11653 11896 -11651
rect 12024 -11623 12056 -11621
rect 12024 -11651 12026 -11623
rect 12026 -11651 12054 -11623
rect 12054 -11651 12056 -11623
rect 12024 -11653 12056 -11651
rect 12184 -11623 12216 -11621
rect 12184 -11651 12186 -11623
rect 12186 -11651 12214 -11623
rect 12214 -11651 12216 -11623
rect 12184 -11653 12216 -11651
rect 12344 -11623 12376 -11621
rect 12344 -11651 12346 -11623
rect 12346 -11651 12374 -11623
rect 12374 -11651 12376 -11623
rect 12344 -11653 12376 -11651
rect 12504 -11623 12536 -11621
rect 12504 -11651 12506 -11623
rect 12506 -11651 12534 -11623
rect 12534 -11651 12536 -11623
rect 12504 -11653 12536 -11651
rect 12664 -11623 12696 -11621
rect 12664 -11651 12666 -11623
rect 12666 -11651 12694 -11623
rect 12694 -11651 12696 -11623
rect 12664 -11653 12696 -11651
rect 9119 -11726 9151 -11724
rect 9119 -11754 9121 -11726
rect 9121 -11754 9149 -11726
rect 9149 -11754 9151 -11726
rect 9119 -11756 9151 -11754
rect 12852 -11726 12884 -11724
rect 12852 -11754 12854 -11726
rect 12854 -11754 12882 -11726
rect 12882 -11754 12884 -11726
rect 12852 -11756 12884 -11754
rect 9119 -11886 9151 -11884
rect 9119 -11914 9121 -11886
rect 9121 -11914 9149 -11886
rect 9149 -11914 9151 -11886
rect 9119 -11916 9151 -11914
rect 9119 -12046 9151 -12044
rect 9119 -12074 9121 -12046
rect 9121 -12074 9149 -12046
rect 9149 -12074 9151 -12046
rect 9119 -12076 9151 -12074
rect 9119 -12206 9151 -12204
rect 9119 -12234 9121 -12206
rect 9121 -12234 9149 -12206
rect 9149 -12234 9151 -12206
rect 9119 -12236 9151 -12234
rect 9119 -12366 9151 -12364
rect 9119 -12394 9121 -12366
rect 9121 -12394 9149 -12366
rect 9149 -12394 9151 -12366
rect 9119 -12396 9151 -12394
rect 9119 -12526 9151 -12524
rect 9119 -12554 9121 -12526
rect 9121 -12554 9149 -12526
rect 9149 -12554 9151 -12526
rect 9119 -12556 9151 -12554
rect 9119 -12686 9151 -12684
rect 9119 -12714 9121 -12686
rect 9121 -12714 9149 -12686
rect 9149 -12714 9151 -12686
rect 9119 -12716 9151 -12714
rect 9119 -12846 9151 -12844
rect 9119 -12874 9121 -12846
rect 9121 -12874 9149 -12846
rect 9149 -12874 9151 -12846
rect 9119 -12876 9151 -12874
rect 6852 -13006 6884 -13004
rect 6852 -13034 6854 -13006
rect 6854 -13034 6882 -13006
rect 6882 -13034 6884 -13006
rect 6852 -13036 6884 -13034
rect 6852 -13166 6884 -13164
rect 6852 -13194 6854 -13166
rect 6854 -13194 6882 -13166
rect 6882 -13194 6884 -13166
rect 6852 -13196 6884 -13194
rect 6852 -13326 6884 -13324
rect 6852 -13354 6854 -13326
rect 6854 -13354 6882 -13326
rect 6882 -13354 6884 -13326
rect 6852 -13356 6884 -13354
rect 6852 -13486 6884 -13484
rect 6852 -13514 6854 -13486
rect 6854 -13514 6882 -13486
rect 6882 -13514 6884 -13486
rect 6852 -13516 6884 -13514
rect 6852 -13646 6884 -13644
rect 6852 -13674 6854 -13646
rect 6854 -13674 6882 -13646
rect 6882 -13674 6884 -13646
rect 6852 -13676 6884 -13674
rect 6852 -13806 6884 -13804
rect 6852 -13834 6854 -13806
rect 6854 -13834 6882 -13806
rect 6882 -13834 6884 -13806
rect 6852 -13836 6884 -13834
rect 6852 -13966 6884 -13964
rect 6852 -13994 6854 -13966
rect 6854 -13994 6882 -13966
rect 6882 -13994 6884 -13966
rect 6852 -13996 6884 -13994
rect 6852 -14126 6884 -14124
rect 6852 -14154 6854 -14126
rect 6854 -14154 6882 -14126
rect 6882 -14154 6884 -14126
rect 6852 -14156 6884 -14154
rect 6852 -14286 6884 -14284
rect 6852 -14314 6854 -14286
rect 6854 -14314 6882 -14286
rect 6882 -14314 6884 -14286
rect 6852 -14316 6884 -14314
rect 6852 -14446 6884 -14444
rect 6852 -14474 6854 -14446
rect 6854 -14474 6882 -14446
rect 6882 -14474 6884 -14446
rect 6852 -14476 6884 -14474
rect 6852 -14606 6884 -14604
rect 6852 -14634 6854 -14606
rect 6854 -14634 6882 -14606
rect 6882 -14634 6884 -14606
rect 6852 -14636 6884 -14634
rect 6852 -14766 6884 -14764
rect 6852 -14794 6854 -14766
rect 6854 -14794 6882 -14766
rect 6882 -14794 6884 -14766
rect 6852 -14796 6884 -14794
rect 6852 -14926 6884 -14924
rect 6852 -14954 6854 -14926
rect 6854 -14954 6882 -14926
rect 6882 -14954 6884 -14926
rect 6852 -14956 6884 -14954
rect 6852 -15086 6884 -15084
rect 6852 -15114 6854 -15086
rect 6854 -15114 6882 -15086
rect 6882 -15114 6884 -15086
rect 6852 -15116 6884 -15114
rect 3119 -15246 3151 -15244
rect 3119 -15274 3121 -15246
rect 3121 -15274 3149 -15246
rect 3149 -15274 3151 -15246
rect 3119 -15276 3151 -15274
rect 6852 -15246 6884 -15244
rect 6852 -15274 6854 -15246
rect 6854 -15274 6882 -15246
rect 6882 -15274 6884 -15246
rect 6852 -15276 6884 -15274
rect 3304 -15351 3336 -15349
rect 3304 -15379 3306 -15351
rect 3306 -15379 3334 -15351
rect 3334 -15379 3336 -15351
rect 3304 -15381 3336 -15379
rect 3464 -15351 3496 -15349
rect 3464 -15379 3466 -15351
rect 3466 -15379 3494 -15351
rect 3494 -15379 3496 -15351
rect 3464 -15381 3496 -15379
rect 3624 -15351 3656 -15349
rect 3624 -15379 3626 -15351
rect 3626 -15379 3654 -15351
rect 3654 -15379 3656 -15351
rect 3624 -15381 3656 -15379
rect 3784 -15351 3816 -15349
rect 3784 -15379 3786 -15351
rect 3786 -15379 3814 -15351
rect 3814 -15379 3816 -15351
rect 3784 -15381 3816 -15379
rect 3944 -15351 3976 -15349
rect 3944 -15379 3946 -15351
rect 3946 -15379 3974 -15351
rect 3974 -15379 3976 -15351
rect 3944 -15381 3976 -15379
rect 4104 -15351 4136 -15349
rect 4104 -15379 4106 -15351
rect 4106 -15379 4134 -15351
rect 4134 -15379 4136 -15351
rect 4104 -15381 4136 -15379
rect 4264 -15351 4296 -15349
rect 4264 -15379 4266 -15351
rect 4266 -15379 4294 -15351
rect 4294 -15379 4296 -15351
rect 4264 -15381 4296 -15379
rect 4424 -15351 4456 -15349
rect 4424 -15379 4426 -15351
rect 4426 -15379 4454 -15351
rect 4454 -15379 4456 -15351
rect 4424 -15381 4456 -15379
rect 4584 -15351 4616 -15349
rect 4584 -15379 4586 -15351
rect 4586 -15379 4614 -15351
rect 4614 -15379 4616 -15351
rect 4584 -15381 4616 -15379
rect 4744 -15351 4776 -15349
rect 4744 -15379 4746 -15351
rect 4746 -15379 4774 -15351
rect 4774 -15379 4776 -15351
rect 4744 -15381 4776 -15379
rect 4904 -15351 4936 -15349
rect 4904 -15379 4906 -15351
rect 4906 -15379 4934 -15351
rect 4934 -15379 4936 -15351
rect 4904 -15381 4936 -15379
rect 5064 -15351 5096 -15349
rect 5064 -15379 5066 -15351
rect 5066 -15379 5094 -15351
rect 5094 -15379 5096 -15351
rect 5064 -15381 5096 -15379
rect 5224 -15351 5256 -15349
rect 5224 -15379 5226 -15351
rect 5226 -15379 5254 -15351
rect 5254 -15379 5256 -15351
rect 5224 -15381 5256 -15379
rect 5384 -15351 5416 -15349
rect 5384 -15379 5386 -15351
rect 5386 -15379 5414 -15351
rect 5414 -15379 5416 -15351
rect 5384 -15381 5416 -15379
rect 5544 -15351 5576 -15349
rect 5544 -15379 5546 -15351
rect 5546 -15379 5574 -15351
rect 5574 -15379 5576 -15351
rect 5544 -15381 5576 -15379
rect 5704 -15351 5736 -15349
rect 5704 -15379 5706 -15351
rect 5706 -15379 5734 -15351
rect 5734 -15379 5736 -15351
rect 5704 -15381 5736 -15379
rect 5864 -15351 5896 -15349
rect 5864 -15379 5866 -15351
rect 5866 -15379 5894 -15351
rect 5894 -15379 5896 -15351
rect 5864 -15381 5896 -15379
rect 6024 -15351 6056 -15349
rect 6024 -15379 6026 -15351
rect 6026 -15379 6054 -15351
rect 6054 -15379 6056 -15351
rect 6024 -15381 6056 -15379
rect 6184 -15351 6216 -15349
rect 6184 -15379 6186 -15351
rect 6186 -15379 6214 -15351
rect 6214 -15379 6216 -15351
rect 6184 -15381 6216 -15379
rect 6344 -15351 6376 -15349
rect 6344 -15379 6346 -15351
rect 6346 -15379 6374 -15351
rect 6374 -15379 6376 -15351
rect 6344 -15381 6376 -15379
rect 6504 -15351 6536 -15349
rect 6504 -15379 6506 -15351
rect 6506 -15379 6534 -15351
rect 6534 -15379 6536 -15351
rect 6504 -15381 6536 -15379
rect 6664 -15351 6696 -15349
rect 6664 -15379 6666 -15351
rect 6666 -15379 6694 -15351
rect 6694 -15379 6696 -15351
rect 6664 -15381 6696 -15379
rect 9119 -13006 9151 -13004
rect 9119 -13034 9121 -13006
rect 9121 -13034 9149 -13006
rect 9149 -13034 9151 -13006
rect 9119 -13036 9151 -13034
rect 9119 -13166 9151 -13164
rect 9119 -13194 9121 -13166
rect 9121 -13194 9149 -13166
rect 9149 -13194 9151 -13166
rect 9119 -13196 9151 -13194
rect 9119 -13326 9151 -13324
rect 9119 -13354 9121 -13326
rect 9121 -13354 9149 -13326
rect 9149 -13354 9151 -13326
rect 9119 -13356 9151 -13354
rect 9119 -13486 9151 -13484
rect 9119 -13514 9121 -13486
rect 9121 -13514 9149 -13486
rect 9149 -13514 9151 -13486
rect 9119 -13516 9151 -13514
rect 9119 -13646 9151 -13644
rect 9119 -13674 9121 -13646
rect 9121 -13674 9149 -13646
rect 9149 -13674 9151 -13646
rect 9119 -13676 9151 -13674
rect 9119 -13806 9151 -13804
rect 9119 -13834 9121 -13806
rect 9121 -13834 9149 -13806
rect 9149 -13834 9151 -13806
rect 9119 -13836 9151 -13834
rect 9119 -13966 9151 -13964
rect 9119 -13994 9121 -13966
rect 9121 -13994 9149 -13966
rect 9149 -13994 9151 -13966
rect 9119 -13996 9151 -13994
rect 9119 -14126 9151 -14124
rect 9119 -14154 9121 -14126
rect 9121 -14154 9149 -14126
rect 9149 -14154 9151 -14126
rect 9119 -14156 9151 -14154
rect 9119 -14286 9151 -14284
rect 9119 -14314 9121 -14286
rect 9121 -14314 9149 -14286
rect 9149 -14314 9151 -14286
rect 9119 -14316 9151 -14314
rect 9119 -14446 9151 -14444
rect 9119 -14474 9121 -14446
rect 9121 -14474 9149 -14446
rect 9149 -14474 9151 -14446
rect 9119 -14476 9151 -14474
rect 9119 -14606 9151 -14604
rect 9119 -14634 9121 -14606
rect 9121 -14634 9149 -14606
rect 9149 -14634 9151 -14606
rect 9119 -14636 9151 -14634
rect 9119 -14766 9151 -14764
rect 9119 -14794 9121 -14766
rect 9121 -14794 9149 -14766
rect 9149 -14794 9151 -14766
rect 9119 -14796 9151 -14794
rect 9119 -14926 9151 -14924
rect 9119 -14954 9121 -14926
rect 9121 -14954 9149 -14926
rect 9149 -14954 9151 -14926
rect 9119 -14956 9151 -14954
rect 9119 -15086 9151 -15084
rect 9119 -15114 9121 -15086
rect 9121 -15114 9149 -15086
rect 9149 -15114 9151 -15086
rect 9119 -15116 9151 -15114
rect 12852 -11886 12884 -11884
rect 12852 -11914 12854 -11886
rect 12854 -11914 12882 -11886
rect 12882 -11914 12884 -11886
rect 12852 -11916 12884 -11914
rect 12852 -12046 12884 -12044
rect 12852 -12074 12854 -12046
rect 12854 -12074 12882 -12046
rect 12882 -12074 12884 -12046
rect 12852 -12076 12884 -12074
rect 12852 -12206 12884 -12204
rect 12852 -12234 12854 -12206
rect 12854 -12234 12882 -12206
rect 12882 -12234 12884 -12206
rect 12852 -12236 12884 -12234
rect 12852 -12366 12884 -12364
rect 12852 -12394 12854 -12366
rect 12854 -12394 12882 -12366
rect 12882 -12394 12884 -12366
rect 12852 -12396 12884 -12394
rect 12852 -12526 12884 -12524
rect 12852 -12554 12854 -12526
rect 12854 -12554 12882 -12526
rect 12882 -12554 12884 -12526
rect 12852 -12556 12884 -12554
rect 12852 -12686 12884 -12684
rect 12852 -12714 12854 -12686
rect 12854 -12714 12882 -12686
rect 12882 -12714 12884 -12686
rect 12852 -12716 12884 -12714
rect 12852 -12846 12884 -12844
rect 12852 -12874 12854 -12846
rect 12854 -12874 12882 -12846
rect 12882 -12874 12884 -12846
rect 12852 -12876 12884 -12874
rect 15304 -11623 15336 -11621
rect 15304 -11651 15306 -11623
rect 15306 -11651 15334 -11623
rect 15334 -11651 15336 -11623
rect 15304 -11653 15336 -11651
rect 15464 -11623 15496 -11621
rect 15464 -11651 15466 -11623
rect 15466 -11651 15494 -11623
rect 15494 -11651 15496 -11623
rect 15464 -11653 15496 -11651
rect 15624 -11623 15656 -11621
rect 15624 -11651 15626 -11623
rect 15626 -11651 15654 -11623
rect 15654 -11651 15656 -11623
rect 15624 -11653 15656 -11651
rect 15784 -11623 15816 -11621
rect 15784 -11651 15786 -11623
rect 15786 -11651 15814 -11623
rect 15814 -11651 15816 -11623
rect 15784 -11653 15816 -11651
rect 15944 -11623 15976 -11621
rect 15944 -11651 15946 -11623
rect 15946 -11651 15974 -11623
rect 15974 -11651 15976 -11623
rect 15944 -11653 15976 -11651
rect 16104 -11623 16136 -11621
rect 16104 -11651 16106 -11623
rect 16106 -11651 16134 -11623
rect 16134 -11651 16136 -11623
rect 16104 -11653 16136 -11651
rect 16264 -11623 16296 -11621
rect 16264 -11651 16266 -11623
rect 16266 -11651 16294 -11623
rect 16294 -11651 16296 -11623
rect 16264 -11653 16296 -11651
rect 16424 -11623 16456 -11621
rect 16424 -11651 16426 -11623
rect 16426 -11651 16454 -11623
rect 16454 -11651 16456 -11623
rect 16424 -11653 16456 -11651
rect 16584 -11623 16616 -11621
rect 16584 -11651 16586 -11623
rect 16586 -11651 16614 -11623
rect 16614 -11651 16616 -11623
rect 16584 -11653 16616 -11651
rect 16744 -11623 16776 -11621
rect 16744 -11651 16746 -11623
rect 16746 -11651 16774 -11623
rect 16774 -11651 16776 -11623
rect 16744 -11653 16776 -11651
rect 16904 -11623 16936 -11621
rect 16904 -11651 16906 -11623
rect 16906 -11651 16934 -11623
rect 16934 -11651 16936 -11623
rect 16904 -11653 16936 -11651
rect 17064 -11623 17096 -11621
rect 17064 -11651 17066 -11623
rect 17066 -11651 17094 -11623
rect 17094 -11651 17096 -11623
rect 17064 -11653 17096 -11651
rect 17224 -11623 17256 -11621
rect 17224 -11651 17226 -11623
rect 17226 -11651 17254 -11623
rect 17254 -11651 17256 -11623
rect 17224 -11653 17256 -11651
rect 17384 -11623 17416 -11621
rect 17384 -11651 17386 -11623
rect 17386 -11651 17414 -11623
rect 17414 -11651 17416 -11623
rect 17384 -11653 17416 -11651
rect 17544 -11623 17576 -11621
rect 17544 -11651 17546 -11623
rect 17546 -11651 17574 -11623
rect 17574 -11651 17576 -11623
rect 17544 -11653 17576 -11651
rect 17704 -11623 17736 -11621
rect 17704 -11651 17706 -11623
rect 17706 -11651 17734 -11623
rect 17734 -11651 17736 -11623
rect 17704 -11653 17736 -11651
rect 17864 -11623 17896 -11621
rect 17864 -11651 17866 -11623
rect 17866 -11651 17894 -11623
rect 17894 -11651 17896 -11623
rect 17864 -11653 17896 -11651
rect 18024 -11623 18056 -11621
rect 18024 -11651 18026 -11623
rect 18026 -11651 18054 -11623
rect 18054 -11651 18056 -11623
rect 18024 -11653 18056 -11651
rect 18184 -11623 18216 -11621
rect 18184 -11651 18186 -11623
rect 18186 -11651 18214 -11623
rect 18214 -11651 18216 -11623
rect 18184 -11653 18216 -11651
rect 18344 -11623 18376 -11621
rect 18344 -11651 18346 -11623
rect 18346 -11651 18374 -11623
rect 18374 -11651 18376 -11623
rect 18344 -11653 18376 -11651
rect 18504 -11623 18536 -11621
rect 18504 -11651 18506 -11623
rect 18506 -11651 18534 -11623
rect 18534 -11651 18536 -11623
rect 18504 -11653 18536 -11651
rect 18664 -11623 18696 -11621
rect 18664 -11651 18666 -11623
rect 18666 -11651 18694 -11623
rect 18694 -11651 18696 -11623
rect 18664 -11653 18696 -11651
rect 15119 -11726 15151 -11724
rect 15119 -11754 15121 -11726
rect 15121 -11754 15149 -11726
rect 15149 -11754 15151 -11726
rect 15119 -11756 15151 -11754
rect 18852 -11726 18884 -11724
rect 18852 -11754 18854 -11726
rect 18854 -11754 18882 -11726
rect 18882 -11754 18884 -11726
rect 18852 -11756 18884 -11754
rect 15119 -11886 15151 -11884
rect 15119 -11914 15121 -11886
rect 15121 -11914 15149 -11886
rect 15149 -11914 15151 -11886
rect 15119 -11916 15151 -11914
rect 15119 -12046 15151 -12044
rect 15119 -12074 15121 -12046
rect 15121 -12074 15149 -12046
rect 15149 -12074 15151 -12046
rect 15119 -12076 15151 -12074
rect 15119 -12206 15151 -12204
rect 15119 -12234 15121 -12206
rect 15121 -12234 15149 -12206
rect 15149 -12234 15151 -12206
rect 15119 -12236 15151 -12234
rect 15119 -12366 15151 -12364
rect 15119 -12394 15121 -12366
rect 15121 -12394 15149 -12366
rect 15149 -12394 15151 -12366
rect 15119 -12396 15151 -12394
rect 15119 -12526 15151 -12524
rect 15119 -12554 15121 -12526
rect 15121 -12554 15149 -12526
rect 15149 -12554 15151 -12526
rect 15119 -12556 15151 -12554
rect 15119 -12686 15151 -12684
rect 15119 -12714 15121 -12686
rect 15121 -12714 15149 -12686
rect 15149 -12714 15151 -12686
rect 15119 -12716 15151 -12714
rect 15119 -12846 15151 -12844
rect 15119 -12874 15121 -12846
rect 15121 -12874 15149 -12846
rect 15149 -12874 15151 -12846
rect 15119 -12876 15151 -12874
rect 12852 -13006 12884 -13004
rect 12852 -13034 12854 -13006
rect 12854 -13034 12882 -13006
rect 12882 -13034 12884 -13006
rect 12852 -13036 12884 -13034
rect 12852 -13166 12884 -13164
rect 12852 -13194 12854 -13166
rect 12854 -13194 12882 -13166
rect 12882 -13194 12884 -13166
rect 12852 -13196 12884 -13194
rect 12852 -13326 12884 -13324
rect 12852 -13354 12854 -13326
rect 12854 -13354 12882 -13326
rect 12882 -13354 12884 -13326
rect 12852 -13356 12884 -13354
rect 12852 -13486 12884 -13484
rect 12852 -13514 12854 -13486
rect 12854 -13514 12882 -13486
rect 12882 -13514 12884 -13486
rect 12852 -13516 12884 -13514
rect 12852 -13646 12884 -13644
rect 12852 -13674 12854 -13646
rect 12854 -13674 12882 -13646
rect 12882 -13674 12884 -13646
rect 12852 -13676 12884 -13674
rect 12852 -13806 12884 -13804
rect 12852 -13834 12854 -13806
rect 12854 -13834 12882 -13806
rect 12882 -13834 12884 -13806
rect 12852 -13836 12884 -13834
rect 12852 -13966 12884 -13964
rect 12852 -13994 12854 -13966
rect 12854 -13994 12882 -13966
rect 12882 -13994 12884 -13966
rect 12852 -13996 12884 -13994
rect 12852 -14126 12884 -14124
rect 12852 -14154 12854 -14126
rect 12854 -14154 12882 -14126
rect 12882 -14154 12884 -14126
rect 12852 -14156 12884 -14154
rect 12852 -14286 12884 -14284
rect 12852 -14314 12854 -14286
rect 12854 -14314 12882 -14286
rect 12882 -14314 12884 -14286
rect 12852 -14316 12884 -14314
rect 12852 -14446 12884 -14444
rect 12852 -14474 12854 -14446
rect 12854 -14474 12882 -14446
rect 12882 -14474 12884 -14446
rect 12852 -14476 12884 -14474
rect 12852 -14606 12884 -14604
rect 12852 -14634 12854 -14606
rect 12854 -14634 12882 -14606
rect 12882 -14634 12884 -14606
rect 12852 -14636 12884 -14634
rect 12852 -14766 12884 -14764
rect 12852 -14794 12854 -14766
rect 12854 -14794 12882 -14766
rect 12882 -14794 12884 -14766
rect 12852 -14796 12884 -14794
rect 12852 -14926 12884 -14924
rect 12852 -14954 12854 -14926
rect 12854 -14954 12882 -14926
rect 12882 -14954 12884 -14926
rect 12852 -14956 12884 -14954
rect 12852 -15086 12884 -15084
rect 12852 -15114 12854 -15086
rect 12854 -15114 12882 -15086
rect 12882 -15114 12884 -15086
rect 12852 -15116 12884 -15114
rect 9119 -15246 9151 -15244
rect 9119 -15274 9121 -15246
rect 9121 -15274 9149 -15246
rect 9149 -15274 9151 -15246
rect 9119 -15276 9151 -15274
rect 12852 -15246 12884 -15244
rect 12852 -15274 12854 -15246
rect 12854 -15274 12882 -15246
rect 12882 -15274 12884 -15246
rect 12852 -15276 12884 -15274
rect 9304 -15351 9336 -15349
rect 9304 -15379 9306 -15351
rect 9306 -15379 9334 -15351
rect 9334 -15379 9336 -15351
rect 9304 -15381 9336 -15379
rect 9464 -15351 9496 -15349
rect 9464 -15379 9466 -15351
rect 9466 -15379 9494 -15351
rect 9494 -15379 9496 -15351
rect 9464 -15381 9496 -15379
rect 9624 -15351 9656 -15349
rect 9624 -15379 9626 -15351
rect 9626 -15379 9654 -15351
rect 9654 -15379 9656 -15351
rect 9624 -15381 9656 -15379
rect 9784 -15351 9816 -15349
rect 9784 -15379 9786 -15351
rect 9786 -15379 9814 -15351
rect 9814 -15379 9816 -15351
rect 9784 -15381 9816 -15379
rect 9944 -15351 9976 -15349
rect 9944 -15379 9946 -15351
rect 9946 -15379 9974 -15351
rect 9974 -15379 9976 -15351
rect 9944 -15381 9976 -15379
rect 10104 -15351 10136 -15349
rect 10104 -15379 10106 -15351
rect 10106 -15379 10134 -15351
rect 10134 -15379 10136 -15351
rect 10104 -15381 10136 -15379
rect 10264 -15351 10296 -15349
rect 10264 -15379 10266 -15351
rect 10266 -15379 10294 -15351
rect 10294 -15379 10296 -15351
rect 10264 -15381 10296 -15379
rect 10424 -15351 10456 -15349
rect 10424 -15379 10426 -15351
rect 10426 -15379 10454 -15351
rect 10454 -15379 10456 -15351
rect 10424 -15381 10456 -15379
rect 10584 -15351 10616 -15349
rect 10584 -15379 10586 -15351
rect 10586 -15379 10614 -15351
rect 10614 -15379 10616 -15351
rect 10584 -15381 10616 -15379
rect 10744 -15351 10776 -15349
rect 10744 -15379 10746 -15351
rect 10746 -15379 10774 -15351
rect 10774 -15379 10776 -15351
rect 10744 -15381 10776 -15379
rect 10904 -15351 10936 -15349
rect 10904 -15379 10906 -15351
rect 10906 -15379 10934 -15351
rect 10934 -15379 10936 -15351
rect 10904 -15381 10936 -15379
rect 11064 -15351 11096 -15349
rect 11064 -15379 11066 -15351
rect 11066 -15379 11094 -15351
rect 11094 -15379 11096 -15351
rect 11064 -15381 11096 -15379
rect 11224 -15351 11256 -15349
rect 11224 -15379 11226 -15351
rect 11226 -15379 11254 -15351
rect 11254 -15379 11256 -15351
rect 11224 -15381 11256 -15379
rect 11384 -15351 11416 -15349
rect 11384 -15379 11386 -15351
rect 11386 -15379 11414 -15351
rect 11414 -15379 11416 -15351
rect 11384 -15381 11416 -15379
rect 11544 -15351 11576 -15349
rect 11544 -15379 11546 -15351
rect 11546 -15379 11574 -15351
rect 11574 -15379 11576 -15351
rect 11544 -15381 11576 -15379
rect 11704 -15351 11736 -15349
rect 11704 -15379 11706 -15351
rect 11706 -15379 11734 -15351
rect 11734 -15379 11736 -15351
rect 11704 -15381 11736 -15379
rect 11864 -15351 11896 -15349
rect 11864 -15379 11866 -15351
rect 11866 -15379 11894 -15351
rect 11894 -15379 11896 -15351
rect 11864 -15381 11896 -15379
rect 12024 -15351 12056 -15349
rect 12024 -15379 12026 -15351
rect 12026 -15379 12054 -15351
rect 12054 -15379 12056 -15351
rect 12024 -15381 12056 -15379
rect 12184 -15351 12216 -15349
rect 12184 -15379 12186 -15351
rect 12186 -15379 12214 -15351
rect 12214 -15379 12216 -15351
rect 12184 -15381 12216 -15379
rect 12344 -15351 12376 -15349
rect 12344 -15379 12346 -15351
rect 12346 -15379 12374 -15351
rect 12374 -15379 12376 -15351
rect 12344 -15381 12376 -15379
rect 12504 -15351 12536 -15349
rect 12504 -15379 12506 -15351
rect 12506 -15379 12534 -15351
rect 12534 -15379 12536 -15351
rect 12504 -15381 12536 -15379
rect 12664 -15351 12696 -15349
rect 12664 -15379 12666 -15351
rect 12666 -15379 12694 -15351
rect 12694 -15379 12696 -15351
rect 12664 -15381 12696 -15379
rect 15119 -13006 15151 -13004
rect 15119 -13034 15121 -13006
rect 15121 -13034 15149 -13006
rect 15149 -13034 15151 -13006
rect 15119 -13036 15151 -13034
rect 15119 -13166 15151 -13164
rect 15119 -13194 15121 -13166
rect 15121 -13194 15149 -13166
rect 15149 -13194 15151 -13166
rect 15119 -13196 15151 -13194
rect 15119 -13326 15151 -13324
rect 15119 -13354 15121 -13326
rect 15121 -13354 15149 -13326
rect 15149 -13354 15151 -13326
rect 15119 -13356 15151 -13354
rect 15119 -13486 15151 -13484
rect 15119 -13514 15121 -13486
rect 15121 -13514 15149 -13486
rect 15149 -13514 15151 -13486
rect 15119 -13516 15151 -13514
rect 15119 -13646 15151 -13644
rect 15119 -13674 15121 -13646
rect 15121 -13674 15149 -13646
rect 15149 -13674 15151 -13646
rect 15119 -13676 15151 -13674
rect 15119 -13806 15151 -13804
rect 15119 -13834 15121 -13806
rect 15121 -13834 15149 -13806
rect 15149 -13834 15151 -13806
rect 15119 -13836 15151 -13834
rect 15119 -13966 15151 -13964
rect 15119 -13994 15121 -13966
rect 15121 -13994 15149 -13966
rect 15149 -13994 15151 -13966
rect 15119 -13996 15151 -13994
rect 15119 -14126 15151 -14124
rect 15119 -14154 15121 -14126
rect 15121 -14154 15149 -14126
rect 15149 -14154 15151 -14126
rect 15119 -14156 15151 -14154
rect 15119 -14286 15151 -14284
rect 15119 -14314 15121 -14286
rect 15121 -14314 15149 -14286
rect 15149 -14314 15151 -14286
rect 15119 -14316 15151 -14314
rect 15119 -14446 15151 -14444
rect 15119 -14474 15121 -14446
rect 15121 -14474 15149 -14446
rect 15149 -14474 15151 -14446
rect 15119 -14476 15151 -14474
rect 15119 -14606 15151 -14604
rect 15119 -14634 15121 -14606
rect 15121 -14634 15149 -14606
rect 15149 -14634 15151 -14606
rect 15119 -14636 15151 -14634
rect 15119 -14766 15151 -14764
rect 15119 -14794 15121 -14766
rect 15121 -14794 15149 -14766
rect 15149 -14794 15151 -14766
rect 15119 -14796 15151 -14794
rect 15119 -14926 15151 -14924
rect 15119 -14954 15121 -14926
rect 15121 -14954 15149 -14926
rect 15149 -14954 15151 -14926
rect 15119 -14956 15151 -14954
rect 15119 -15086 15151 -15084
rect 15119 -15114 15121 -15086
rect 15121 -15114 15149 -15086
rect 15149 -15114 15151 -15086
rect 15119 -15116 15151 -15114
rect 18852 -11886 18884 -11884
rect 18852 -11914 18854 -11886
rect 18854 -11914 18882 -11886
rect 18882 -11914 18884 -11886
rect 18852 -11916 18884 -11914
rect 18852 -12046 18884 -12044
rect 18852 -12074 18854 -12046
rect 18854 -12074 18882 -12046
rect 18882 -12074 18884 -12046
rect 18852 -12076 18884 -12074
rect 18852 -12206 18884 -12204
rect 18852 -12234 18854 -12206
rect 18854 -12234 18882 -12206
rect 18882 -12234 18884 -12206
rect 18852 -12236 18884 -12234
rect 18852 -12366 18884 -12364
rect 18852 -12394 18854 -12366
rect 18854 -12394 18882 -12366
rect 18882 -12394 18884 -12366
rect 18852 -12396 18884 -12394
rect 18852 -12526 18884 -12524
rect 18852 -12554 18854 -12526
rect 18854 -12554 18882 -12526
rect 18882 -12554 18884 -12526
rect 18852 -12556 18884 -12554
rect 18852 -12686 18884 -12684
rect 18852 -12714 18854 -12686
rect 18854 -12714 18882 -12686
rect 18882 -12714 18884 -12686
rect 18852 -12716 18884 -12714
rect 18852 -12846 18884 -12844
rect 18852 -12874 18854 -12846
rect 18854 -12874 18882 -12846
rect 18882 -12874 18884 -12846
rect 18852 -12876 18884 -12874
rect 18852 -13006 18884 -13004
rect 18852 -13034 18854 -13006
rect 18854 -13034 18882 -13006
rect 18882 -13034 18884 -13006
rect 18852 -13036 18884 -13034
rect 18852 -13166 18884 -13164
rect 18852 -13194 18854 -13166
rect 18854 -13194 18882 -13166
rect 18882 -13194 18884 -13166
rect 18852 -13196 18884 -13194
rect 18852 -13326 18884 -13324
rect 18852 -13354 18854 -13326
rect 18854 -13354 18882 -13326
rect 18882 -13354 18884 -13326
rect 18852 -13356 18884 -13354
rect 18852 -13486 18884 -13484
rect 18852 -13514 18854 -13486
rect 18854 -13514 18882 -13486
rect 18882 -13514 18884 -13486
rect 18852 -13516 18884 -13514
rect 18852 -13646 18884 -13644
rect 18852 -13674 18854 -13646
rect 18854 -13674 18882 -13646
rect 18882 -13674 18884 -13646
rect 18852 -13676 18884 -13674
rect 18852 -13806 18884 -13804
rect 18852 -13834 18854 -13806
rect 18854 -13834 18882 -13806
rect 18882 -13834 18884 -13806
rect 18852 -13836 18884 -13834
rect 18852 -13966 18884 -13964
rect 18852 -13994 18854 -13966
rect 18854 -13994 18882 -13966
rect 18882 -13994 18884 -13966
rect 18852 -13996 18884 -13994
rect 18852 -14126 18884 -14124
rect 18852 -14154 18854 -14126
rect 18854 -14154 18882 -14126
rect 18882 -14154 18884 -14126
rect 18852 -14156 18884 -14154
rect 18852 -14286 18884 -14284
rect 18852 -14314 18854 -14286
rect 18854 -14314 18882 -14286
rect 18882 -14314 18884 -14286
rect 18852 -14316 18884 -14314
rect 18852 -14446 18884 -14444
rect 18852 -14474 18854 -14446
rect 18854 -14474 18882 -14446
rect 18882 -14474 18884 -14446
rect 18852 -14476 18884 -14474
rect 18852 -14606 18884 -14604
rect 18852 -14634 18854 -14606
rect 18854 -14634 18882 -14606
rect 18882 -14634 18884 -14606
rect 18852 -14636 18884 -14634
rect 18852 -14766 18884 -14764
rect 18852 -14794 18854 -14766
rect 18854 -14794 18882 -14766
rect 18882 -14794 18884 -14766
rect 18852 -14796 18884 -14794
rect 18852 -14926 18884 -14924
rect 18852 -14954 18854 -14926
rect 18854 -14954 18882 -14926
rect 18882 -14954 18884 -14926
rect 18852 -14956 18884 -14954
rect 18852 -15086 18884 -15084
rect 18852 -15114 18854 -15086
rect 18854 -15114 18882 -15086
rect 18882 -15114 18884 -15086
rect 18852 -15116 18884 -15114
rect 15119 -15246 15151 -15244
rect 15119 -15274 15121 -15246
rect 15121 -15274 15149 -15246
rect 15149 -15274 15151 -15246
rect 15119 -15276 15151 -15274
rect 18852 -15246 18884 -15244
rect 18852 -15274 18854 -15246
rect 18854 -15274 18882 -15246
rect 18882 -15274 18884 -15246
rect 18852 -15276 18884 -15274
rect 15304 -15351 15336 -15349
rect 15304 -15379 15306 -15351
rect 15306 -15379 15334 -15351
rect 15334 -15379 15336 -15351
rect 15304 -15381 15336 -15379
rect 15464 -15351 15496 -15349
rect 15464 -15379 15466 -15351
rect 15466 -15379 15494 -15351
rect 15494 -15379 15496 -15351
rect 15464 -15381 15496 -15379
rect 15624 -15351 15656 -15349
rect 15624 -15379 15626 -15351
rect 15626 -15379 15654 -15351
rect 15654 -15379 15656 -15351
rect 15624 -15381 15656 -15379
rect 15784 -15351 15816 -15349
rect 15784 -15379 15786 -15351
rect 15786 -15379 15814 -15351
rect 15814 -15379 15816 -15351
rect 15784 -15381 15816 -15379
rect 15944 -15351 15976 -15349
rect 15944 -15379 15946 -15351
rect 15946 -15379 15974 -15351
rect 15974 -15379 15976 -15351
rect 15944 -15381 15976 -15379
rect 16104 -15351 16136 -15349
rect 16104 -15379 16106 -15351
rect 16106 -15379 16134 -15351
rect 16134 -15379 16136 -15351
rect 16104 -15381 16136 -15379
rect 16264 -15351 16296 -15349
rect 16264 -15379 16266 -15351
rect 16266 -15379 16294 -15351
rect 16294 -15379 16296 -15351
rect 16264 -15381 16296 -15379
rect 16424 -15351 16456 -15349
rect 16424 -15379 16426 -15351
rect 16426 -15379 16454 -15351
rect 16454 -15379 16456 -15351
rect 16424 -15381 16456 -15379
rect 16584 -15351 16616 -15349
rect 16584 -15379 16586 -15351
rect 16586 -15379 16614 -15351
rect 16614 -15379 16616 -15351
rect 16584 -15381 16616 -15379
rect 16744 -15351 16776 -15349
rect 16744 -15379 16746 -15351
rect 16746 -15379 16774 -15351
rect 16774 -15379 16776 -15351
rect 16744 -15381 16776 -15379
rect 16904 -15351 16936 -15349
rect 16904 -15379 16906 -15351
rect 16906 -15379 16934 -15351
rect 16934 -15379 16936 -15351
rect 16904 -15381 16936 -15379
rect 17064 -15351 17096 -15349
rect 17064 -15379 17066 -15351
rect 17066 -15379 17094 -15351
rect 17094 -15379 17096 -15351
rect 17064 -15381 17096 -15379
rect 17224 -15351 17256 -15349
rect 17224 -15379 17226 -15351
rect 17226 -15379 17254 -15351
rect 17254 -15379 17256 -15351
rect 17224 -15381 17256 -15379
rect 17384 -15351 17416 -15349
rect 17384 -15379 17386 -15351
rect 17386 -15379 17414 -15351
rect 17414 -15379 17416 -15351
rect 17384 -15381 17416 -15379
rect 17544 -15351 17576 -15349
rect 17544 -15379 17546 -15351
rect 17546 -15379 17574 -15351
rect 17574 -15379 17576 -15351
rect 17544 -15381 17576 -15379
rect 17704 -15351 17736 -15349
rect 17704 -15379 17706 -15351
rect 17706 -15379 17734 -15351
rect 17734 -15379 17736 -15351
rect 17704 -15381 17736 -15379
rect 17864 -15351 17896 -15349
rect 17864 -15379 17866 -15351
rect 17866 -15379 17894 -15351
rect 17894 -15379 17896 -15351
rect 17864 -15381 17896 -15379
rect 18024 -15351 18056 -15349
rect 18024 -15379 18026 -15351
rect 18026 -15379 18054 -15351
rect 18054 -15379 18056 -15351
rect 18024 -15381 18056 -15379
rect 18184 -15351 18216 -15349
rect 18184 -15379 18186 -15351
rect 18186 -15379 18214 -15351
rect 18214 -15379 18216 -15351
rect 18184 -15381 18216 -15379
rect 18344 -15351 18376 -15349
rect 18344 -15379 18346 -15351
rect 18346 -15379 18374 -15351
rect 18374 -15379 18376 -15351
rect 18344 -15381 18376 -15379
rect 18504 -15351 18536 -15349
rect 18504 -15379 18506 -15351
rect 18506 -15379 18534 -15351
rect 18534 -15379 18536 -15351
rect 18504 -15381 18536 -15379
rect 18664 -15351 18696 -15349
rect 18664 -15379 18666 -15351
rect 18666 -15379 18694 -15351
rect 18694 -15379 18696 -15351
rect 18664 -15381 18696 -15379
rect 21304 -11623 21336 -11621
rect 21304 -11651 21306 -11623
rect 21306 -11651 21334 -11623
rect 21334 -11651 21336 -11623
rect 21304 -11653 21336 -11651
rect 21464 -11623 21496 -11621
rect 21464 -11651 21466 -11623
rect 21466 -11651 21494 -11623
rect 21494 -11651 21496 -11623
rect 21464 -11653 21496 -11651
rect 21624 -11623 21656 -11621
rect 21624 -11651 21626 -11623
rect 21626 -11651 21654 -11623
rect 21654 -11651 21656 -11623
rect 21624 -11653 21656 -11651
rect 21784 -11623 21816 -11621
rect 21784 -11651 21786 -11623
rect 21786 -11651 21814 -11623
rect 21814 -11651 21816 -11623
rect 21784 -11653 21816 -11651
rect 21944 -11623 21976 -11621
rect 21944 -11651 21946 -11623
rect 21946 -11651 21974 -11623
rect 21974 -11651 21976 -11623
rect 21944 -11653 21976 -11651
rect 22104 -11623 22136 -11621
rect 22104 -11651 22106 -11623
rect 22106 -11651 22134 -11623
rect 22134 -11651 22136 -11623
rect 22104 -11653 22136 -11651
rect 22264 -11623 22296 -11621
rect 22264 -11651 22266 -11623
rect 22266 -11651 22294 -11623
rect 22294 -11651 22296 -11623
rect 22264 -11653 22296 -11651
rect 22424 -11623 22456 -11621
rect 22424 -11651 22426 -11623
rect 22426 -11651 22454 -11623
rect 22454 -11651 22456 -11623
rect 22424 -11653 22456 -11651
rect 22584 -11623 22616 -11621
rect 22584 -11651 22586 -11623
rect 22586 -11651 22614 -11623
rect 22614 -11651 22616 -11623
rect 22584 -11653 22616 -11651
rect 22744 -11623 22776 -11621
rect 22744 -11651 22746 -11623
rect 22746 -11651 22774 -11623
rect 22774 -11651 22776 -11623
rect 22744 -11653 22776 -11651
rect 22904 -11623 22936 -11621
rect 22904 -11651 22906 -11623
rect 22906 -11651 22934 -11623
rect 22934 -11651 22936 -11623
rect 22904 -11653 22936 -11651
rect 23064 -11623 23096 -11621
rect 23064 -11651 23066 -11623
rect 23066 -11651 23094 -11623
rect 23094 -11651 23096 -11623
rect 23064 -11653 23096 -11651
rect 23224 -11623 23256 -11621
rect 23224 -11651 23226 -11623
rect 23226 -11651 23254 -11623
rect 23254 -11651 23256 -11623
rect 23224 -11653 23256 -11651
rect 23384 -11623 23416 -11621
rect 23384 -11651 23386 -11623
rect 23386 -11651 23414 -11623
rect 23414 -11651 23416 -11623
rect 23384 -11653 23416 -11651
rect 23544 -11623 23576 -11621
rect 23544 -11651 23546 -11623
rect 23546 -11651 23574 -11623
rect 23574 -11651 23576 -11623
rect 23544 -11653 23576 -11651
rect 23704 -11623 23736 -11621
rect 23704 -11651 23706 -11623
rect 23706 -11651 23734 -11623
rect 23734 -11651 23736 -11623
rect 23704 -11653 23736 -11651
rect 23864 -11623 23896 -11621
rect 23864 -11651 23866 -11623
rect 23866 -11651 23894 -11623
rect 23894 -11651 23896 -11623
rect 23864 -11653 23896 -11651
rect 24024 -11623 24056 -11621
rect 24024 -11651 24026 -11623
rect 24026 -11651 24054 -11623
rect 24054 -11651 24056 -11623
rect 24024 -11653 24056 -11651
rect 24184 -11623 24216 -11621
rect 24184 -11651 24186 -11623
rect 24186 -11651 24214 -11623
rect 24214 -11651 24216 -11623
rect 24184 -11653 24216 -11651
rect 24344 -11623 24376 -11621
rect 24344 -11651 24346 -11623
rect 24346 -11651 24374 -11623
rect 24374 -11651 24376 -11623
rect 24344 -11653 24376 -11651
rect 24504 -11623 24536 -11621
rect 24504 -11651 24506 -11623
rect 24506 -11651 24534 -11623
rect 24534 -11651 24536 -11623
rect 24504 -11653 24536 -11651
rect 24664 -11623 24696 -11621
rect 24664 -11651 24666 -11623
rect 24666 -11651 24694 -11623
rect 24694 -11651 24696 -11623
rect 24664 -11653 24696 -11651
rect 21119 -11726 21151 -11724
rect 21119 -11754 21121 -11726
rect 21121 -11754 21149 -11726
rect 21149 -11754 21151 -11726
rect 21119 -11756 21151 -11754
rect 24852 -11726 24884 -11724
rect 24852 -11754 24854 -11726
rect 24854 -11754 24882 -11726
rect 24882 -11754 24884 -11726
rect 24852 -11756 24884 -11754
rect 21119 -11886 21151 -11884
rect 21119 -11914 21121 -11886
rect 21121 -11914 21149 -11886
rect 21149 -11914 21151 -11886
rect 21119 -11916 21151 -11914
rect 21119 -12046 21151 -12044
rect 21119 -12074 21121 -12046
rect 21121 -12074 21149 -12046
rect 21149 -12074 21151 -12046
rect 21119 -12076 21151 -12074
rect 21119 -12206 21151 -12204
rect 21119 -12234 21121 -12206
rect 21121 -12234 21149 -12206
rect 21149 -12234 21151 -12206
rect 21119 -12236 21151 -12234
rect 21119 -12366 21151 -12364
rect 21119 -12394 21121 -12366
rect 21121 -12394 21149 -12366
rect 21149 -12394 21151 -12366
rect 21119 -12396 21151 -12394
rect 21119 -12526 21151 -12524
rect 21119 -12554 21121 -12526
rect 21121 -12554 21149 -12526
rect 21149 -12554 21151 -12526
rect 21119 -12556 21151 -12554
rect 21119 -12686 21151 -12684
rect 21119 -12714 21121 -12686
rect 21121 -12714 21149 -12686
rect 21149 -12714 21151 -12686
rect 21119 -12716 21151 -12714
rect 21119 -12846 21151 -12844
rect 21119 -12874 21121 -12846
rect 21121 -12874 21149 -12846
rect 21149 -12874 21151 -12846
rect 21119 -12876 21151 -12874
rect 21119 -13006 21151 -13004
rect 21119 -13034 21121 -13006
rect 21121 -13034 21149 -13006
rect 21149 -13034 21151 -13006
rect 21119 -13036 21151 -13034
rect 21119 -13166 21151 -13164
rect 21119 -13194 21121 -13166
rect 21121 -13194 21149 -13166
rect 21149 -13194 21151 -13166
rect 21119 -13196 21151 -13194
rect 21119 -13326 21151 -13324
rect 21119 -13354 21121 -13326
rect 21121 -13354 21149 -13326
rect 21149 -13354 21151 -13326
rect 21119 -13356 21151 -13354
rect 21119 -13486 21151 -13484
rect 21119 -13514 21121 -13486
rect 21121 -13514 21149 -13486
rect 21149 -13514 21151 -13486
rect 21119 -13516 21151 -13514
rect 21119 -13646 21151 -13644
rect 21119 -13674 21121 -13646
rect 21121 -13674 21149 -13646
rect 21149 -13674 21151 -13646
rect 21119 -13676 21151 -13674
rect 21119 -13806 21151 -13804
rect 21119 -13834 21121 -13806
rect 21121 -13834 21149 -13806
rect 21149 -13834 21151 -13806
rect 21119 -13836 21151 -13834
rect 21119 -13966 21151 -13964
rect 21119 -13994 21121 -13966
rect 21121 -13994 21149 -13966
rect 21149 -13994 21151 -13966
rect 21119 -13996 21151 -13994
rect 21119 -14126 21151 -14124
rect 21119 -14154 21121 -14126
rect 21121 -14154 21149 -14126
rect 21149 -14154 21151 -14126
rect 21119 -14156 21151 -14154
rect 21119 -14286 21151 -14284
rect 21119 -14314 21121 -14286
rect 21121 -14314 21149 -14286
rect 21149 -14314 21151 -14286
rect 21119 -14316 21151 -14314
rect 21119 -14446 21151 -14444
rect 21119 -14474 21121 -14446
rect 21121 -14474 21149 -14446
rect 21149 -14474 21151 -14446
rect 21119 -14476 21151 -14474
rect 21119 -14606 21151 -14604
rect 21119 -14634 21121 -14606
rect 21121 -14634 21149 -14606
rect 21149 -14634 21151 -14606
rect 21119 -14636 21151 -14634
rect 21119 -14766 21151 -14764
rect 21119 -14794 21121 -14766
rect 21121 -14794 21149 -14766
rect 21149 -14794 21151 -14766
rect 21119 -14796 21151 -14794
rect 21119 -14926 21151 -14924
rect 21119 -14954 21121 -14926
rect 21121 -14954 21149 -14926
rect 21149 -14954 21151 -14926
rect 21119 -14956 21151 -14954
rect 21119 -15086 21151 -15084
rect 21119 -15114 21121 -15086
rect 21121 -15114 21149 -15086
rect 21149 -15114 21151 -15086
rect 21119 -15116 21151 -15114
rect 24852 -11886 24884 -11884
rect 24852 -11914 24854 -11886
rect 24854 -11914 24882 -11886
rect 24882 -11914 24884 -11886
rect 24852 -11916 24884 -11914
rect 24852 -12046 24884 -12044
rect 24852 -12074 24854 -12046
rect 24854 -12074 24882 -12046
rect 24882 -12074 24884 -12046
rect 24852 -12076 24884 -12074
rect 24852 -12206 24884 -12204
rect 24852 -12234 24854 -12206
rect 24854 -12234 24882 -12206
rect 24882 -12234 24884 -12206
rect 24852 -12236 24884 -12234
rect 24852 -12366 24884 -12364
rect 24852 -12394 24854 -12366
rect 24854 -12394 24882 -12366
rect 24882 -12394 24884 -12366
rect 24852 -12396 24884 -12394
rect 24852 -12526 24884 -12524
rect 24852 -12554 24854 -12526
rect 24854 -12554 24882 -12526
rect 24882 -12554 24884 -12526
rect 24852 -12556 24884 -12554
rect 24852 -12686 24884 -12684
rect 24852 -12714 24854 -12686
rect 24854 -12714 24882 -12686
rect 24882 -12714 24884 -12686
rect 24852 -12716 24884 -12714
rect 24852 -12846 24884 -12844
rect 24852 -12874 24854 -12846
rect 24854 -12874 24882 -12846
rect 24882 -12874 24884 -12846
rect 24852 -12876 24884 -12874
rect 24852 -13006 24884 -13004
rect 24852 -13034 24854 -13006
rect 24854 -13034 24882 -13006
rect 24882 -13034 24884 -13006
rect 24852 -13036 24884 -13034
rect 24852 -13166 24884 -13164
rect 24852 -13194 24854 -13166
rect 24854 -13194 24882 -13166
rect 24882 -13194 24884 -13166
rect 24852 -13196 24884 -13194
rect 24852 -13326 24884 -13324
rect 24852 -13354 24854 -13326
rect 24854 -13354 24882 -13326
rect 24882 -13354 24884 -13326
rect 24852 -13356 24884 -13354
rect 24852 -13486 24884 -13484
rect 24852 -13514 24854 -13486
rect 24854 -13514 24882 -13486
rect 24882 -13514 24884 -13486
rect 24852 -13516 24884 -13514
rect 24852 -13646 24884 -13644
rect 24852 -13674 24854 -13646
rect 24854 -13674 24882 -13646
rect 24882 -13674 24884 -13646
rect 24852 -13676 24884 -13674
rect 24852 -13806 24884 -13804
rect 24852 -13834 24854 -13806
rect 24854 -13834 24882 -13806
rect 24882 -13834 24884 -13806
rect 24852 -13836 24884 -13834
rect 24852 -13966 24884 -13964
rect 24852 -13994 24854 -13966
rect 24854 -13994 24882 -13966
rect 24882 -13994 24884 -13966
rect 24852 -13996 24884 -13994
rect 24852 -14126 24884 -14124
rect 24852 -14154 24854 -14126
rect 24854 -14154 24882 -14126
rect 24882 -14154 24884 -14126
rect 24852 -14156 24884 -14154
rect 24852 -14286 24884 -14284
rect 24852 -14314 24854 -14286
rect 24854 -14314 24882 -14286
rect 24882 -14314 24884 -14286
rect 24852 -14316 24884 -14314
rect 24852 -14446 24884 -14444
rect 24852 -14474 24854 -14446
rect 24854 -14474 24882 -14446
rect 24882 -14474 24884 -14446
rect 24852 -14476 24884 -14474
rect 24852 -14606 24884 -14604
rect 24852 -14634 24854 -14606
rect 24854 -14634 24882 -14606
rect 24882 -14634 24884 -14606
rect 24852 -14636 24884 -14634
rect 24852 -14766 24884 -14764
rect 24852 -14794 24854 -14766
rect 24854 -14794 24882 -14766
rect 24882 -14794 24884 -14766
rect 24852 -14796 24884 -14794
rect 24852 -14926 24884 -14924
rect 24852 -14954 24854 -14926
rect 24854 -14954 24882 -14926
rect 24882 -14954 24884 -14926
rect 24852 -14956 24884 -14954
rect 24852 -15086 24884 -15084
rect 24852 -15114 24854 -15086
rect 24854 -15114 24882 -15086
rect 24882 -15114 24884 -15086
rect 24852 -15116 24884 -15114
rect 21119 -15246 21151 -15244
rect 21119 -15274 21121 -15246
rect 21121 -15274 21149 -15246
rect 21149 -15274 21151 -15246
rect 21119 -15276 21151 -15274
rect 24852 -15246 24884 -15244
rect 24852 -15274 24854 -15246
rect 24854 -15274 24882 -15246
rect 24882 -15274 24884 -15246
rect 24852 -15276 24884 -15274
rect 21304 -15351 21336 -15349
rect 21304 -15379 21306 -15351
rect 21306 -15379 21334 -15351
rect 21334 -15379 21336 -15351
rect 21304 -15381 21336 -15379
rect 21464 -15351 21496 -15349
rect 21464 -15379 21466 -15351
rect 21466 -15379 21494 -15351
rect 21494 -15379 21496 -15351
rect 21464 -15381 21496 -15379
rect 21624 -15351 21656 -15349
rect 21624 -15379 21626 -15351
rect 21626 -15379 21654 -15351
rect 21654 -15379 21656 -15351
rect 21624 -15381 21656 -15379
rect 21784 -15351 21816 -15349
rect 21784 -15379 21786 -15351
rect 21786 -15379 21814 -15351
rect 21814 -15379 21816 -15351
rect 21784 -15381 21816 -15379
rect 21944 -15351 21976 -15349
rect 21944 -15379 21946 -15351
rect 21946 -15379 21974 -15351
rect 21974 -15379 21976 -15351
rect 21944 -15381 21976 -15379
rect 22104 -15351 22136 -15349
rect 22104 -15379 22106 -15351
rect 22106 -15379 22134 -15351
rect 22134 -15379 22136 -15351
rect 22104 -15381 22136 -15379
rect 22264 -15351 22296 -15349
rect 22264 -15379 22266 -15351
rect 22266 -15379 22294 -15351
rect 22294 -15379 22296 -15351
rect 22264 -15381 22296 -15379
rect 22424 -15351 22456 -15349
rect 22424 -15379 22426 -15351
rect 22426 -15379 22454 -15351
rect 22454 -15379 22456 -15351
rect 22424 -15381 22456 -15379
rect 22584 -15351 22616 -15349
rect 22584 -15379 22586 -15351
rect 22586 -15379 22614 -15351
rect 22614 -15379 22616 -15351
rect 22584 -15381 22616 -15379
rect 22744 -15351 22776 -15349
rect 22744 -15379 22746 -15351
rect 22746 -15379 22774 -15351
rect 22774 -15379 22776 -15351
rect 22744 -15381 22776 -15379
rect 22904 -15351 22936 -15349
rect 22904 -15379 22906 -15351
rect 22906 -15379 22934 -15351
rect 22934 -15379 22936 -15351
rect 22904 -15381 22936 -15379
rect 23064 -15351 23096 -15349
rect 23064 -15379 23066 -15351
rect 23066 -15379 23094 -15351
rect 23094 -15379 23096 -15351
rect 23064 -15381 23096 -15379
rect 23224 -15351 23256 -15349
rect 23224 -15379 23226 -15351
rect 23226 -15379 23254 -15351
rect 23254 -15379 23256 -15351
rect 23224 -15381 23256 -15379
rect 23384 -15351 23416 -15349
rect 23384 -15379 23386 -15351
rect 23386 -15379 23414 -15351
rect 23414 -15379 23416 -15351
rect 23384 -15381 23416 -15379
rect 23544 -15351 23576 -15349
rect 23544 -15379 23546 -15351
rect 23546 -15379 23574 -15351
rect 23574 -15379 23576 -15351
rect 23544 -15381 23576 -15379
rect 23704 -15351 23736 -15349
rect 23704 -15379 23706 -15351
rect 23706 -15379 23734 -15351
rect 23734 -15379 23736 -15351
rect 23704 -15381 23736 -15379
rect 23864 -15351 23896 -15349
rect 23864 -15379 23866 -15351
rect 23866 -15379 23894 -15351
rect 23894 -15379 23896 -15351
rect 23864 -15381 23896 -15379
rect 24024 -15351 24056 -15349
rect 24024 -15379 24026 -15351
rect 24026 -15379 24054 -15351
rect 24054 -15379 24056 -15351
rect 24024 -15381 24056 -15379
rect 24184 -15351 24216 -15349
rect 24184 -15379 24186 -15351
rect 24186 -15379 24214 -15351
rect 24214 -15379 24216 -15351
rect 24184 -15381 24216 -15379
rect 24344 -15351 24376 -15349
rect 24344 -15379 24346 -15351
rect 24346 -15379 24374 -15351
rect 24374 -15379 24376 -15351
rect 24344 -15381 24376 -15379
rect 24504 -15351 24536 -15349
rect 24504 -15379 24506 -15351
rect 24506 -15379 24534 -15351
rect 24534 -15379 24536 -15351
rect 24504 -15381 24536 -15379
rect 24664 -15351 24696 -15349
rect 24664 -15379 24666 -15351
rect 24666 -15379 24694 -15351
rect 24694 -15379 24696 -15351
rect 24664 -15381 24696 -15379
<< metal4 >>
rect 3000 9424 7000 9500
rect 3000 9319 3261 9424
rect 3000 9201 3073 9319
rect 3191 9306 3261 9319
rect 3379 9306 3421 9424
rect 3539 9306 3581 9424
rect 3699 9306 3741 9424
rect 3859 9306 3901 9424
rect 4019 9306 4061 9424
rect 4179 9306 4221 9424
rect 4339 9306 4381 9424
rect 4499 9306 4541 9424
rect 4659 9306 4701 9424
rect 4819 9306 4861 9424
rect 4979 9306 5021 9424
rect 5139 9306 5181 9424
rect 5299 9306 5341 9424
rect 5459 9306 5501 9424
rect 5619 9306 5661 9424
rect 5779 9306 5821 9424
rect 5939 9306 5981 9424
rect 6099 9306 6141 9424
rect 6259 9306 6301 9424
rect 6419 9306 6461 9424
rect 6579 9306 6621 9424
rect 6739 9319 7000 9424
rect 6739 9306 6806 9319
rect 3191 9230 6806 9306
rect 3191 9201 3270 9230
rect 3000 9159 3270 9201
rect 3000 9041 3073 9159
rect 3191 9041 3270 9159
rect 3000 8999 3270 9041
rect 3000 8881 3073 8999
rect 3191 8881 3270 8999
rect 3000 8839 3270 8881
rect 3000 8721 3073 8839
rect 3191 8721 3270 8839
rect 3000 8679 3270 8721
rect 3000 8561 3073 8679
rect 3191 8561 3270 8679
rect 3000 8519 3270 8561
rect 3000 8401 3073 8519
rect 3191 8401 3270 8519
rect 3000 8359 3270 8401
rect 3000 8241 3073 8359
rect 3191 8241 3270 8359
rect 3000 8199 3270 8241
rect 3000 8081 3073 8199
rect 3191 8081 3270 8199
rect 3000 8039 3270 8081
rect 3000 7921 3073 8039
rect 3191 7921 3270 8039
rect 3000 7879 3270 7921
rect 3000 7761 3073 7879
rect 3191 7761 3270 7879
rect 3000 7719 3270 7761
rect 3000 7601 3073 7719
rect 3191 7601 3270 7719
rect 3000 7559 3270 7601
rect 3000 7441 3073 7559
rect 3191 7441 3270 7559
rect 3000 7399 3270 7441
rect 3000 7281 3073 7399
rect 3191 7281 3270 7399
rect 3000 7239 3270 7281
rect 3000 7121 3073 7239
rect 3191 7121 3270 7239
rect 3000 7079 3270 7121
rect 3000 6961 3073 7079
rect 3191 6961 3270 7079
rect 3000 6919 3270 6961
rect 3000 6801 3073 6919
rect 3191 6801 3270 6919
rect 3000 6759 3270 6801
rect 3000 6641 3073 6759
rect 3191 6641 3270 6759
rect 3000 6599 3270 6641
rect 3000 6481 3073 6599
rect 3191 6481 3270 6599
rect 3000 6439 3270 6481
rect 3000 6321 3073 6439
rect 3191 6321 3270 6439
rect 3000 6279 3270 6321
rect 3000 6161 3073 6279
rect 3191 6161 3270 6279
rect 3000 6119 3270 6161
rect 3000 6001 3073 6119
rect 3191 6001 3270 6119
rect 3000 5959 3270 6001
rect 3000 5841 3073 5959
rect 3191 5841 3270 5959
rect 3000 5799 3270 5841
rect 3000 5681 3073 5799
rect 3191 5770 3270 5799
rect 6730 9201 6806 9230
rect 6924 9201 7000 9319
rect 6730 9159 7000 9201
rect 6730 9041 6806 9159
rect 6924 9041 7000 9159
rect 6730 8999 7000 9041
rect 6730 8881 6806 8999
rect 6924 8881 7000 8999
rect 6730 8839 7000 8881
rect 6730 8721 6806 8839
rect 6924 8721 7000 8839
rect 6730 8679 7000 8721
rect 6730 8561 6806 8679
rect 6924 8561 7000 8679
rect 6730 8519 7000 8561
rect 6730 8401 6806 8519
rect 6924 8401 7000 8519
rect 6730 8359 7000 8401
rect 6730 8241 6806 8359
rect 6924 8241 7000 8359
rect 6730 8199 7000 8241
rect 6730 8081 6806 8199
rect 6924 8081 7000 8199
rect 6730 8039 7000 8081
rect 6730 7921 6806 8039
rect 6924 7921 7000 8039
rect 6730 7879 7000 7921
rect 6730 7761 6806 7879
rect 6924 7761 7000 7879
rect 6730 7719 7000 7761
rect 6730 7601 6806 7719
rect 6924 7601 7000 7719
rect 6730 7559 7000 7601
rect 6730 7441 6806 7559
rect 6924 7441 7000 7559
rect 6730 7399 7000 7441
rect 6730 7281 6806 7399
rect 6924 7281 7000 7399
rect 6730 7239 7000 7281
rect 6730 7121 6806 7239
rect 6924 7121 7000 7239
rect 6730 7079 7000 7121
rect 6730 6961 6806 7079
rect 6924 6961 7000 7079
rect 6730 6919 7000 6961
rect 6730 6801 6806 6919
rect 6924 6801 7000 6919
rect 6730 6759 7000 6801
rect 6730 6641 6806 6759
rect 6924 6641 7000 6759
rect 6730 6599 7000 6641
rect 6730 6481 6806 6599
rect 6924 6481 7000 6599
rect 6730 6439 7000 6481
rect 6730 6321 6806 6439
rect 6924 6321 7000 6439
rect 6730 6279 7000 6321
rect 6730 6161 6806 6279
rect 6924 6161 7000 6279
rect 6730 6119 7000 6161
rect 6730 6001 6806 6119
rect 6924 6001 7000 6119
rect 6730 5959 7000 6001
rect 6730 5841 6806 5959
rect 6924 5841 7000 5959
rect 6730 5799 7000 5841
rect 6730 5770 6806 5799
rect 3191 5696 6806 5770
rect 3191 5681 3261 5696
rect 3000 5578 3261 5681
rect 3379 5578 3421 5696
rect 3539 5578 3581 5696
rect 3699 5578 3741 5696
rect 3859 5578 3901 5696
rect 4019 5578 4061 5696
rect 4179 5578 4221 5696
rect 4339 5578 4381 5696
rect 4499 5578 4541 5696
rect 4659 5578 4701 5696
rect 4819 5578 4861 5696
rect 4979 5578 5021 5696
rect 5139 5578 5181 5696
rect 5299 5578 5341 5696
rect 5459 5578 5501 5696
rect 5619 5578 5661 5696
rect 5779 5578 5821 5696
rect 5939 5578 5981 5696
rect 6099 5578 6141 5696
rect 6259 5578 6301 5696
rect 6419 5578 6461 5696
rect 6579 5578 6621 5696
rect 6739 5681 6806 5696
rect 6924 5681 7000 5799
rect 6739 5578 7000 5681
rect 3000 5500 7000 5578
rect 9000 9424 13000 9500
rect 9000 9319 9261 9424
rect 9000 9201 9073 9319
rect 9191 9306 9261 9319
rect 9379 9306 9421 9424
rect 9539 9306 9581 9424
rect 9699 9306 9741 9424
rect 9859 9306 9901 9424
rect 10019 9306 10061 9424
rect 10179 9306 10221 9424
rect 10339 9306 10381 9424
rect 10499 9306 10541 9424
rect 10659 9306 10701 9424
rect 10819 9306 10861 9424
rect 10979 9306 11021 9424
rect 11139 9306 11181 9424
rect 11299 9306 11341 9424
rect 11459 9306 11501 9424
rect 11619 9306 11661 9424
rect 11779 9306 11821 9424
rect 11939 9306 11981 9424
rect 12099 9306 12141 9424
rect 12259 9306 12301 9424
rect 12419 9306 12461 9424
rect 12579 9306 12621 9424
rect 12739 9319 13000 9424
rect 12739 9306 12806 9319
rect 9191 9230 12806 9306
rect 9191 9201 9270 9230
rect 9000 9159 9270 9201
rect 9000 9041 9073 9159
rect 9191 9041 9270 9159
rect 9000 8999 9270 9041
rect 9000 8881 9073 8999
rect 9191 8881 9270 8999
rect 9000 8839 9270 8881
rect 9000 8721 9073 8839
rect 9191 8721 9270 8839
rect 9000 8679 9270 8721
rect 9000 8561 9073 8679
rect 9191 8561 9270 8679
rect 9000 8519 9270 8561
rect 9000 8401 9073 8519
rect 9191 8401 9270 8519
rect 9000 8359 9270 8401
rect 9000 8241 9073 8359
rect 9191 8241 9270 8359
rect 9000 8199 9270 8241
rect 9000 8081 9073 8199
rect 9191 8081 9270 8199
rect 9000 8039 9270 8081
rect 9000 7921 9073 8039
rect 9191 7921 9270 8039
rect 9000 7879 9270 7921
rect 9000 7761 9073 7879
rect 9191 7761 9270 7879
rect 9000 7719 9270 7761
rect 9000 7601 9073 7719
rect 9191 7601 9270 7719
rect 9000 7559 9270 7601
rect 9000 7441 9073 7559
rect 9191 7441 9270 7559
rect 9000 7399 9270 7441
rect 9000 7281 9073 7399
rect 9191 7281 9270 7399
rect 9000 7239 9270 7281
rect 9000 7121 9073 7239
rect 9191 7121 9270 7239
rect 9000 7079 9270 7121
rect 9000 6961 9073 7079
rect 9191 6961 9270 7079
rect 9000 6919 9270 6961
rect 9000 6801 9073 6919
rect 9191 6801 9270 6919
rect 9000 6759 9270 6801
rect 9000 6641 9073 6759
rect 9191 6641 9270 6759
rect 9000 6599 9270 6641
rect 9000 6481 9073 6599
rect 9191 6481 9270 6599
rect 9000 6439 9270 6481
rect 9000 6321 9073 6439
rect 9191 6321 9270 6439
rect 9000 6279 9270 6321
rect 9000 6161 9073 6279
rect 9191 6161 9270 6279
rect 9000 6119 9270 6161
rect 9000 6001 9073 6119
rect 9191 6001 9270 6119
rect 9000 5959 9270 6001
rect 9000 5841 9073 5959
rect 9191 5841 9270 5959
rect 9000 5799 9270 5841
rect 9000 5681 9073 5799
rect 9191 5770 9270 5799
rect 12730 9201 12806 9230
rect 12924 9201 13000 9319
rect 12730 9159 13000 9201
rect 12730 9041 12806 9159
rect 12924 9041 13000 9159
rect 12730 8999 13000 9041
rect 12730 8881 12806 8999
rect 12924 8881 13000 8999
rect 12730 8839 13000 8881
rect 12730 8721 12806 8839
rect 12924 8721 13000 8839
rect 12730 8679 13000 8721
rect 12730 8561 12806 8679
rect 12924 8561 13000 8679
rect 12730 8519 13000 8561
rect 12730 8401 12806 8519
rect 12924 8401 13000 8519
rect 12730 8359 13000 8401
rect 12730 8241 12806 8359
rect 12924 8241 13000 8359
rect 12730 8199 13000 8241
rect 12730 8081 12806 8199
rect 12924 8081 13000 8199
rect 12730 8039 13000 8081
rect 12730 7921 12806 8039
rect 12924 7921 13000 8039
rect 12730 7879 13000 7921
rect 12730 7761 12806 7879
rect 12924 7761 13000 7879
rect 12730 7719 13000 7761
rect 12730 7601 12806 7719
rect 12924 7601 13000 7719
rect 12730 7559 13000 7601
rect 12730 7441 12806 7559
rect 12924 7441 13000 7559
rect 12730 7399 13000 7441
rect 12730 7281 12806 7399
rect 12924 7281 13000 7399
rect 12730 7239 13000 7281
rect 12730 7121 12806 7239
rect 12924 7121 13000 7239
rect 12730 7079 13000 7121
rect 12730 6961 12806 7079
rect 12924 6961 13000 7079
rect 12730 6919 13000 6961
rect 12730 6801 12806 6919
rect 12924 6801 13000 6919
rect 12730 6759 13000 6801
rect 12730 6641 12806 6759
rect 12924 6641 13000 6759
rect 12730 6599 13000 6641
rect 12730 6481 12806 6599
rect 12924 6481 13000 6599
rect 12730 6439 13000 6481
rect 12730 6321 12806 6439
rect 12924 6321 13000 6439
rect 12730 6279 13000 6321
rect 12730 6161 12806 6279
rect 12924 6161 13000 6279
rect 12730 6119 13000 6161
rect 12730 6001 12806 6119
rect 12924 6001 13000 6119
rect 12730 5959 13000 6001
rect 12730 5841 12806 5959
rect 12924 5841 13000 5959
rect 12730 5799 13000 5841
rect 12730 5770 12806 5799
rect 9191 5696 12806 5770
rect 9191 5681 9261 5696
rect 9000 5578 9261 5681
rect 9379 5578 9421 5696
rect 9539 5578 9581 5696
rect 9699 5578 9741 5696
rect 9859 5578 9901 5696
rect 10019 5578 10061 5696
rect 10179 5578 10221 5696
rect 10339 5578 10381 5696
rect 10499 5578 10541 5696
rect 10659 5578 10701 5696
rect 10819 5578 10861 5696
rect 10979 5578 11021 5696
rect 11139 5578 11181 5696
rect 11299 5578 11341 5696
rect 11459 5578 11501 5696
rect 11619 5578 11661 5696
rect 11779 5578 11821 5696
rect 11939 5578 11981 5696
rect 12099 5578 12141 5696
rect 12259 5578 12301 5696
rect 12419 5578 12461 5696
rect 12579 5578 12621 5696
rect 12739 5681 12806 5696
rect 12924 5681 13000 5799
rect 12739 5578 13000 5681
rect 9000 5500 13000 5578
rect 15000 9424 19000 9500
rect 15000 9319 15261 9424
rect 15000 9201 15073 9319
rect 15191 9306 15261 9319
rect 15379 9306 15421 9424
rect 15539 9306 15581 9424
rect 15699 9306 15741 9424
rect 15859 9306 15901 9424
rect 16019 9306 16061 9424
rect 16179 9306 16221 9424
rect 16339 9306 16381 9424
rect 16499 9306 16541 9424
rect 16659 9306 16701 9424
rect 16819 9306 16861 9424
rect 16979 9306 17021 9424
rect 17139 9306 17181 9424
rect 17299 9306 17341 9424
rect 17459 9306 17501 9424
rect 17619 9306 17661 9424
rect 17779 9306 17821 9424
rect 17939 9306 17981 9424
rect 18099 9306 18141 9424
rect 18259 9306 18301 9424
rect 18419 9306 18461 9424
rect 18579 9306 18621 9424
rect 18739 9319 19000 9424
rect 18739 9306 18806 9319
rect 15191 9230 18806 9306
rect 15191 9201 15270 9230
rect 15000 9159 15270 9201
rect 15000 9041 15073 9159
rect 15191 9041 15270 9159
rect 15000 8999 15270 9041
rect 15000 8881 15073 8999
rect 15191 8881 15270 8999
rect 15000 8839 15270 8881
rect 15000 8721 15073 8839
rect 15191 8721 15270 8839
rect 15000 8679 15270 8721
rect 15000 8561 15073 8679
rect 15191 8561 15270 8679
rect 15000 8519 15270 8561
rect 15000 8401 15073 8519
rect 15191 8401 15270 8519
rect 15000 8359 15270 8401
rect 15000 8241 15073 8359
rect 15191 8241 15270 8359
rect 15000 8199 15270 8241
rect 15000 8081 15073 8199
rect 15191 8081 15270 8199
rect 15000 8039 15270 8081
rect 15000 7921 15073 8039
rect 15191 7921 15270 8039
rect 15000 7879 15270 7921
rect 15000 7761 15073 7879
rect 15191 7761 15270 7879
rect 15000 7719 15270 7761
rect 15000 7601 15073 7719
rect 15191 7601 15270 7719
rect 15000 7559 15270 7601
rect 15000 7441 15073 7559
rect 15191 7441 15270 7559
rect 15000 7399 15270 7441
rect 15000 7281 15073 7399
rect 15191 7281 15270 7399
rect 15000 7239 15270 7281
rect 15000 7121 15073 7239
rect 15191 7121 15270 7239
rect 15000 7079 15270 7121
rect 15000 6961 15073 7079
rect 15191 6961 15270 7079
rect 15000 6919 15270 6961
rect 15000 6801 15073 6919
rect 15191 6801 15270 6919
rect 15000 6759 15270 6801
rect 15000 6641 15073 6759
rect 15191 6641 15270 6759
rect 15000 6599 15270 6641
rect 15000 6481 15073 6599
rect 15191 6481 15270 6599
rect 15000 6439 15270 6481
rect 15000 6321 15073 6439
rect 15191 6321 15270 6439
rect 15000 6279 15270 6321
rect 15000 6161 15073 6279
rect 15191 6161 15270 6279
rect 15000 6119 15270 6161
rect 15000 6001 15073 6119
rect 15191 6001 15270 6119
rect 15000 5959 15270 6001
rect 15000 5841 15073 5959
rect 15191 5841 15270 5959
rect 15000 5799 15270 5841
rect 15000 5681 15073 5799
rect 15191 5770 15270 5799
rect 18730 9201 18806 9230
rect 18924 9201 19000 9319
rect 18730 9159 19000 9201
rect 18730 9041 18806 9159
rect 18924 9041 19000 9159
rect 18730 8999 19000 9041
rect 18730 8881 18806 8999
rect 18924 8881 19000 8999
rect 18730 8839 19000 8881
rect 18730 8721 18806 8839
rect 18924 8721 19000 8839
rect 18730 8679 19000 8721
rect 18730 8561 18806 8679
rect 18924 8561 19000 8679
rect 18730 8519 19000 8561
rect 18730 8401 18806 8519
rect 18924 8401 19000 8519
rect 18730 8359 19000 8401
rect 18730 8241 18806 8359
rect 18924 8241 19000 8359
rect 18730 8199 19000 8241
rect 18730 8081 18806 8199
rect 18924 8081 19000 8199
rect 18730 8039 19000 8081
rect 18730 7921 18806 8039
rect 18924 7921 19000 8039
rect 18730 7879 19000 7921
rect 18730 7761 18806 7879
rect 18924 7761 19000 7879
rect 18730 7719 19000 7761
rect 18730 7601 18806 7719
rect 18924 7601 19000 7719
rect 18730 7559 19000 7601
rect 18730 7441 18806 7559
rect 18924 7441 19000 7559
rect 18730 7399 19000 7441
rect 18730 7281 18806 7399
rect 18924 7281 19000 7399
rect 18730 7239 19000 7281
rect 18730 7121 18806 7239
rect 18924 7121 19000 7239
rect 18730 7079 19000 7121
rect 18730 6961 18806 7079
rect 18924 6961 19000 7079
rect 18730 6919 19000 6961
rect 18730 6801 18806 6919
rect 18924 6801 19000 6919
rect 18730 6759 19000 6801
rect 18730 6641 18806 6759
rect 18924 6641 19000 6759
rect 18730 6599 19000 6641
rect 18730 6481 18806 6599
rect 18924 6481 19000 6599
rect 18730 6439 19000 6481
rect 18730 6321 18806 6439
rect 18924 6321 19000 6439
rect 18730 6279 19000 6321
rect 18730 6161 18806 6279
rect 18924 6161 19000 6279
rect 18730 6119 19000 6161
rect 18730 6001 18806 6119
rect 18924 6001 19000 6119
rect 18730 5959 19000 6001
rect 18730 5841 18806 5959
rect 18924 5841 19000 5959
rect 18730 5799 19000 5841
rect 18730 5770 18806 5799
rect 15191 5696 18806 5770
rect 15191 5681 15261 5696
rect 15000 5578 15261 5681
rect 15379 5578 15421 5696
rect 15539 5578 15581 5696
rect 15699 5578 15741 5696
rect 15859 5578 15901 5696
rect 16019 5578 16061 5696
rect 16179 5578 16221 5696
rect 16339 5578 16381 5696
rect 16499 5578 16541 5696
rect 16659 5578 16701 5696
rect 16819 5578 16861 5696
rect 16979 5578 17021 5696
rect 17139 5578 17181 5696
rect 17299 5578 17341 5696
rect 17459 5578 17501 5696
rect 17619 5578 17661 5696
rect 17779 5578 17821 5696
rect 17939 5578 17981 5696
rect 18099 5578 18141 5696
rect 18259 5578 18301 5696
rect 18419 5578 18461 5696
rect 18579 5578 18621 5696
rect 18739 5681 18806 5696
rect 18924 5681 19000 5799
rect 18739 5578 19000 5681
rect 15000 5500 19000 5578
rect 21000 9424 25000 9500
rect 21000 9319 21261 9424
rect 21000 9201 21073 9319
rect 21191 9306 21261 9319
rect 21379 9306 21421 9424
rect 21539 9306 21581 9424
rect 21699 9306 21741 9424
rect 21859 9306 21901 9424
rect 22019 9306 22061 9424
rect 22179 9306 22221 9424
rect 22339 9306 22381 9424
rect 22499 9306 22541 9424
rect 22659 9306 22701 9424
rect 22819 9306 22861 9424
rect 22979 9306 23021 9424
rect 23139 9306 23181 9424
rect 23299 9306 23341 9424
rect 23459 9306 23501 9424
rect 23619 9306 23661 9424
rect 23779 9306 23821 9424
rect 23939 9306 23981 9424
rect 24099 9306 24141 9424
rect 24259 9306 24301 9424
rect 24419 9306 24461 9424
rect 24579 9306 24621 9424
rect 24739 9319 25000 9424
rect 24739 9306 24806 9319
rect 21191 9230 24806 9306
rect 21191 9201 21270 9230
rect 21000 9159 21270 9201
rect 21000 9041 21073 9159
rect 21191 9041 21270 9159
rect 21000 8999 21270 9041
rect 21000 8881 21073 8999
rect 21191 8881 21270 8999
rect 21000 8839 21270 8881
rect 21000 8721 21073 8839
rect 21191 8721 21270 8839
rect 21000 8679 21270 8721
rect 21000 8561 21073 8679
rect 21191 8561 21270 8679
rect 21000 8519 21270 8561
rect 21000 8401 21073 8519
rect 21191 8401 21270 8519
rect 21000 8359 21270 8401
rect 21000 8241 21073 8359
rect 21191 8241 21270 8359
rect 21000 8199 21270 8241
rect 21000 8081 21073 8199
rect 21191 8081 21270 8199
rect 21000 8039 21270 8081
rect 21000 7921 21073 8039
rect 21191 7921 21270 8039
rect 21000 7879 21270 7921
rect 21000 7761 21073 7879
rect 21191 7761 21270 7879
rect 21000 7719 21270 7761
rect 21000 7601 21073 7719
rect 21191 7601 21270 7719
rect 21000 7559 21270 7601
rect 21000 7441 21073 7559
rect 21191 7441 21270 7559
rect 21000 7399 21270 7441
rect 21000 7281 21073 7399
rect 21191 7281 21270 7399
rect 21000 7239 21270 7281
rect 21000 7121 21073 7239
rect 21191 7121 21270 7239
rect 21000 7079 21270 7121
rect 21000 6961 21073 7079
rect 21191 6961 21270 7079
rect 21000 6919 21270 6961
rect 21000 6801 21073 6919
rect 21191 6801 21270 6919
rect 21000 6759 21270 6801
rect 21000 6641 21073 6759
rect 21191 6641 21270 6759
rect 21000 6599 21270 6641
rect 21000 6481 21073 6599
rect 21191 6481 21270 6599
rect 21000 6439 21270 6481
rect 21000 6321 21073 6439
rect 21191 6321 21270 6439
rect 21000 6279 21270 6321
rect 21000 6161 21073 6279
rect 21191 6161 21270 6279
rect 21000 6119 21270 6161
rect 21000 6001 21073 6119
rect 21191 6001 21270 6119
rect 21000 5959 21270 6001
rect 21000 5841 21073 5959
rect 21191 5841 21270 5959
rect 21000 5799 21270 5841
rect 21000 5681 21073 5799
rect 21191 5770 21270 5799
rect 24730 9201 24806 9230
rect 24924 9201 25000 9319
rect 24730 9159 25000 9201
rect 24730 9041 24806 9159
rect 24924 9041 25000 9159
rect 24730 8999 25000 9041
rect 24730 8881 24806 8999
rect 24924 8881 25000 8999
rect 24730 8839 25000 8881
rect 24730 8721 24806 8839
rect 24924 8721 25000 8839
rect 24730 8679 25000 8721
rect 24730 8561 24806 8679
rect 24924 8561 25000 8679
rect 24730 8519 25000 8561
rect 24730 8401 24806 8519
rect 24924 8401 25000 8519
rect 24730 8359 25000 8401
rect 24730 8241 24806 8359
rect 24924 8241 25000 8359
rect 24730 8199 25000 8241
rect 24730 8081 24806 8199
rect 24924 8081 25000 8199
rect 24730 8039 25000 8081
rect 24730 7921 24806 8039
rect 24924 7921 25000 8039
rect 24730 7879 25000 7921
rect 24730 7761 24806 7879
rect 24924 7761 25000 7879
rect 24730 7719 25000 7761
rect 24730 7601 24806 7719
rect 24924 7601 25000 7719
rect 24730 7559 25000 7601
rect 24730 7441 24806 7559
rect 24924 7441 25000 7559
rect 24730 7399 25000 7441
rect 24730 7281 24806 7399
rect 24924 7281 25000 7399
rect 24730 7239 25000 7281
rect 24730 7121 24806 7239
rect 24924 7121 25000 7239
rect 24730 7079 25000 7121
rect 24730 6961 24806 7079
rect 24924 6961 25000 7079
rect 24730 6919 25000 6961
rect 24730 6801 24806 6919
rect 24924 6801 25000 6919
rect 24730 6759 25000 6801
rect 24730 6641 24806 6759
rect 24924 6641 25000 6759
rect 24730 6599 25000 6641
rect 24730 6481 24806 6599
rect 24924 6481 25000 6599
rect 24730 6439 25000 6481
rect 24730 6321 24806 6439
rect 24924 6321 25000 6439
rect 24730 6279 25000 6321
rect 24730 6161 24806 6279
rect 24924 6161 25000 6279
rect 24730 6119 25000 6161
rect 24730 6001 24806 6119
rect 24924 6001 25000 6119
rect 24730 5959 25000 6001
rect 24730 5841 24806 5959
rect 24924 5841 25000 5959
rect 24730 5799 25000 5841
rect 24730 5770 24806 5799
rect 21191 5696 24806 5770
rect 21191 5681 21261 5696
rect 21000 5578 21261 5681
rect 21379 5578 21421 5696
rect 21539 5578 21581 5696
rect 21699 5578 21741 5696
rect 21859 5578 21901 5696
rect 22019 5578 22061 5696
rect 22179 5578 22221 5696
rect 22339 5578 22381 5696
rect 22499 5578 22541 5696
rect 22659 5578 22701 5696
rect 22819 5578 22861 5696
rect 22979 5578 23021 5696
rect 23139 5578 23181 5696
rect 23299 5578 23341 5696
rect 23459 5578 23501 5696
rect 23619 5578 23661 5696
rect 23779 5578 23821 5696
rect 23939 5578 23981 5696
rect 24099 5578 24141 5696
rect 24259 5578 24301 5696
rect 24419 5578 24461 5696
rect 24579 5578 24621 5696
rect 24739 5681 24806 5696
rect 24924 5681 25000 5799
rect 24739 5578 25000 5681
rect 21000 5500 25000 5578
rect 6250 5350 6550 5450
rect 6750 5400 6850 5450
rect 6700 5350 6900 5400
rect 5850 5200 6150 5300
rect 6350 5150 6450 5350
rect 6650 5300 6950 5350
rect 11650 5300 11750 5450
rect 11850 5350 12150 5450
rect 12250 5350 12350 5450
rect 12450 5350 12550 5450
rect 12750 5400 12850 5450
rect 12700 5350 12900 5400
rect 18650 5350 18950 5450
rect 24650 5350 24950 5450
rect 12050 5300 12150 5350
rect 6250 5050 6550 5150
rect 6650 5050 6750 5300
rect 6850 5050 6950 5300
rect 11500 5200 11750 5300
rect 11900 5200 12150 5300
rect 12300 5250 12550 5350
rect 11650 5150 11750 5200
rect 12050 5150 12150 5200
rect 11450 5050 11750 5150
rect 11850 5050 12150 5150
rect 12250 5150 12350 5250
rect 12450 5150 12550 5250
rect 12250 5100 12550 5150
rect 12300 5050 12550 5100
rect 12650 5300 12950 5350
rect 12650 5050 12750 5300
rect 12850 5050 12950 5300
rect 18650 5300 18750 5350
rect 24650 5300 24750 5350
rect 18650 5250 18900 5300
rect 24650 5250 24900 5300
rect 18700 5200 18950 5250
rect 24700 5200 24950 5250
rect 18850 5150 18950 5200
rect 24850 5150 24950 5200
rect 18650 5050 18950 5150
rect 24650 5050 24950 5150
rect 18650 4950 18950 5000
rect 6300 3900 6500 3950
rect 6750 3900 6850 3950
rect 5950 3800 6050 3900
rect 6250 3850 6550 3900
rect 6700 3850 6900 3900
rect 5850 3700 6150 3800
rect 5950 3600 6050 3700
rect 6250 3650 6350 3850
rect 6450 3650 6550 3850
rect 6250 3600 6550 3650
rect 6650 3800 6950 3850
rect 11950 3800 12050 3900
rect 12250 3850 12550 3950
rect 12750 3900 12850 3950
rect 12700 3850 12900 3900
rect 17850 3850 18150 3950
rect 18250 3850 18550 3950
rect 18750 3900 18850 3950
rect 23900 3900 24150 3950
rect 24300 3900 24550 3950
rect 24750 3900 24850 3950
rect 18700 3850 18900 3900
rect 23850 3850 24150 3900
rect 6300 3550 6500 3600
rect 6650 3550 6750 3800
rect 6850 3550 6950 3800
rect 11850 3700 12150 3800
rect 11950 3600 12050 3700
rect 12350 3650 12450 3850
rect 12650 3800 12950 3850
rect 12250 3550 12550 3650
rect 12650 3550 12750 3800
rect 12850 3550 12950 3800
rect 17850 3800 17950 3850
rect 18250 3800 18350 3850
rect 18650 3800 18950 3850
rect 17850 3750 18100 3800
rect 18250 3750 18500 3800
rect 17900 3700 18150 3750
rect 18300 3700 18550 3750
rect 18050 3650 18150 3700
rect 18450 3650 18550 3700
rect 17850 3550 18150 3650
rect 18250 3550 18550 3650
rect 18650 3550 18750 3800
rect 18850 3550 18950 3800
rect 23850 3650 23950 3850
rect 24050 3650 24150 3850
rect 23850 3600 24150 3650
rect 24250 3850 24550 3900
rect 24700 3850 24900 3900
rect 24250 3650 24350 3850
rect 24450 3650 24550 3850
rect 24250 3600 24550 3650
rect 23900 3550 24150 3600
rect 24300 3550 24550 3600
rect 24650 3800 24950 3850
rect 24650 3550 24750 3800
rect 24850 3550 24950 3800
rect 3000 3424 7000 3500
rect 3000 3319 3261 3424
rect 3000 3201 3073 3319
rect 3191 3306 3261 3319
rect 3379 3306 3421 3424
rect 3539 3306 3581 3424
rect 3699 3306 3741 3424
rect 3859 3306 3901 3424
rect 4019 3306 4061 3424
rect 4179 3306 4221 3424
rect 4339 3306 4381 3424
rect 4499 3306 4541 3424
rect 4659 3306 4701 3424
rect 4819 3306 4861 3424
rect 4979 3306 5021 3424
rect 5139 3306 5181 3424
rect 5299 3306 5341 3424
rect 5459 3306 5501 3424
rect 5619 3306 5661 3424
rect 5779 3306 5821 3424
rect 5939 3306 5981 3424
rect 6099 3306 6141 3424
rect 6259 3306 6301 3424
rect 6419 3306 6461 3424
rect 6579 3306 6621 3424
rect 6739 3319 7000 3424
rect 6739 3306 6806 3319
rect 3191 3230 6806 3306
rect 3191 3201 3270 3230
rect 3000 3159 3270 3201
rect 3000 3041 3073 3159
rect 3191 3041 3270 3159
rect 3000 2999 3270 3041
rect 3000 2881 3073 2999
rect 3191 2881 3270 2999
rect 3000 2839 3270 2881
rect 3000 2721 3073 2839
rect 3191 2721 3270 2839
rect 3000 2679 3270 2721
rect 3000 2561 3073 2679
rect 3191 2561 3270 2679
rect 3000 2519 3270 2561
rect 3000 2401 3073 2519
rect 3191 2401 3270 2519
rect 3000 2359 3270 2401
rect 3000 2241 3073 2359
rect 3191 2241 3270 2359
rect 3000 2199 3270 2241
rect 3000 2081 3073 2199
rect 3191 2081 3270 2199
rect 3000 2039 3270 2081
rect 3000 1921 3073 2039
rect 3191 1921 3270 2039
rect 3000 1879 3270 1921
rect 3000 1761 3073 1879
rect 3191 1761 3270 1879
rect 3000 1719 3270 1761
rect 3000 1601 3073 1719
rect 3191 1601 3270 1719
rect 3000 1559 3270 1601
rect 3000 1441 3073 1559
rect 3191 1441 3270 1559
rect 3000 1399 3270 1441
rect 3000 1281 3073 1399
rect 3191 1281 3270 1399
rect 3000 1239 3270 1281
rect 3000 1121 3073 1239
rect 3191 1121 3270 1239
rect 3000 1079 3270 1121
rect 3000 961 3073 1079
rect 3191 961 3270 1079
rect 3000 919 3270 961
rect 3000 801 3073 919
rect 3191 801 3270 919
rect 3000 759 3270 801
rect 3000 641 3073 759
rect 3191 641 3270 759
rect 3000 599 3270 641
rect 3000 481 3073 599
rect 3191 481 3270 599
rect 3000 439 3270 481
rect 3000 321 3073 439
rect 3191 321 3270 439
rect 3000 279 3270 321
rect 3000 161 3073 279
rect 3191 161 3270 279
rect 3000 119 3270 161
rect 3000 1 3073 119
rect 3191 1 3270 119
rect 3000 -41 3270 1
rect 3000 -159 3073 -41
rect 3191 -159 3270 -41
rect 3000 -201 3270 -159
rect 3000 -319 3073 -201
rect 3191 -230 3270 -201
rect 6730 3201 6806 3230
rect 6924 3201 7000 3319
rect 6730 3159 7000 3201
rect 6730 3041 6806 3159
rect 6924 3041 7000 3159
rect 6730 2999 7000 3041
rect 6730 2881 6806 2999
rect 6924 2881 7000 2999
rect 6730 2839 7000 2881
rect 6730 2721 6806 2839
rect 6924 2721 7000 2839
rect 6730 2679 7000 2721
rect 6730 2561 6806 2679
rect 6924 2561 7000 2679
rect 6730 2519 7000 2561
rect 6730 2401 6806 2519
rect 6924 2401 7000 2519
rect 6730 2359 7000 2401
rect 6730 2241 6806 2359
rect 6924 2241 7000 2359
rect 6730 2199 7000 2241
rect 6730 2081 6806 2199
rect 6924 2081 7000 2199
rect 6730 2039 7000 2081
rect 6730 1921 6806 2039
rect 6924 1921 7000 2039
rect 6730 1879 7000 1921
rect 6730 1761 6806 1879
rect 6924 1761 7000 1879
rect 6730 1719 7000 1761
rect 6730 1601 6806 1719
rect 6924 1601 7000 1719
rect 6730 1559 7000 1601
rect 6730 1441 6806 1559
rect 6924 1441 7000 1559
rect 6730 1399 7000 1441
rect 6730 1281 6806 1399
rect 6924 1281 7000 1399
rect 6730 1239 7000 1281
rect 6730 1121 6806 1239
rect 6924 1121 7000 1239
rect 6730 1079 7000 1121
rect 6730 961 6806 1079
rect 6924 961 7000 1079
rect 6730 919 7000 961
rect 6730 801 6806 919
rect 6924 801 7000 919
rect 6730 759 7000 801
rect 6730 641 6806 759
rect 6924 641 7000 759
rect 6730 599 7000 641
rect 6730 481 6806 599
rect 6924 481 7000 599
rect 6730 439 7000 481
rect 6730 321 6806 439
rect 6924 321 7000 439
rect 6730 279 7000 321
rect 6730 161 6806 279
rect 6924 161 7000 279
rect 6730 119 7000 161
rect 6730 1 6806 119
rect 6924 1 7000 119
rect 6730 -41 7000 1
rect 6730 -159 6806 -41
rect 6924 -159 7000 -41
rect 6730 -201 7000 -159
rect 6730 -230 6806 -201
rect 3191 -304 6806 -230
rect 6924 -250 7000 -201
rect 9000 3424 13000 3500
rect 9000 3319 9261 3424
rect 9000 3201 9073 3319
rect 9191 3306 9261 3319
rect 9379 3306 9421 3424
rect 9539 3306 9581 3424
rect 9699 3306 9741 3424
rect 9859 3306 9901 3424
rect 10019 3306 10061 3424
rect 10179 3306 10221 3424
rect 10339 3306 10381 3424
rect 10499 3306 10541 3424
rect 10659 3306 10701 3424
rect 10819 3306 10861 3424
rect 10979 3306 11021 3424
rect 11139 3306 11181 3424
rect 11299 3306 11341 3424
rect 11459 3306 11501 3424
rect 11619 3306 11661 3424
rect 11779 3306 11821 3424
rect 11939 3306 11981 3424
rect 12099 3306 12141 3424
rect 12259 3306 12301 3424
rect 12419 3306 12461 3424
rect 12579 3306 12621 3424
rect 12739 3319 13000 3424
rect 12739 3306 12806 3319
rect 9191 3230 12806 3306
rect 9191 3201 9270 3230
rect 9000 3159 9270 3201
rect 9000 3041 9073 3159
rect 9191 3041 9270 3159
rect 9000 2999 9270 3041
rect 9000 2881 9073 2999
rect 9191 2881 9270 2999
rect 9000 2839 9270 2881
rect 9000 2721 9073 2839
rect 9191 2721 9270 2839
rect 9000 2679 9270 2721
rect 9000 2561 9073 2679
rect 9191 2561 9270 2679
rect 9000 2519 9270 2561
rect 9000 2401 9073 2519
rect 9191 2401 9270 2519
rect 9000 2359 9270 2401
rect 9000 2241 9073 2359
rect 9191 2241 9270 2359
rect 9000 2199 9270 2241
rect 9000 2081 9073 2199
rect 9191 2081 9270 2199
rect 9000 2039 9270 2081
rect 9000 1921 9073 2039
rect 9191 1921 9270 2039
rect 9000 1879 9270 1921
rect 9000 1761 9073 1879
rect 9191 1761 9270 1879
rect 9000 1719 9270 1761
rect 9000 1601 9073 1719
rect 9191 1601 9270 1719
rect 9000 1559 9270 1601
rect 9000 1441 9073 1559
rect 9191 1441 9270 1559
rect 9000 1399 9270 1441
rect 9000 1281 9073 1399
rect 9191 1281 9270 1399
rect 9000 1239 9270 1281
rect 9000 1121 9073 1239
rect 9191 1121 9270 1239
rect 9000 1079 9270 1121
rect 9000 961 9073 1079
rect 9191 961 9270 1079
rect 9000 919 9270 961
rect 9000 801 9073 919
rect 9191 801 9270 919
rect 9000 759 9270 801
rect 9000 641 9073 759
rect 9191 641 9270 759
rect 9000 599 9270 641
rect 9000 481 9073 599
rect 9191 481 9270 599
rect 9000 439 9270 481
rect 9000 321 9073 439
rect 9191 321 9270 439
rect 9000 279 9270 321
rect 9000 161 9073 279
rect 9191 161 9270 279
rect 9000 119 9270 161
rect 9000 1 9073 119
rect 9191 1 9270 119
rect 9000 -41 9270 1
rect 9000 -159 9073 -41
rect 9191 -159 9270 -41
rect 9000 -201 9270 -159
rect 3191 -319 3261 -304
rect 3000 -422 3261 -319
rect 3379 -422 3421 -304
rect 3539 -422 3581 -304
rect 3699 -422 3741 -304
rect 3859 -422 3901 -304
rect 4019 -422 4061 -304
rect 4179 -422 4221 -304
rect 4339 -422 4381 -304
rect 4499 -422 4541 -304
rect 4659 -422 4701 -304
rect 4819 -422 4861 -304
rect 4979 -422 5021 -304
rect 5139 -422 5181 -304
rect 5299 -422 5341 -304
rect 5459 -422 5501 -304
rect 5619 -422 5661 -304
rect 5779 -422 5821 -304
rect 5939 -422 5981 -304
rect 6099 -422 6141 -304
rect 6259 -422 6301 -304
rect 6419 -422 6461 -304
rect 6579 -422 6621 -304
rect 6739 -319 6806 -304
rect 6924 -319 8750 -250
rect 6739 -350 8750 -319
rect 6739 -422 7000 -350
rect 3000 -500 7000 -422
rect 8650 -550 8750 -350
rect 9000 -319 9073 -201
rect 9191 -230 9270 -201
rect 12730 3201 12806 3230
rect 12924 3201 13000 3319
rect 12730 3159 13000 3201
rect 12730 3041 12806 3159
rect 12924 3041 13000 3159
rect 12730 2999 13000 3041
rect 12730 2881 12806 2999
rect 12924 2881 13000 2999
rect 12730 2839 13000 2881
rect 12730 2721 12806 2839
rect 12924 2721 13000 2839
rect 12730 2679 13000 2721
rect 12730 2561 12806 2679
rect 12924 2561 13000 2679
rect 12730 2519 13000 2561
rect 12730 2401 12806 2519
rect 12924 2401 13000 2519
rect 12730 2359 13000 2401
rect 12730 2241 12806 2359
rect 12924 2241 13000 2359
rect 12730 2199 13000 2241
rect 12730 2081 12806 2199
rect 12924 2081 13000 2199
rect 12730 2039 13000 2081
rect 12730 1921 12806 2039
rect 12924 1921 13000 2039
rect 12730 1879 13000 1921
rect 12730 1761 12806 1879
rect 12924 1761 13000 1879
rect 12730 1719 13000 1761
rect 12730 1601 12806 1719
rect 12924 1601 13000 1719
rect 12730 1559 13000 1601
rect 12730 1441 12806 1559
rect 12924 1441 13000 1559
rect 12730 1399 13000 1441
rect 12730 1281 12806 1399
rect 12924 1281 13000 1399
rect 12730 1239 13000 1281
rect 12730 1121 12806 1239
rect 12924 1121 13000 1239
rect 12730 1079 13000 1121
rect 12730 961 12806 1079
rect 12924 961 13000 1079
rect 12730 919 13000 961
rect 12730 801 12806 919
rect 12924 801 13000 919
rect 12730 759 13000 801
rect 12730 641 12806 759
rect 12924 641 13000 759
rect 12730 599 13000 641
rect 12730 481 12806 599
rect 12924 481 13000 599
rect 12730 439 13000 481
rect 12730 321 12806 439
rect 12924 321 13000 439
rect 12730 279 13000 321
rect 12730 161 12806 279
rect 12924 161 13000 279
rect 12730 119 13000 161
rect 12730 1 12806 119
rect 12924 1 13000 119
rect 12730 -41 13000 1
rect 12730 -159 12806 -41
rect 12924 -159 13000 -41
rect 12730 -201 13000 -159
rect 12730 -230 12806 -201
rect 9191 -304 12806 -230
rect 9191 -319 9261 -304
rect 9000 -422 9261 -319
rect 9379 -422 9421 -304
rect 9539 -422 9581 -304
rect 9699 -422 9741 -304
rect 9859 -422 9901 -304
rect 10019 -422 10061 -304
rect 10179 -422 10221 -304
rect 10339 -422 10381 -304
rect 10499 -422 10541 -304
rect 10659 -422 10701 -304
rect 10819 -422 10861 -304
rect 10979 -422 11021 -304
rect 11139 -422 11181 -304
rect 11299 -422 11341 -304
rect 11459 -422 11501 -304
rect 11619 -422 11661 -304
rect 11779 -422 11821 -304
rect 11939 -422 11981 -304
rect 12099 -422 12141 -304
rect 12259 -422 12301 -304
rect 12419 -422 12461 -304
rect 12579 -422 12621 -304
rect 12739 -319 12806 -304
rect 12924 -319 13000 -201
rect 12739 -422 13000 -319
rect 9000 -500 13000 -422
rect 15000 3424 19000 3500
rect 15000 3319 15261 3424
rect 15000 3201 15073 3319
rect 15191 3306 15261 3319
rect 15379 3306 15421 3424
rect 15539 3306 15581 3424
rect 15699 3306 15741 3424
rect 15859 3306 15901 3424
rect 16019 3306 16061 3424
rect 16179 3306 16221 3424
rect 16339 3306 16381 3424
rect 16499 3306 16541 3424
rect 16659 3306 16701 3424
rect 16819 3306 16861 3424
rect 16979 3306 17021 3424
rect 17139 3306 17181 3424
rect 17299 3306 17341 3424
rect 17459 3306 17501 3424
rect 17619 3306 17661 3424
rect 17779 3306 17821 3424
rect 17939 3306 17981 3424
rect 18099 3306 18141 3424
rect 18259 3306 18301 3424
rect 18419 3306 18461 3424
rect 18579 3306 18621 3424
rect 18739 3319 19000 3424
rect 18739 3306 18806 3319
rect 15191 3230 18806 3306
rect 15191 3201 15270 3230
rect 15000 3159 15270 3201
rect 15000 3041 15073 3159
rect 15191 3041 15270 3159
rect 15000 2999 15270 3041
rect 15000 2881 15073 2999
rect 15191 2881 15270 2999
rect 15000 2839 15270 2881
rect 15000 2721 15073 2839
rect 15191 2721 15270 2839
rect 15000 2679 15270 2721
rect 15000 2561 15073 2679
rect 15191 2561 15270 2679
rect 15000 2519 15270 2561
rect 15000 2401 15073 2519
rect 15191 2401 15270 2519
rect 15000 2359 15270 2401
rect 15000 2241 15073 2359
rect 15191 2241 15270 2359
rect 15000 2199 15270 2241
rect 15000 2081 15073 2199
rect 15191 2081 15270 2199
rect 15000 2039 15270 2081
rect 15000 1921 15073 2039
rect 15191 1921 15270 2039
rect 15000 1879 15270 1921
rect 15000 1761 15073 1879
rect 15191 1761 15270 1879
rect 15000 1719 15270 1761
rect 15000 1601 15073 1719
rect 15191 1601 15270 1719
rect 15000 1559 15270 1601
rect 15000 1441 15073 1559
rect 15191 1441 15270 1559
rect 15000 1399 15270 1441
rect 15000 1281 15073 1399
rect 15191 1281 15270 1399
rect 15000 1239 15270 1281
rect 15000 1121 15073 1239
rect 15191 1121 15270 1239
rect 15000 1079 15270 1121
rect 15000 961 15073 1079
rect 15191 961 15270 1079
rect 15000 919 15270 961
rect 15000 801 15073 919
rect 15191 801 15270 919
rect 15000 759 15270 801
rect 15000 641 15073 759
rect 15191 641 15270 759
rect 15000 599 15270 641
rect 15000 481 15073 599
rect 15191 481 15270 599
rect 15000 439 15270 481
rect 15000 321 15073 439
rect 15191 321 15270 439
rect 15000 279 15270 321
rect 15000 161 15073 279
rect 15191 161 15270 279
rect 15000 119 15270 161
rect 15000 1 15073 119
rect 15191 1 15270 119
rect 15000 -41 15270 1
rect 15000 -159 15073 -41
rect 15191 -159 15270 -41
rect 15000 -201 15270 -159
rect 15000 -319 15073 -201
rect 15191 -230 15270 -201
rect 18730 3201 18806 3230
rect 18924 3201 19000 3319
rect 18730 3159 19000 3201
rect 18730 3041 18806 3159
rect 18924 3041 19000 3159
rect 18730 2999 19000 3041
rect 18730 2881 18806 2999
rect 18924 2881 19000 2999
rect 18730 2839 19000 2881
rect 18730 2721 18806 2839
rect 18924 2721 19000 2839
rect 18730 2679 19000 2721
rect 18730 2561 18806 2679
rect 18924 2561 19000 2679
rect 18730 2519 19000 2561
rect 18730 2401 18806 2519
rect 18924 2401 19000 2519
rect 18730 2359 19000 2401
rect 18730 2241 18806 2359
rect 18924 2241 19000 2359
rect 18730 2199 19000 2241
rect 18730 2081 18806 2199
rect 18924 2081 19000 2199
rect 18730 2039 19000 2081
rect 18730 1921 18806 2039
rect 18924 1921 19000 2039
rect 18730 1879 19000 1921
rect 18730 1761 18806 1879
rect 18924 1761 19000 1879
rect 18730 1719 19000 1761
rect 18730 1601 18806 1719
rect 18924 1601 19000 1719
rect 18730 1559 19000 1601
rect 18730 1441 18806 1559
rect 18924 1441 19000 1559
rect 18730 1399 19000 1441
rect 18730 1281 18806 1399
rect 18924 1281 19000 1399
rect 18730 1239 19000 1281
rect 18730 1121 18806 1239
rect 18924 1121 19000 1239
rect 18730 1079 19000 1121
rect 18730 961 18806 1079
rect 18924 961 19000 1079
rect 18730 919 19000 961
rect 18730 801 18806 919
rect 18924 801 19000 919
rect 18730 759 19000 801
rect 18730 641 18806 759
rect 18924 641 19000 759
rect 18730 599 19000 641
rect 18730 481 18806 599
rect 18924 481 19000 599
rect 18730 439 19000 481
rect 18730 321 18806 439
rect 18924 321 19000 439
rect 18730 279 19000 321
rect 18730 161 18806 279
rect 18924 161 19000 279
rect 18730 119 19000 161
rect 18730 1 18806 119
rect 18924 1 19000 119
rect 18730 -41 19000 1
rect 18730 -159 18806 -41
rect 18924 -159 19000 -41
rect 18730 -201 19000 -159
rect 18730 -230 18806 -201
rect 15191 -304 18806 -230
rect 15191 -319 15261 -304
rect 15000 -422 15261 -319
rect 15379 -422 15421 -304
rect 15539 -422 15581 -304
rect 15699 -422 15741 -304
rect 15859 -422 15901 -304
rect 16019 -422 16061 -304
rect 16179 -422 16221 -304
rect 16339 -422 16381 -304
rect 16499 -422 16541 -304
rect 16659 -422 16701 -304
rect 16819 -422 16861 -304
rect 16979 -422 17021 -304
rect 17139 -422 17181 -304
rect 17299 -422 17341 -304
rect 17459 -422 17501 -304
rect 17619 -422 17661 -304
rect 17779 -422 17821 -304
rect 17939 -422 17981 -304
rect 18099 -422 18141 -304
rect 18259 -422 18301 -304
rect 18419 -422 18461 -304
rect 18579 -422 18621 -304
rect 18739 -319 18806 -304
rect 18924 -319 19000 -201
rect 18739 -422 19000 -319
rect 15000 -500 19000 -422
rect 21000 3424 25000 3500
rect 21000 3319 21261 3424
rect 21000 3201 21073 3319
rect 21191 3306 21261 3319
rect 21379 3306 21421 3424
rect 21539 3306 21581 3424
rect 21699 3306 21741 3424
rect 21859 3306 21901 3424
rect 22019 3306 22061 3424
rect 22179 3306 22221 3424
rect 22339 3306 22381 3424
rect 22499 3306 22541 3424
rect 22659 3306 22701 3424
rect 22819 3306 22861 3424
rect 22979 3306 23021 3424
rect 23139 3306 23181 3424
rect 23299 3306 23341 3424
rect 23459 3306 23501 3424
rect 23619 3306 23661 3424
rect 23779 3306 23821 3424
rect 23939 3306 23981 3424
rect 24099 3306 24141 3424
rect 24259 3306 24301 3424
rect 24419 3306 24461 3424
rect 24579 3306 24621 3424
rect 24739 3319 25000 3424
rect 24739 3306 24806 3319
rect 21191 3230 24806 3306
rect 21191 3201 21270 3230
rect 21000 3159 21270 3201
rect 21000 3041 21073 3159
rect 21191 3041 21270 3159
rect 21000 2999 21270 3041
rect 21000 2881 21073 2999
rect 21191 2881 21270 2999
rect 21000 2839 21270 2881
rect 21000 2721 21073 2839
rect 21191 2721 21270 2839
rect 21000 2679 21270 2721
rect 21000 2561 21073 2679
rect 21191 2561 21270 2679
rect 21000 2519 21270 2561
rect 21000 2401 21073 2519
rect 21191 2401 21270 2519
rect 21000 2359 21270 2401
rect 21000 2241 21073 2359
rect 21191 2241 21270 2359
rect 21000 2199 21270 2241
rect 21000 2081 21073 2199
rect 21191 2081 21270 2199
rect 21000 2039 21270 2081
rect 21000 1921 21073 2039
rect 21191 1921 21270 2039
rect 21000 1879 21270 1921
rect 21000 1761 21073 1879
rect 21191 1761 21270 1879
rect 21000 1719 21270 1761
rect 21000 1601 21073 1719
rect 21191 1601 21270 1719
rect 21000 1559 21270 1601
rect 21000 1441 21073 1559
rect 21191 1441 21270 1559
rect 21000 1399 21270 1441
rect 21000 1281 21073 1399
rect 21191 1281 21270 1399
rect 21000 1239 21270 1281
rect 21000 1121 21073 1239
rect 21191 1121 21270 1239
rect 21000 1079 21270 1121
rect 21000 961 21073 1079
rect 21191 961 21270 1079
rect 21000 919 21270 961
rect 21000 801 21073 919
rect 21191 801 21270 919
rect 21000 759 21270 801
rect 21000 641 21073 759
rect 21191 641 21270 759
rect 21000 599 21270 641
rect 21000 481 21073 599
rect 21191 481 21270 599
rect 21000 439 21270 481
rect 21000 321 21073 439
rect 21191 321 21270 439
rect 21000 279 21270 321
rect 21000 161 21073 279
rect 21191 161 21270 279
rect 21000 119 21270 161
rect 21000 1 21073 119
rect 21191 1 21270 119
rect 21000 -41 21270 1
rect 21000 -159 21073 -41
rect 21191 -159 21270 -41
rect 21000 -201 21270 -159
rect 21000 -319 21073 -201
rect 21191 -230 21270 -201
rect 24730 3201 24806 3230
rect 24924 3201 25000 3319
rect 24730 3159 25000 3201
rect 24730 3041 24806 3159
rect 24924 3041 25000 3159
rect 24730 2999 25000 3041
rect 24730 2881 24806 2999
rect 24924 2881 25000 2999
rect 24730 2839 25000 2881
rect 24730 2721 24806 2839
rect 24924 2721 25000 2839
rect 24730 2679 25000 2721
rect 24730 2561 24806 2679
rect 24924 2561 25000 2679
rect 24730 2519 25000 2561
rect 24730 2401 24806 2519
rect 24924 2401 25000 2519
rect 24730 2359 25000 2401
rect 24730 2241 24806 2359
rect 24924 2241 25000 2359
rect 24730 2199 25000 2241
rect 24730 2081 24806 2199
rect 24924 2081 25000 2199
rect 24730 2039 25000 2081
rect 24730 1921 24806 2039
rect 24924 1921 25000 2039
rect 24730 1879 25000 1921
rect 24730 1761 24806 1879
rect 24924 1761 25000 1879
rect 24730 1719 25000 1761
rect 24730 1601 24806 1719
rect 24924 1601 25000 1719
rect 24730 1559 25000 1601
rect 24730 1441 24806 1559
rect 24924 1441 25000 1559
rect 24730 1399 25000 1441
rect 24730 1281 24806 1399
rect 24924 1281 25000 1399
rect 24730 1239 25000 1281
rect 24730 1121 24806 1239
rect 24924 1121 25000 1239
rect 24730 1079 25000 1121
rect 24730 961 24806 1079
rect 24924 961 25000 1079
rect 24730 919 25000 961
rect 24730 801 24806 919
rect 24924 801 25000 919
rect 24730 759 25000 801
rect 24730 641 24806 759
rect 24924 641 25000 759
rect 24730 599 25000 641
rect 24730 481 24806 599
rect 24924 481 25000 599
rect 24730 439 25000 481
rect 24730 321 24806 439
rect 24924 321 25000 439
rect 24730 279 25000 321
rect 24730 161 24806 279
rect 24924 161 25000 279
rect 24730 119 25000 161
rect 24730 1 24806 119
rect 24924 1 25000 119
rect 24730 -41 25000 1
rect 24730 -159 24806 -41
rect 24924 -159 25000 -41
rect 24730 -201 25000 -159
rect 24730 -230 24806 -201
rect 21191 -304 24806 -230
rect 21191 -319 21261 -304
rect 21000 -422 21261 -319
rect 21379 -422 21421 -304
rect 21539 -422 21581 -304
rect 21699 -422 21741 -304
rect 21859 -422 21901 -304
rect 22019 -422 22061 -304
rect 22179 -422 22221 -304
rect 22339 -422 22381 -304
rect 22499 -422 22541 -304
rect 22659 -422 22701 -304
rect 22819 -422 22861 -304
rect 22979 -422 23021 -304
rect 23139 -422 23181 -304
rect 23299 -422 23341 -304
rect 23459 -422 23501 -304
rect 23619 -422 23661 -304
rect 23779 -422 23821 -304
rect 23939 -422 23981 -304
rect 24099 -422 24141 -304
rect 24259 -422 24301 -304
rect 24419 -422 24461 -304
rect 24579 -422 24621 -304
rect 24739 -319 24806 -304
rect 24924 -319 25000 -201
rect 24739 -422 25000 -319
rect 21000 -500 25000 -422
rect 8650 -650 14550 -550
rect 14450 -750 14550 -650
rect 14450 -850 15650 -750
rect 16900 -850 19000 -500
rect 11750 -2770 12450 -2750
rect 11065 -2800 12450 -2770
rect 11750 -2850 12450 -2800
rect 5500 -4550 6600 -3950
rect 5500 -5500 6150 -4550
rect 12350 -5150 12450 -2850
rect 15550 -3200 15650 -850
rect 21850 -1450 22500 -500
rect 21400 -2050 22500 -1450
rect 15550 -3250 15750 -3200
rect 9000 -5500 11100 -5150
rect 12350 -5250 13550 -5150
rect 13450 -5350 13550 -5250
rect 13450 -5450 19350 -5350
rect 3000 -5578 7000 -5500
rect 3000 -5681 3261 -5578
rect 3000 -5799 3076 -5681
rect 3194 -5696 3261 -5681
rect 3379 -5696 3421 -5578
rect 3539 -5696 3581 -5578
rect 3699 -5696 3741 -5578
rect 3859 -5696 3901 -5578
rect 4019 -5696 4061 -5578
rect 4179 -5696 4221 -5578
rect 4339 -5696 4381 -5578
rect 4499 -5696 4541 -5578
rect 4659 -5696 4701 -5578
rect 4819 -5696 4861 -5578
rect 4979 -5696 5021 -5578
rect 5139 -5696 5181 -5578
rect 5299 -5696 5341 -5578
rect 5459 -5696 5501 -5578
rect 5619 -5696 5661 -5578
rect 5779 -5696 5821 -5578
rect 5939 -5696 5981 -5578
rect 6099 -5696 6141 -5578
rect 6259 -5696 6301 -5578
rect 6419 -5696 6461 -5578
rect 6579 -5696 6621 -5578
rect 6739 -5681 7000 -5578
rect 6739 -5696 6809 -5681
rect 3194 -5770 6809 -5696
rect 3194 -5799 3270 -5770
rect 3000 -5841 3270 -5799
rect 3000 -5959 3076 -5841
rect 3194 -5959 3270 -5841
rect 3000 -6001 3270 -5959
rect 3000 -6119 3076 -6001
rect 3194 -6119 3270 -6001
rect 3000 -6161 3270 -6119
rect 3000 -6279 3076 -6161
rect 3194 -6279 3270 -6161
rect 3000 -6321 3270 -6279
rect 3000 -6439 3076 -6321
rect 3194 -6439 3270 -6321
rect 3000 -6481 3270 -6439
rect 3000 -6599 3076 -6481
rect 3194 -6599 3270 -6481
rect 3000 -6641 3270 -6599
rect 3000 -6759 3076 -6641
rect 3194 -6759 3270 -6641
rect 3000 -6801 3270 -6759
rect 3000 -6919 3076 -6801
rect 3194 -6919 3270 -6801
rect 3000 -6961 3270 -6919
rect 3000 -7079 3076 -6961
rect 3194 -7079 3270 -6961
rect 3000 -7121 3270 -7079
rect 3000 -7239 3076 -7121
rect 3194 -7239 3270 -7121
rect 3000 -7281 3270 -7239
rect 3000 -7399 3076 -7281
rect 3194 -7399 3270 -7281
rect 3000 -7441 3270 -7399
rect 3000 -7559 3076 -7441
rect 3194 -7559 3270 -7441
rect 3000 -7601 3270 -7559
rect 3000 -7719 3076 -7601
rect 3194 -7719 3270 -7601
rect 3000 -7761 3270 -7719
rect 3000 -7879 3076 -7761
rect 3194 -7879 3270 -7761
rect 3000 -7921 3270 -7879
rect 3000 -8039 3076 -7921
rect 3194 -8039 3270 -7921
rect 3000 -8081 3270 -8039
rect 3000 -8199 3076 -8081
rect 3194 -8199 3270 -8081
rect 3000 -8241 3270 -8199
rect 3000 -8359 3076 -8241
rect 3194 -8359 3270 -8241
rect 3000 -8401 3270 -8359
rect 3000 -8519 3076 -8401
rect 3194 -8519 3270 -8401
rect 3000 -8561 3270 -8519
rect 3000 -8679 3076 -8561
rect 3194 -8679 3270 -8561
rect 3000 -8721 3270 -8679
rect 3000 -8839 3076 -8721
rect 3194 -8839 3270 -8721
rect 3000 -8881 3270 -8839
rect 3000 -8999 3076 -8881
rect 3194 -8999 3270 -8881
rect 3000 -9041 3270 -8999
rect 3000 -9159 3076 -9041
rect 3194 -9159 3270 -9041
rect 3000 -9201 3270 -9159
rect 3000 -9319 3076 -9201
rect 3194 -9230 3270 -9201
rect 6730 -5799 6809 -5770
rect 6927 -5799 7000 -5681
rect 6730 -5841 7000 -5799
rect 6730 -5959 6809 -5841
rect 6927 -5959 7000 -5841
rect 6730 -6001 7000 -5959
rect 6730 -6119 6809 -6001
rect 6927 -6119 7000 -6001
rect 6730 -6161 7000 -6119
rect 6730 -6279 6809 -6161
rect 6927 -6279 7000 -6161
rect 6730 -6321 7000 -6279
rect 6730 -6439 6809 -6321
rect 6927 -6439 7000 -6321
rect 6730 -6481 7000 -6439
rect 6730 -6599 6809 -6481
rect 6927 -6599 7000 -6481
rect 6730 -6641 7000 -6599
rect 6730 -6759 6809 -6641
rect 6927 -6759 7000 -6641
rect 6730 -6801 7000 -6759
rect 6730 -6919 6809 -6801
rect 6927 -6919 7000 -6801
rect 6730 -6961 7000 -6919
rect 6730 -7079 6809 -6961
rect 6927 -7079 7000 -6961
rect 6730 -7121 7000 -7079
rect 6730 -7239 6809 -7121
rect 6927 -7239 7000 -7121
rect 6730 -7281 7000 -7239
rect 6730 -7399 6809 -7281
rect 6927 -7399 7000 -7281
rect 6730 -7441 7000 -7399
rect 6730 -7559 6809 -7441
rect 6927 -7559 7000 -7441
rect 6730 -7601 7000 -7559
rect 6730 -7719 6809 -7601
rect 6927 -7719 7000 -7601
rect 6730 -7761 7000 -7719
rect 6730 -7879 6809 -7761
rect 6927 -7879 7000 -7761
rect 6730 -7921 7000 -7879
rect 6730 -8039 6809 -7921
rect 6927 -8039 7000 -7921
rect 6730 -8081 7000 -8039
rect 6730 -8199 6809 -8081
rect 6927 -8199 7000 -8081
rect 6730 -8241 7000 -8199
rect 6730 -8359 6809 -8241
rect 6927 -8359 7000 -8241
rect 6730 -8401 7000 -8359
rect 6730 -8519 6809 -8401
rect 6927 -8519 7000 -8401
rect 6730 -8561 7000 -8519
rect 6730 -8679 6809 -8561
rect 6927 -8679 7000 -8561
rect 6730 -8721 7000 -8679
rect 6730 -8839 6809 -8721
rect 6927 -8839 7000 -8721
rect 6730 -8881 7000 -8839
rect 6730 -8999 6809 -8881
rect 6927 -8999 7000 -8881
rect 6730 -9041 7000 -8999
rect 6730 -9159 6809 -9041
rect 6927 -9159 7000 -9041
rect 6730 -9201 7000 -9159
rect 6730 -9230 6809 -9201
rect 3194 -9306 6809 -9230
rect 3194 -9319 3261 -9306
rect 3000 -9424 3261 -9319
rect 3379 -9424 3421 -9306
rect 3539 -9424 3581 -9306
rect 3699 -9424 3741 -9306
rect 3859 -9424 3901 -9306
rect 4019 -9424 4061 -9306
rect 4179 -9424 4221 -9306
rect 4339 -9424 4381 -9306
rect 4499 -9424 4541 -9306
rect 4659 -9424 4701 -9306
rect 4819 -9424 4861 -9306
rect 4979 -9424 5021 -9306
rect 5139 -9424 5181 -9306
rect 5299 -9424 5341 -9306
rect 5459 -9424 5501 -9306
rect 5619 -9424 5661 -9306
rect 5779 -9424 5821 -9306
rect 5939 -9424 5981 -9306
rect 6099 -9424 6141 -9306
rect 6259 -9424 6301 -9306
rect 6419 -9424 6461 -9306
rect 6579 -9424 6621 -9306
rect 6739 -9319 6809 -9306
rect 6927 -9319 7000 -9201
rect 6739 -9424 7000 -9319
rect 3000 -9500 7000 -9424
rect 9000 -5578 13000 -5500
rect 9000 -5681 9261 -5578
rect 9000 -5799 9076 -5681
rect 9194 -5696 9261 -5681
rect 9379 -5696 9421 -5578
rect 9539 -5696 9581 -5578
rect 9699 -5696 9741 -5578
rect 9859 -5696 9901 -5578
rect 10019 -5696 10061 -5578
rect 10179 -5696 10221 -5578
rect 10339 -5696 10381 -5578
rect 10499 -5696 10541 -5578
rect 10659 -5696 10701 -5578
rect 10819 -5696 10861 -5578
rect 10979 -5696 11021 -5578
rect 11139 -5696 11181 -5578
rect 11299 -5696 11341 -5578
rect 11459 -5696 11501 -5578
rect 11619 -5696 11661 -5578
rect 11779 -5696 11821 -5578
rect 11939 -5696 11981 -5578
rect 12099 -5696 12141 -5578
rect 12259 -5696 12301 -5578
rect 12419 -5696 12461 -5578
rect 12579 -5696 12621 -5578
rect 12739 -5681 13000 -5578
rect 12739 -5696 12809 -5681
rect 9194 -5770 12809 -5696
rect 9194 -5799 9270 -5770
rect 9000 -5841 9270 -5799
rect 9000 -5959 9076 -5841
rect 9194 -5959 9270 -5841
rect 9000 -6001 9270 -5959
rect 9000 -6119 9076 -6001
rect 9194 -6119 9270 -6001
rect 9000 -6161 9270 -6119
rect 9000 -6279 9076 -6161
rect 9194 -6279 9270 -6161
rect 9000 -6321 9270 -6279
rect 9000 -6439 9076 -6321
rect 9194 -6439 9270 -6321
rect 9000 -6481 9270 -6439
rect 9000 -6599 9076 -6481
rect 9194 -6599 9270 -6481
rect 9000 -6641 9270 -6599
rect 9000 -6759 9076 -6641
rect 9194 -6759 9270 -6641
rect 9000 -6801 9270 -6759
rect 9000 -6919 9076 -6801
rect 9194 -6919 9270 -6801
rect 9000 -6961 9270 -6919
rect 9000 -7079 9076 -6961
rect 9194 -7079 9270 -6961
rect 9000 -7121 9270 -7079
rect 9000 -7239 9076 -7121
rect 9194 -7239 9270 -7121
rect 9000 -7281 9270 -7239
rect 9000 -7399 9076 -7281
rect 9194 -7399 9270 -7281
rect 9000 -7441 9270 -7399
rect 9000 -7559 9076 -7441
rect 9194 -7559 9270 -7441
rect 9000 -7601 9270 -7559
rect 9000 -7719 9076 -7601
rect 9194 -7719 9270 -7601
rect 9000 -7761 9270 -7719
rect 9000 -7879 9076 -7761
rect 9194 -7879 9270 -7761
rect 9000 -7921 9270 -7879
rect 9000 -8039 9076 -7921
rect 9194 -8039 9270 -7921
rect 9000 -8081 9270 -8039
rect 9000 -8199 9076 -8081
rect 9194 -8199 9270 -8081
rect 9000 -8241 9270 -8199
rect 9000 -8359 9076 -8241
rect 9194 -8359 9270 -8241
rect 9000 -8401 9270 -8359
rect 9000 -8519 9076 -8401
rect 9194 -8519 9270 -8401
rect 9000 -8561 9270 -8519
rect 9000 -8679 9076 -8561
rect 9194 -8679 9270 -8561
rect 9000 -8721 9270 -8679
rect 9000 -8839 9076 -8721
rect 9194 -8839 9270 -8721
rect 9000 -8881 9270 -8839
rect 9000 -8999 9076 -8881
rect 9194 -8999 9270 -8881
rect 9000 -9041 9270 -8999
rect 9000 -9159 9076 -9041
rect 9194 -9159 9270 -9041
rect 9000 -9201 9270 -9159
rect 9000 -9319 9076 -9201
rect 9194 -9230 9270 -9201
rect 12730 -5799 12809 -5770
rect 12927 -5799 13000 -5681
rect 12730 -5841 13000 -5799
rect 12730 -5959 12809 -5841
rect 12927 -5959 13000 -5841
rect 12730 -6001 13000 -5959
rect 12730 -6119 12809 -6001
rect 12927 -6119 13000 -6001
rect 12730 -6161 13000 -6119
rect 12730 -6279 12809 -6161
rect 12927 -6279 13000 -6161
rect 12730 -6321 13000 -6279
rect 12730 -6439 12809 -6321
rect 12927 -6439 13000 -6321
rect 12730 -6481 13000 -6439
rect 12730 -6599 12809 -6481
rect 12927 -6599 13000 -6481
rect 12730 -6641 13000 -6599
rect 12730 -6759 12809 -6641
rect 12927 -6759 13000 -6641
rect 12730 -6801 13000 -6759
rect 12730 -6919 12809 -6801
rect 12927 -6919 13000 -6801
rect 12730 -6961 13000 -6919
rect 12730 -7079 12809 -6961
rect 12927 -7079 13000 -6961
rect 12730 -7121 13000 -7079
rect 12730 -7239 12809 -7121
rect 12927 -7239 13000 -7121
rect 12730 -7281 13000 -7239
rect 12730 -7399 12809 -7281
rect 12927 -7399 13000 -7281
rect 12730 -7441 13000 -7399
rect 12730 -7559 12809 -7441
rect 12927 -7559 13000 -7441
rect 12730 -7601 13000 -7559
rect 12730 -7719 12809 -7601
rect 12927 -7719 13000 -7601
rect 12730 -7761 13000 -7719
rect 12730 -7879 12809 -7761
rect 12927 -7879 13000 -7761
rect 12730 -7921 13000 -7879
rect 12730 -8039 12809 -7921
rect 12927 -8039 13000 -7921
rect 12730 -8081 13000 -8039
rect 12730 -8199 12809 -8081
rect 12927 -8199 13000 -8081
rect 12730 -8241 13000 -8199
rect 12730 -8359 12809 -8241
rect 12927 -8359 13000 -8241
rect 12730 -8401 13000 -8359
rect 12730 -8519 12809 -8401
rect 12927 -8519 13000 -8401
rect 12730 -8561 13000 -8519
rect 12730 -8679 12809 -8561
rect 12927 -8679 13000 -8561
rect 12730 -8721 13000 -8679
rect 12730 -8839 12809 -8721
rect 12927 -8839 13000 -8721
rect 12730 -8881 13000 -8839
rect 12730 -8999 12809 -8881
rect 12927 -8999 13000 -8881
rect 12730 -9041 13000 -8999
rect 12730 -9159 12809 -9041
rect 12927 -9159 13000 -9041
rect 12730 -9201 13000 -9159
rect 12730 -9230 12809 -9201
rect 9194 -9306 12809 -9230
rect 9194 -9319 9261 -9306
rect 9000 -9424 9261 -9319
rect 9379 -9424 9421 -9306
rect 9539 -9424 9581 -9306
rect 9699 -9424 9741 -9306
rect 9859 -9424 9901 -9306
rect 10019 -9424 10061 -9306
rect 10179 -9424 10221 -9306
rect 10339 -9424 10381 -9306
rect 10499 -9424 10541 -9306
rect 10659 -9424 10701 -9306
rect 10819 -9424 10861 -9306
rect 10979 -9424 11021 -9306
rect 11139 -9424 11181 -9306
rect 11299 -9424 11341 -9306
rect 11459 -9424 11501 -9306
rect 11619 -9424 11661 -9306
rect 11779 -9424 11821 -9306
rect 11939 -9424 11981 -9306
rect 12099 -9424 12141 -9306
rect 12259 -9424 12301 -9306
rect 12419 -9424 12461 -9306
rect 12579 -9424 12621 -9306
rect 12739 -9319 12809 -9306
rect 12927 -9319 13000 -9201
rect 12739 -9424 13000 -9319
rect 9000 -9500 13000 -9424
rect 15000 -5578 19000 -5500
rect 15000 -5681 15261 -5578
rect 15000 -5799 15076 -5681
rect 15194 -5696 15261 -5681
rect 15379 -5696 15421 -5578
rect 15539 -5696 15581 -5578
rect 15699 -5696 15741 -5578
rect 15859 -5696 15901 -5578
rect 16019 -5696 16061 -5578
rect 16179 -5696 16221 -5578
rect 16339 -5696 16381 -5578
rect 16499 -5696 16541 -5578
rect 16659 -5696 16701 -5578
rect 16819 -5696 16861 -5578
rect 16979 -5696 17021 -5578
rect 17139 -5696 17181 -5578
rect 17299 -5696 17341 -5578
rect 17459 -5696 17501 -5578
rect 17619 -5696 17661 -5578
rect 17779 -5696 17821 -5578
rect 17939 -5696 17981 -5578
rect 18099 -5696 18141 -5578
rect 18259 -5696 18301 -5578
rect 18419 -5696 18461 -5578
rect 18579 -5696 18621 -5578
rect 18739 -5681 19000 -5578
rect 18739 -5696 18809 -5681
rect 15194 -5770 18809 -5696
rect 15194 -5799 15270 -5770
rect 15000 -5841 15270 -5799
rect 15000 -5959 15076 -5841
rect 15194 -5959 15270 -5841
rect 15000 -6001 15270 -5959
rect 15000 -6119 15076 -6001
rect 15194 -6119 15270 -6001
rect 15000 -6161 15270 -6119
rect 15000 -6279 15076 -6161
rect 15194 -6279 15270 -6161
rect 15000 -6321 15270 -6279
rect 15000 -6439 15076 -6321
rect 15194 -6439 15270 -6321
rect 15000 -6481 15270 -6439
rect 15000 -6599 15076 -6481
rect 15194 -6599 15270 -6481
rect 15000 -6641 15270 -6599
rect 15000 -6759 15076 -6641
rect 15194 -6759 15270 -6641
rect 15000 -6801 15270 -6759
rect 15000 -6919 15076 -6801
rect 15194 -6919 15270 -6801
rect 15000 -6961 15270 -6919
rect 15000 -7079 15076 -6961
rect 15194 -7079 15270 -6961
rect 15000 -7121 15270 -7079
rect 15000 -7239 15076 -7121
rect 15194 -7239 15270 -7121
rect 15000 -7281 15270 -7239
rect 15000 -7399 15076 -7281
rect 15194 -7399 15270 -7281
rect 15000 -7441 15270 -7399
rect 15000 -7559 15076 -7441
rect 15194 -7559 15270 -7441
rect 15000 -7601 15270 -7559
rect 15000 -7719 15076 -7601
rect 15194 -7719 15270 -7601
rect 15000 -7761 15270 -7719
rect 15000 -7879 15076 -7761
rect 15194 -7879 15270 -7761
rect 15000 -7921 15270 -7879
rect 15000 -8039 15076 -7921
rect 15194 -8039 15270 -7921
rect 15000 -8081 15270 -8039
rect 15000 -8199 15076 -8081
rect 15194 -8199 15270 -8081
rect 15000 -8241 15270 -8199
rect 15000 -8359 15076 -8241
rect 15194 -8359 15270 -8241
rect 15000 -8401 15270 -8359
rect 15000 -8519 15076 -8401
rect 15194 -8519 15270 -8401
rect 15000 -8561 15270 -8519
rect 15000 -8679 15076 -8561
rect 15194 -8679 15270 -8561
rect 15000 -8721 15270 -8679
rect 15000 -8839 15076 -8721
rect 15194 -8839 15270 -8721
rect 15000 -8881 15270 -8839
rect 15000 -8999 15076 -8881
rect 15194 -8999 15270 -8881
rect 15000 -9041 15270 -8999
rect 15000 -9159 15076 -9041
rect 15194 -9159 15270 -9041
rect 15000 -9201 15270 -9159
rect 15000 -9319 15076 -9201
rect 15194 -9230 15270 -9201
rect 18730 -5799 18809 -5770
rect 18927 -5799 19000 -5681
rect 19250 -5650 19350 -5450
rect 21000 -5578 25000 -5500
rect 21000 -5650 21261 -5578
rect 19250 -5681 21261 -5650
rect 19250 -5750 21076 -5681
rect 21194 -5696 21261 -5681
rect 21379 -5696 21421 -5578
rect 21539 -5696 21581 -5578
rect 21699 -5696 21741 -5578
rect 21859 -5696 21901 -5578
rect 22019 -5696 22061 -5578
rect 22179 -5696 22221 -5578
rect 22339 -5696 22381 -5578
rect 22499 -5696 22541 -5578
rect 22659 -5696 22701 -5578
rect 22819 -5696 22861 -5578
rect 22979 -5696 23021 -5578
rect 23139 -5696 23181 -5578
rect 23299 -5696 23341 -5578
rect 23459 -5696 23501 -5578
rect 23619 -5696 23661 -5578
rect 23779 -5696 23821 -5578
rect 23939 -5696 23981 -5578
rect 24099 -5696 24141 -5578
rect 24259 -5696 24301 -5578
rect 24419 -5696 24461 -5578
rect 24579 -5696 24621 -5578
rect 24739 -5681 25000 -5578
rect 24739 -5696 24809 -5681
rect 18730 -5841 19000 -5799
rect 18730 -5959 18809 -5841
rect 18927 -5959 19000 -5841
rect 18730 -6001 19000 -5959
rect 18730 -6119 18809 -6001
rect 18927 -6119 19000 -6001
rect 18730 -6161 19000 -6119
rect 18730 -6279 18809 -6161
rect 18927 -6279 19000 -6161
rect 18730 -6321 19000 -6279
rect 18730 -6439 18809 -6321
rect 18927 -6439 19000 -6321
rect 18730 -6481 19000 -6439
rect 18730 -6599 18809 -6481
rect 18927 -6599 19000 -6481
rect 18730 -6641 19000 -6599
rect 18730 -6759 18809 -6641
rect 18927 -6759 19000 -6641
rect 18730 -6801 19000 -6759
rect 18730 -6919 18809 -6801
rect 18927 -6919 19000 -6801
rect 18730 -6961 19000 -6919
rect 18730 -7079 18809 -6961
rect 18927 -7079 19000 -6961
rect 18730 -7121 19000 -7079
rect 18730 -7239 18809 -7121
rect 18927 -7239 19000 -7121
rect 18730 -7281 19000 -7239
rect 18730 -7399 18809 -7281
rect 18927 -7399 19000 -7281
rect 18730 -7441 19000 -7399
rect 18730 -7559 18809 -7441
rect 18927 -7559 19000 -7441
rect 18730 -7601 19000 -7559
rect 18730 -7719 18809 -7601
rect 18927 -7719 19000 -7601
rect 18730 -7761 19000 -7719
rect 18730 -7879 18809 -7761
rect 18927 -7879 19000 -7761
rect 18730 -7921 19000 -7879
rect 18730 -8039 18809 -7921
rect 18927 -8039 19000 -7921
rect 18730 -8081 19000 -8039
rect 18730 -8199 18809 -8081
rect 18927 -8199 19000 -8081
rect 18730 -8241 19000 -8199
rect 18730 -8359 18809 -8241
rect 18927 -8359 19000 -8241
rect 18730 -8401 19000 -8359
rect 18730 -8519 18809 -8401
rect 18927 -8519 19000 -8401
rect 18730 -8561 19000 -8519
rect 18730 -8679 18809 -8561
rect 18927 -8679 19000 -8561
rect 18730 -8721 19000 -8679
rect 18730 -8839 18809 -8721
rect 18927 -8839 19000 -8721
rect 18730 -8881 19000 -8839
rect 18730 -8999 18809 -8881
rect 18927 -8999 19000 -8881
rect 18730 -9041 19000 -8999
rect 18730 -9159 18809 -9041
rect 18927 -9159 19000 -9041
rect 18730 -9201 19000 -9159
rect 18730 -9230 18809 -9201
rect 15194 -9306 18809 -9230
rect 15194 -9319 15261 -9306
rect 15000 -9424 15261 -9319
rect 15379 -9424 15421 -9306
rect 15539 -9424 15581 -9306
rect 15699 -9424 15741 -9306
rect 15859 -9424 15901 -9306
rect 16019 -9424 16061 -9306
rect 16179 -9424 16221 -9306
rect 16339 -9424 16381 -9306
rect 16499 -9424 16541 -9306
rect 16659 -9424 16701 -9306
rect 16819 -9424 16861 -9306
rect 16979 -9424 17021 -9306
rect 17139 -9424 17181 -9306
rect 17299 -9424 17341 -9306
rect 17459 -9424 17501 -9306
rect 17619 -9424 17661 -9306
rect 17779 -9424 17821 -9306
rect 17939 -9424 17981 -9306
rect 18099 -9424 18141 -9306
rect 18259 -9424 18301 -9306
rect 18419 -9424 18461 -9306
rect 18579 -9424 18621 -9306
rect 18739 -9319 18809 -9306
rect 18927 -9319 19000 -9201
rect 18739 -9424 19000 -9319
rect 15000 -9500 19000 -9424
rect 21000 -5799 21076 -5750
rect 21194 -5770 24809 -5696
rect 21194 -5799 21270 -5770
rect 21000 -5841 21270 -5799
rect 21000 -5959 21076 -5841
rect 21194 -5959 21270 -5841
rect 21000 -6001 21270 -5959
rect 21000 -6119 21076 -6001
rect 21194 -6119 21270 -6001
rect 21000 -6161 21270 -6119
rect 21000 -6279 21076 -6161
rect 21194 -6279 21270 -6161
rect 21000 -6321 21270 -6279
rect 21000 -6439 21076 -6321
rect 21194 -6439 21270 -6321
rect 21000 -6481 21270 -6439
rect 21000 -6599 21076 -6481
rect 21194 -6599 21270 -6481
rect 21000 -6641 21270 -6599
rect 21000 -6759 21076 -6641
rect 21194 -6759 21270 -6641
rect 21000 -6801 21270 -6759
rect 21000 -6919 21076 -6801
rect 21194 -6919 21270 -6801
rect 21000 -6961 21270 -6919
rect 21000 -7079 21076 -6961
rect 21194 -7079 21270 -6961
rect 21000 -7121 21270 -7079
rect 21000 -7239 21076 -7121
rect 21194 -7239 21270 -7121
rect 21000 -7281 21270 -7239
rect 21000 -7399 21076 -7281
rect 21194 -7399 21270 -7281
rect 21000 -7441 21270 -7399
rect 21000 -7559 21076 -7441
rect 21194 -7559 21270 -7441
rect 21000 -7601 21270 -7559
rect 21000 -7719 21076 -7601
rect 21194 -7719 21270 -7601
rect 21000 -7761 21270 -7719
rect 21000 -7879 21076 -7761
rect 21194 -7879 21270 -7761
rect 21000 -7921 21270 -7879
rect 21000 -8039 21076 -7921
rect 21194 -8039 21270 -7921
rect 21000 -8081 21270 -8039
rect 21000 -8199 21076 -8081
rect 21194 -8199 21270 -8081
rect 21000 -8241 21270 -8199
rect 21000 -8359 21076 -8241
rect 21194 -8359 21270 -8241
rect 21000 -8401 21270 -8359
rect 21000 -8519 21076 -8401
rect 21194 -8519 21270 -8401
rect 21000 -8561 21270 -8519
rect 21000 -8679 21076 -8561
rect 21194 -8679 21270 -8561
rect 21000 -8721 21270 -8679
rect 21000 -8839 21076 -8721
rect 21194 -8839 21270 -8721
rect 21000 -8881 21270 -8839
rect 21000 -8999 21076 -8881
rect 21194 -8999 21270 -8881
rect 21000 -9041 21270 -8999
rect 21000 -9159 21076 -9041
rect 21194 -9159 21270 -9041
rect 21000 -9201 21270 -9159
rect 21000 -9319 21076 -9201
rect 21194 -9230 21270 -9201
rect 24730 -5799 24809 -5770
rect 24927 -5799 25000 -5681
rect 24730 -5841 25000 -5799
rect 24730 -5959 24809 -5841
rect 24927 -5959 25000 -5841
rect 24730 -6001 25000 -5959
rect 24730 -6119 24809 -6001
rect 24927 -6119 25000 -6001
rect 24730 -6161 25000 -6119
rect 24730 -6279 24809 -6161
rect 24927 -6279 25000 -6161
rect 24730 -6321 25000 -6279
rect 24730 -6439 24809 -6321
rect 24927 -6439 25000 -6321
rect 24730 -6481 25000 -6439
rect 24730 -6599 24809 -6481
rect 24927 -6599 25000 -6481
rect 24730 -6641 25000 -6599
rect 24730 -6759 24809 -6641
rect 24927 -6759 25000 -6641
rect 24730 -6801 25000 -6759
rect 24730 -6919 24809 -6801
rect 24927 -6919 25000 -6801
rect 24730 -6961 25000 -6919
rect 24730 -7079 24809 -6961
rect 24927 -7079 25000 -6961
rect 24730 -7121 25000 -7079
rect 24730 -7239 24809 -7121
rect 24927 -7239 25000 -7121
rect 24730 -7281 25000 -7239
rect 24730 -7399 24809 -7281
rect 24927 -7399 25000 -7281
rect 24730 -7441 25000 -7399
rect 24730 -7559 24809 -7441
rect 24927 -7559 25000 -7441
rect 24730 -7601 25000 -7559
rect 24730 -7719 24809 -7601
rect 24927 -7719 25000 -7601
rect 24730 -7761 25000 -7719
rect 24730 -7879 24809 -7761
rect 24927 -7879 25000 -7761
rect 24730 -7921 25000 -7879
rect 24730 -8039 24809 -7921
rect 24927 -8039 25000 -7921
rect 24730 -8081 25000 -8039
rect 24730 -8199 24809 -8081
rect 24927 -8199 25000 -8081
rect 24730 -8241 25000 -8199
rect 24730 -8359 24809 -8241
rect 24927 -8359 25000 -8241
rect 24730 -8401 25000 -8359
rect 24730 -8519 24809 -8401
rect 24927 -8519 25000 -8401
rect 24730 -8561 25000 -8519
rect 24730 -8679 24809 -8561
rect 24927 -8679 25000 -8561
rect 24730 -8721 25000 -8679
rect 24730 -8839 24809 -8721
rect 24927 -8839 25000 -8721
rect 24730 -8881 25000 -8839
rect 24730 -8999 24809 -8881
rect 24927 -8999 25000 -8881
rect 24730 -9041 25000 -8999
rect 24730 -9159 24809 -9041
rect 24927 -9159 25000 -9041
rect 24730 -9201 25000 -9159
rect 24730 -9230 24809 -9201
rect 21194 -9306 24809 -9230
rect 21194 -9319 21261 -9306
rect 21000 -9424 21261 -9319
rect 21379 -9424 21421 -9306
rect 21539 -9424 21581 -9306
rect 21699 -9424 21741 -9306
rect 21859 -9424 21901 -9306
rect 22019 -9424 22061 -9306
rect 22179 -9424 22221 -9306
rect 22339 -9424 22381 -9306
rect 22499 -9424 22541 -9306
rect 22659 -9424 22701 -9306
rect 22819 -9424 22861 -9306
rect 22979 -9424 23021 -9306
rect 23139 -9424 23181 -9306
rect 23299 -9424 23341 -9306
rect 23459 -9424 23501 -9306
rect 23619 -9424 23661 -9306
rect 23779 -9424 23821 -9306
rect 23939 -9424 23981 -9306
rect 24099 -9424 24141 -9306
rect 24259 -9424 24301 -9306
rect 24419 -9424 24461 -9306
rect 24579 -9424 24621 -9306
rect 24739 -9319 24809 -9306
rect 24927 -9319 25000 -9201
rect 24739 -9424 25000 -9319
rect 21000 -9500 25000 -9424
rect 3050 -9800 3150 -9550
rect 3250 -9800 3350 -9550
rect 3050 -9850 3350 -9800
rect 3450 -9600 3700 -9550
rect 3850 -9600 4100 -9550
rect 3450 -9650 3750 -9600
rect 3450 -9850 3550 -9650
rect 3650 -9850 3750 -9650
rect 3100 -9900 3300 -9850
rect 3450 -9900 3750 -9850
rect 3850 -9650 4150 -9600
rect 3850 -9850 3950 -9650
rect 4050 -9850 4150 -9650
rect 9050 -9800 9150 -9550
rect 9250 -9800 9350 -9550
rect 9450 -9650 9750 -9550
rect 9850 -9650 10150 -9550
rect 9450 -9700 9550 -9650
rect 9850 -9700 9950 -9650
rect 9450 -9750 9700 -9700
rect 9850 -9750 10100 -9700
rect 9500 -9800 9750 -9750
rect 9900 -9800 10150 -9750
rect 9050 -9850 9350 -9800
rect 9650 -9850 9750 -9800
rect 10050 -9850 10150 -9800
rect 15050 -9800 15150 -9550
rect 15250 -9800 15350 -9550
rect 15450 -9650 15750 -9550
rect 15050 -9850 15350 -9800
rect 15550 -9850 15650 -9650
rect 15950 -9700 16050 -9600
rect 15850 -9800 16150 -9700
rect 21050 -9800 21150 -9550
rect 21250 -9800 21350 -9550
rect 21500 -9600 21700 -9550
rect 3850 -9900 4150 -9850
rect 9100 -9900 9300 -9850
rect 3150 -9950 3250 -9900
rect 3450 -9950 3700 -9900
rect 3850 -9950 4100 -9900
rect 9150 -9950 9250 -9900
rect 9450 -9950 9750 -9850
rect 9850 -9950 10150 -9850
rect 15100 -9900 15300 -9850
rect 15150 -9950 15250 -9900
rect 15450 -9950 15750 -9850
rect 15950 -9900 16050 -9800
rect 21050 -9850 21350 -9800
rect 21450 -9650 21750 -9600
rect 21450 -9850 21550 -9650
rect 21650 -9850 21750 -9650
rect 21950 -9700 22050 -9600
rect 21850 -9800 22150 -9700
rect 21100 -9900 21300 -9850
rect 21450 -9900 21750 -9850
rect 21950 -9900 22050 -9800
rect 21150 -9950 21250 -9900
rect 21500 -9950 21700 -9900
rect 9050 -11000 9350 -10950
rect 3050 -11150 3350 -11050
rect 9050 -11150 9350 -11050
rect 3050 -11200 3150 -11150
rect 9050 -11200 9150 -11150
rect 3050 -11250 3300 -11200
rect 9050 -11250 9300 -11200
rect 3100 -11300 3350 -11250
rect 9100 -11300 9350 -11250
rect 3250 -11350 3350 -11300
rect 9250 -11350 9350 -11300
rect 15050 -11300 15150 -11050
rect 15250 -11300 15350 -11050
rect 15050 -11350 15350 -11300
rect 15450 -11100 15700 -11050
rect 15450 -11150 15750 -11100
rect 15450 -11250 15550 -11150
rect 15650 -11250 15750 -11150
rect 15850 -11150 16150 -11050
rect 16250 -11150 16550 -11050
rect 15850 -11200 15950 -11150
rect 16250 -11200 16350 -11150
rect 15450 -11350 15700 -11250
rect 15850 -11300 16100 -11200
rect 16250 -11300 16500 -11200
rect 21050 -11300 21150 -11050
rect 21250 -11300 21350 -11050
rect 21450 -11150 21750 -11050
rect 15850 -11350 15950 -11300
rect 3050 -11450 3350 -11350
rect 9050 -11450 9350 -11350
rect 15100 -11400 15300 -11350
rect 15150 -11450 15250 -11400
rect 15450 -11450 15550 -11350
rect 15650 -11450 15750 -11350
rect 15850 -11450 16150 -11350
rect 16250 -11450 16350 -11300
rect 21050 -11350 21350 -11300
rect 21550 -11350 21650 -11150
rect 21850 -11300 22150 -11200
rect 21100 -11400 21300 -11350
rect 21150 -11450 21250 -11400
rect 21450 -11450 21750 -11350
rect 3000 -11578 7000 -11500
rect 3000 -11681 3261 -11578
rect 3000 -11799 3076 -11681
rect 3194 -11696 3261 -11681
rect 3379 -11696 3421 -11578
rect 3539 -11696 3581 -11578
rect 3699 -11696 3741 -11578
rect 3859 -11696 3901 -11578
rect 4019 -11696 4061 -11578
rect 4179 -11696 4221 -11578
rect 4339 -11696 4381 -11578
rect 4499 -11696 4541 -11578
rect 4659 -11696 4701 -11578
rect 4819 -11696 4861 -11578
rect 4979 -11696 5021 -11578
rect 5139 -11696 5181 -11578
rect 5299 -11696 5341 -11578
rect 5459 -11696 5501 -11578
rect 5619 -11696 5661 -11578
rect 5779 -11696 5821 -11578
rect 5939 -11696 5981 -11578
rect 6099 -11696 6141 -11578
rect 6259 -11696 6301 -11578
rect 6419 -11696 6461 -11578
rect 6579 -11696 6621 -11578
rect 6739 -11681 7000 -11578
rect 6739 -11696 6809 -11681
rect 3194 -11770 6809 -11696
rect 3194 -11799 3270 -11770
rect 3000 -11841 3270 -11799
rect 3000 -11959 3076 -11841
rect 3194 -11959 3270 -11841
rect 3000 -12001 3270 -11959
rect 3000 -12119 3076 -12001
rect 3194 -12119 3270 -12001
rect 3000 -12161 3270 -12119
rect 3000 -12279 3076 -12161
rect 3194 -12279 3270 -12161
rect 3000 -12321 3270 -12279
rect 3000 -12439 3076 -12321
rect 3194 -12439 3270 -12321
rect 3000 -12481 3270 -12439
rect 3000 -12599 3076 -12481
rect 3194 -12599 3270 -12481
rect 3000 -12641 3270 -12599
rect 3000 -12759 3076 -12641
rect 3194 -12759 3270 -12641
rect 3000 -12801 3270 -12759
rect 3000 -12919 3076 -12801
rect 3194 -12919 3270 -12801
rect 3000 -12961 3270 -12919
rect 3000 -13079 3076 -12961
rect 3194 -13079 3270 -12961
rect 3000 -13121 3270 -13079
rect 3000 -13239 3076 -13121
rect 3194 -13239 3270 -13121
rect 3000 -13281 3270 -13239
rect 3000 -13399 3076 -13281
rect 3194 -13399 3270 -13281
rect 3000 -13441 3270 -13399
rect 3000 -13559 3076 -13441
rect 3194 -13559 3270 -13441
rect 3000 -13601 3270 -13559
rect 3000 -13719 3076 -13601
rect 3194 -13719 3270 -13601
rect 3000 -13761 3270 -13719
rect 3000 -13879 3076 -13761
rect 3194 -13879 3270 -13761
rect 3000 -13921 3270 -13879
rect 3000 -14039 3076 -13921
rect 3194 -14039 3270 -13921
rect 3000 -14081 3270 -14039
rect 3000 -14199 3076 -14081
rect 3194 -14199 3270 -14081
rect 3000 -14241 3270 -14199
rect 3000 -14359 3076 -14241
rect 3194 -14359 3270 -14241
rect 3000 -14401 3270 -14359
rect 3000 -14519 3076 -14401
rect 3194 -14519 3270 -14401
rect 3000 -14561 3270 -14519
rect 3000 -14679 3076 -14561
rect 3194 -14679 3270 -14561
rect 3000 -14721 3270 -14679
rect 3000 -14839 3076 -14721
rect 3194 -14839 3270 -14721
rect 3000 -14881 3270 -14839
rect 3000 -14999 3076 -14881
rect 3194 -14999 3270 -14881
rect 3000 -15041 3270 -14999
rect 3000 -15159 3076 -15041
rect 3194 -15159 3270 -15041
rect 3000 -15201 3270 -15159
rect 3000 -15319 3076 -15201
rect 3194 -15230 3270 -15201
rect 6730 -11799 6809 -11770
rect 6927 -11799 7000 -11681
rect 6730 -11841 7000 -11799
rect 6730 -11959 6809 -11841
rect 6927 -11959 7000 -11841
rect 6730 -12001 7000 -11959
rect 6730 -12119 6809 -12001
rect 6927 -12119 7000 -12001
rect 6730 -12161 7000 -12119
rect 6730 -12279 6809 -12161
rect 6927 -12279 7000 -12161
rect 6730 -12321 7000 -12279
rect 6730 -12439 6809 -12321
rect 6927 -12439 7000 -12321
rect 6730 -12481 7000 -12439
rect 6730 -12599 6809 -12481
rect 6927 -12599 7000 -12481
rect 6730 -12641 7000 -12599
rect 6730 -12759 6809 -12641
rect 6927 -12759 7000 -12641
rect 6730 -12801 7000 -12759
rect 6730 -12919 6809 -12801
rect 6927 -12919 7000 -12801
rect 6730 -12961 7000 -12919
rect 6730 -13079 6809 -12961
rect 6927 -13079 7000 -12961
rect 6730 -13121 7000 -13079
rect 6730 -13239 6809 -13121
rect 6927 -13239 7000 -13121
rect 6730 -13281 7000 -13239
rect 6730 -13399 6809 -13281
rect 6927 -13399 7000 -13281
rect 6730 -13441 7000 -13399
rect 6730 -13559 6809 -13441
rect 6927 -13559 7000 -13441
rect 6730 -13601 7000 -13559
rect 6730 -13719 6809 -13601
rect 6927 -13719 7000 -13601
rect 6730 -13761 7000 -13719
rect 6730 -13879 6809 -13761
rect 6927 -13879 7000 -13761
rect 6730 -13921 7000 -13879
rect 6730 -14039 6809 -13921
rect 6927 -14039 7000 -13921
rect 6730 -14081 7000 -14039
rect 6730 -14199 6809 -14081
rect 6927 -14199 7000 -14081
rect 6730 -14241 7000 -14199
rect 6730 -14359 6809 -14241
rect 6927 -14359 7000 -14241
rect 6730 -14401 7000 -14359
rect 6730 -14519 6809 -14401
rect 6927 -14519 7000 -14401
rect 6730 -14561 7000 -14519
rect 6730 -14679 6809 -14561
rect 6927 -14679 7000 -14561
rect 6730 -14721 7000 -14679
rect 6730 -14839 6809 -14721
rect 6927 -14839 7000 -14721
rect 6730 -14881 7000 -14839
rect 6730 -14999 6809 -14881
rect 6927 -14999 7000 -14881
rect 6730 -15041 7000 -14999
rect 6730 -15159 6809 -15041
rect 6927 -15159 7000 -15041
rect 6730 -15201 7000 -15159
rect 6730 -15230 6809 -15201
rect 3194 -15306 6809 -15230
rect 3194 -15319 3261 -15306
rect 3000 -15424 3261 -15319
rect 3379 -15424 3421 -15306
rect 3539 -15424 3581 -15306
rect 3699 -15424 3741 -15306
rect 3859 -15424 3901 -15306
rect 4019 -15424 4061 -15306
rect 4179 -15424 4221 -15306
rect 4339 -15424 4381 -15306
rect 4499 -15424 4541 -15306
rect 4659 -15424 4701 -15306
rect 4819 -15424 4861 -15306
rect 4979 -15424 5021 -15306
rect 5139 -15424 5181 -15306
rect 5299 -15424 5341 -15306
rect 5459 -15424 5501 -15306
rect 5619 -15424 5661 -15306
rect 5779 -15424 5821 -15306
rect 5939 -15424 5981 -15306
rect 6099 -15424 6141 -15306
rect 6259 -15424 6301 -15306
rect 6419 -15424 6461 -15306
rect 6579 -15424 6621 -15306
rect 6739 -15319 6809 -15306
rect 6927 -15319 7000 -15201
rect 6739 -15424 7000 -15319
rect 3000 -15500 7000 -15424
rect 9000 -11578 13000 -11500
rect 9000 -11681 9261 -11578
rect 9000 -11799 9076 -11681
rect 9194 -11696 9261 -11681
rect 9379 -11696 9421 -11578
rect 9539 -11696 9581 -11578
rect 9699 -11696 9741 -11578
rect 9859 -11696 9901 -11578
rect 10019 -11696 10061 -11578
rect 10179 -11696 10221 -11578
rect 10339 -11696 10381 -11578
rect 10499 -11696 10541 -11578
rect 10659 -11696 10701 -11578
rect 10819 -11696 10861 -11578
rect 10979 -11696 11021 -11578
rect 11139 -11696 11181 -11578
rect 11299 -11696 11341 -11578
rect 11459 -11696 11501 -11578
rect 11619 -11696 11661 -11578
rect 11779 -11696 11821 -11578
rect 11939 -11696 11981 -11578
rect 12099 -11696 12141 -11578
rect 12259 -11696 12301 -11578
rect 12419 -11696 12461 -11578
rect 12579 -11696 12621 -11578
rect 12739 -11681 13000 -11578
rect 12739 -11696 12809 -11681
rect 9194 -11770 12809 -11696
rect 9194 -11799 9270 -11770
rect 9000 -11841 9270 -11799
rect 9000 -11959 9076 -11841
rect 9194 -11959 9270 -11841
rect 9000 -12001 9270 -11959
rect 9000 -12119 9076 -12001
rect 9194 -12119 9270 -12001
rect 9000 -12161 9270 -12119
rect 9000 -12279 9076 -12161
rect 9194 -12279 9270 -12161
rect 9000 -12321 9270 -12279
rect 9000 -12439 9076 -12321
rect 9194 -12439 9270 -12321
rect 9000 -12481 9270 -12439
rect 9000 -12599 9076 -12481
rect 9194 -12599 9270 -12481
rect 9000 -12641 9270 -12599
rect 9000 -12759 9076 -12641
rect 9194 -12759 9270 -12641
rect 9000 -12801 9270 -12759
rect 9000 -12919 9076 -12801
rect 9194 -12919 9270 -12801
rect 9000 -12961 9270 -12919
rect 9000 -13079 9076 -12961
rect 9194 -13079 9270 -12961
rect 9000 -13121 9270 -13079
rect 9000 -13239 9076 -13121
rect 9194 -13239 9270 -13121
rect 9000 -13281 9270 -13239
rect 9000 -13399 9076 -13281
rect 9194 -13399 9270 -13281
rect 9000 -13441 9270 -13399
rect 9000 -13559 9076 -13441
rect 9194 -13559 9270 -13441
rect 9000 -13601 9270 -13559
rect 9000 -13719 9076 -13601
rect 9194 -13719 9270 -13601
rect 9000 -13761 9270 -13719
rect 9000 -13879 9076 -13761
rect 9194 -13879 9270 -13761
rect 9000 -13921 9270 -13879
rect 9000 -14039 9076 -13921
rect 9194 -14039 9270 -13921
rect 9000 -14081 9270 -14039
rect 9000 -14199 9076 -14081
rect 9194 -14199 9270 -14081
rect 9000 -14241 9270 -14199
rect 9000 -14359 9076 -14241
rect 9194 -14359 9270 -14241
rect 9000 -14401 9270 -14359
rect 9000 -14519 9076 -14401
rect 9194 -14519 9270 -14401
rect 9000 -14561 9270 -14519
rect 9000 -14679 9076 -14561
rect 9194 -14679 9270 -14561
rect 9000 -14721 9270 -14679
rect 9000 -14839 9076 -14721
rect 9194 -14839 9270 -14721
rect 9000 -14881 9270 -14839
rect 9000 -14999 9076 -14881
rect 9194 -14999 9270 -14881
rect 9000 -15041 9270 -14999
rect 9000 -15159 9076 -15041
rect 9194 -15159 9270 -15041
rect 9000 -15201 9270 -15159
rect 9000 -15319 9076 -15201
rect 9194 -15230 9270 -15201
rect 12730 -11799 12809 -11770
rect 12927 -11799 13000 -11681
rect 12730 -11841 13000 -11799
rect 12730 -11959 12809 -11841
rect 12927 -11959 13000 -11841
rect 12730 -12001 13000 -11959
rect 12730 -12119 12809 -12001
rect 12927 -12119 13000 -12001
rect 12730 -12161 13000 -12119
rect 12730 -12279 12809 -12161
rect 12927 -12279 13000 -12161
rect 12730 -12321 13000 -12279
rect 12730 -12439 12809 -12321
rect 12927 -12439 13000 -12321
rect 12730 -12481 13000 -12439
rect 12730 -12599 12809 -12481
rect 12927 -12599 13000 -12481
rect 12730 -12641 13000 -12599
rect 12730 -12759 12809 -12641
rect 12927 -12759 13000 -12641
rect 12730 -12801 13000 -12759
rect 12730 -12919 12809 -12801
rect 12927 -12919 13000 -12801
rect 12730 -12961 13000 -12919
rect 12730 -13079 12809 -12961
rect 12927 -13079 13000 -12961
rect 12730 -13121 13000 -13079
rect 12730 -13239 12809 -13121
rect 12927 -13239 13000 -13121
rect 12730 -13281 13000 -13239
rect 12730 -13399 12809 -13281
rect 12927 -13399 13000 -13281
rect 12730 -13441 13000 -13399
rect 12730 -13559 12809 -13441
rect 12927 -13559 13000 -13441
rect 12730 -13601 13000 -13559
rect 12730 -13719 12809 -13601
rect 12927 -13719 13000 -13601
rect 12730 -13761 13000 -13719
rect 12730 -13879 12809 -13761
rect 12927 -13879 13000 -13761
rect 12730 -13921 13000 -13879
rect 12730 -14039 12809 -13921
rect 12927 -14039 13000 -13921
rect 12730 -14081 13000 -14039
rect 12730 -14199 12809 -14081
rect 12927 -14199 13000 -14081
rect 12730 -14241 13000 -14199
rect 12730 -14359 12809 -14241
rect 12927 -14359 13000 -14241
rect 12730 -14401 13000 -14359
rect 12730 -14519 12809 -14401
rect 12927 -14519 13000 -14401
rect 12730 -14561 13000 -14519
rect 12730 -14679 12809 -14561
rect 12927 -14679 13000 -14561
rect 12730 -14721 13000 -14679
rect 12730 -14839 12809 -14721
rect 12927 -14839 13000 -14721
rect 12730 -14881 13000 -14839
rect 12730 -14999 12809 -14881
rect 12927 -14999 13000 -14881
rect 12730 -15041 13000 -14999
rect 12730 -15159 12809 -15041
rect 12927 -15159 13000 -15041
rect 12730 -15201 13000 -15159
rect 12730 -15230 12809 -15201
rect 9194 -15306 12809 -15230
rect 9194 -15319 9261 -15306
rect 9000 -15424 9261 -15319
rect 9379 -15424 9421 -15306
rect 9539 -15424 9581 -15306
rect 9699 -15424 9741 -15306
rect 9859 -15424 9901 -15306
rect 10019 -15424 10061 -15306
rect 10179 -15424 10221 -15306
rect 10339 -15424 10381 -15306
rect 10499 -15424 10541 -15306
rect 10659 -15424 10701 -15306
rect 10819 -15424 10861 -15306
rect 10979 -15424 11021 -15306
rect 11139 -15424 11181 -15306
rect 11299 -15424 11341 -15306
rect 11459 -15424 11501 -15306
rect 11619 -15424 11661 -15306
rect 11779 -15424 11821 -15306
rect 11939 -15424 11981 -15306
rect 12099 -15424 12141 -15306
rect 12259 -15424 12301 -15306
rect 12419 -15424 12461 -15306
rect 12579 -15424 12621 -15306
rect 12739 -15319 12809 -15306
rect 12927 -15319 13000 -15201
rect 12739 -15424 13000 -15319
rect 9000 -15500 13000 -15424
rect 15000 -11578 19000 -11500
rect 15000 -11681 15261 -11578
rect 15000 -11799 15076 -11681
rect 15194 -11696 15261 -11681
rect 15379 -11696 15421 -11578
rect 15539 -11696 15581 -11578
rect 15699 -11696 15741 -11578
rect 15859 -11696 15901 -11578
rect 16019 -11696 16061 -11578
rect 16179 -11696 16221 -11578
rect 16339 -11696 16381 -11578
rect 16499 -11696 16541 -11578
rect 16659 -11696 16701 -11578
rect 16819 -11696 16861 -11578
rect 16979 -11696 17021 -11578
rect 17139 -11696 17181 -11578
rect 17299 -11696 17341 -11578
rect 17459 -11696 17501 -11578
rect 17619 -11696 17661 -11578
rect 17779 -11696 17821 -11578
rect 17939 -11696 17981 -11578
rect 18099 -11696 18141 -11578
rect 18259 -11696 18301 -11578
rect 18419 -11696 18461 -11578
rect 18579 -11696 18621 -11578
rect 18739 -11681 19000 -11578
rect 18739 -11696 18809 -11681
rect 15194 -11770 18809 -11696
rect 15194 -11799 15270 -11770
rect 15000 -11841 15270 -11799
rect 15000 -11959 15076 -11841
rect 15194 -11959 15270 -11841
rect 15000 -12001 15270 -11959
rect 15000 -12119 15076 -12001
rect 15194 -12119 15270 -12001
rect 15000 -12161 15270 -12119
rect 15000 -12279 15076 -12161
rect 15194 -12279 15270 -12161
rect 15000 -12321 15270 -12279
rect 15000 -12439 15076 -12321
rect 15194 -12439 15270 -12321
rect 15000 -12481 15270 -12439
rect 15000 -12599 15076 -12481
rect 15194 -12599 15270 -12481
rect 15000 -12641 15270 -12599
rect 15000 -12759 15076 -12641
rect 15194 -12759 15270 -12641
rect 15000 -12801 15270 -12759
rect 15000 -12919 15076 -12801
rect 15194 -12919 15270 -12801
rect 15000 -12961 15270 -12919
rect 15000 -13079 15076 -12961
rect 15194 -13079 15270 -12961
rect 15000 -13121 15270 -13079
rect 15000 -13239 15076 -13121
rect 15194 -13239 15270 -13121
rect 15000 -13281 15270 -13239
rect 15000 -13399 15076 -13281
rect 15194 -13399 15270 -13281
rect 15000 -13441 15270 -13399
rect 15000 -13559 15076 -13441
rect 15194 -13559 15270 -13441
rect 15000 -13601 15270 -13559
rect 15000 -13719 15076 -13601
rect 15194 -13719 15270 -13601
rect 15000 -13761 15270 -13719
rect 15000 -13879 15076 -13761
rect 15194 -13879 15270 -13761
rect 15000 -13921 15270 -13879
rect 15000 -14039 15076 -13921
rect 15194 -14039 15270 -13921
rect 15000 -14081 15270 -14039
rect 15000 -14199 15076 -14081
rect 15194 -14199 15270 -14081
rect 15000 -14241 15270 -14199
rect 15000 -14359 15076 -14241
rect 15194 -14359 15270 -14241
rect 15000 -14401 15270 -14359
rect 15000 -14519 15076 -14401
rect 15194 -14519 15270 -14401
rect 15000 -14561 15270 -14519
rect 15000 -14679 15076 -14561
rect 15194 -14679 15270 -14561
rect 15000 -14721 15270 -14679
rect 15000 -14839 15076 -14721
rect 15194 -14839 15270 -14721
rect 15000 -14881 15270 -14839
rect 15000 -14999 15076 -14881
rect 15194 -14999 15270 -14881
rect 15000 -15041 15270 -14999
rect 15000 -15159 15076 -15041
rect 15194 -15159 15270 -15041
rect 15000 -15201 15270 -15159
rect 15000 -15319 15076 -15201
rect 15194 -15230 15270 -15201
rect 18730 -11799 18809 -11770
rect 18927 -11799 19000 -11681
rect 18730 -11841 19000 -11799
rect 18730 -11959 18809 -11841
rect 18927 -11959 19000 -11841
rect 18730 -12001 19000 -11959
rect 18730 -12119 18809 -12001
rect 18927 -12119 19000 -12001
rect 18730 -12161 19000 -12119
rect 18730 -12279 18809 -12161
rect 18927 -12279 19000 -12161
rect 18730 -12321 19000 -12279
rect 18730 -12439 18809 -12321
rect 18927 -12439 19000 -12321
rect 18730 -12481 19000 -12439
rect 18730 -12599 18809 -12481
rect 18927 -12599 19000 -12481
rect 18730 -12641 19000 -12599
rect 18730 -12759 18809 -12641
rect 18927 -12759 19000 -12641
rect 18730 -12801 19000 -12759
rect 18730 -12919 18809 -12801
rect 18927 -12919 19000 -12801
rect 18730 -12961 19000 -12919
rect 18730 -13079 18809 -12961
rect 18927 -13079 19000 -12961
rect 18730 -13121 19000 -13079
rect 18730 -13239 18809 -13121
rect 18927 -13239 19000 -13121
rect 18730 -13281 19000 -13239
rect 18730 -13399 18809 -13281
rect 18927 -13399 19000 -13281
rect 18730 -13441 19000 -13399
rect 18730 -13559 18809 -13441
rect 18927 -13559 19000 -13441
rect 18730 -13601 19000 -13559
rect 18730 -13719 18809 -13601
rect 18927 -13719 19000 -13601
rect 18730 -13761 19000 -13719
rect 18730 -13879 18809 -13761
rect 18927 -13879 19000 -13761
rect 18730 -13921 19000 -13879
rect 18730 -14039 18809 -13921
rect 18927 -14039 19000 -13921
rect 18730 -14081 19000 -14039
rect 18730 -14199 18809 -14081
rect 18927 -14199 19000 -14081
rect 18730 -14241 19000 -14199
rect 18730 -14359 18809 -14241
rect 18927 -14359 19000 -14241
rect 18730 -14401 19000 -14359
rect 18730 -14519 18809 -14401
rect 18927 -14519 19000 -14401
rect 18730 -14561 19000 -14519
rect 18730 -14679 18809 -14561
rect 18927 -14679 19000 -14561
rect 18730 -14721 19000 -14679
rect 18730 -14839 18809 -14721
rect 18927 -14839 19000 -14721
rect 18730 -14881 19000 -14839
rect 18730 -14999 18809 -14881
rect 18927 -14999 19000 -14881
rect 18730 -15041 19000 -14999
rect 18730 -15159 18809 -15041
rect 18927 -15159 19000 -15041
rect 18730 -15201 19000 -15159
rect 18730 -15230 18809 -15201
rect 15194 -15306 18809 -15230
rect 15194 -15319 15261 -15306
rect 15000 -15424 15261 -15319
rect 15379 -15424 15421 -15306
rect 15539 -15424 15581 -15306
rect 15699 -15424 15741 -15306
rect 15859 -15424 15901 -15306
rect 16019 -15424 16061 -15306
rect 16179 -15424 16221 -15306
rect 16339 -15424 16381 -15306
rect 16499 -15424 16541 -15306
rect 16659 -15424 16701 -15306
rect 16819 -15424 16861 -15306
rect 16979 -15424 17021 -15306
rect 17139 -15424 17181 -15306
rect 17299 -15424 17341 -15306
rect 17459 -15424 17501 -15306
rect 17619 -15424 17661 -15306
rect 17779 -15424 17821 -15306
rect 17939 -15424 17981 -15306
rect 18099 -15424 18141 -15306
rect 18259 -15424 18301 -15306
rect 18419 -15424 18461 -15306
rect 18579 -15424 18621 -15306
rect 18739 -15319 18809 -15306
rect 18927 -15319 19000 -15201
rect 18739 -15424 19000 -15319
rect 15000 -15500 19000 -15424
rect 21000 -11578 25000 -11500
rect 21000 -11681 21261 -11578
rect 21000 -11799 21076 -11681
rect 21194 -11696 21261 -11681
rect 21379 -11696 21421 -11578
rect 21539 -11696 21581 -11578
rect 21699 -11696 21741 -11578
rect 21859 -11696 21901 -11578
rect 22019 -11696 22061 -11578
rect 22179 -11696 22221 -11578
rect 22339 -11696 22381 -11578
rect 22499 -11696 22541 -11578
rect 22659 -11696 22701 -11578
rect 22819 -11696 22861 -11578
rect 22979 -11696 23021 -11578
rect 23139 -11696 23181 -11578
rect 23299 -11696 23341 -11578
rect 23459 -11696 23501 -11578
rect 23619 -11696 23661 -11578
rect 23779 -11696 23821 -11578
rect 23939 -11696 23981 -11578
rect 24099 -11696 24141 -11578
rect 24259 -11696 24301 -11578
rect 24419 -11696 24461 -11578
rect 24579 -11696 24621 -11578
rect 24739 -11681 25000 -11578
rect 24739 -11696 24809 -11681
rect 21194 -11770 24809 -11696
rect 21194 -11799 21270 -11770
rect 21000 -11841 21270 -11799
rect 21000 -11959 21076 -11841
rect 21194 -11959 21270 -11841
rect 21000 -12001 21270 -11959
rect 21000 -12119 21076 -12001
rect 21194 -12119 21270 -12001
rect 21000 -12161 21270 -12119
rect 21000 -12279 21076 -12161
rect 21194 -12279 21270 -12161
rect 21000 -12321 21270 -12279
rect 21000 -12439 21076 -12321
rect 21194 -12439 21270 -12321
rect 21000 -12481 21270 -12439
rect 21000 -12599 21076 -12481
rect 21194 -12599 21270 -12481
rect 21000 -12641 21270 -12599
rect 21000 -12759 21076 -12641
rect 21194 -12759 21270 -12641
rect 21000 -12801 21270 -12759
rect 21000 -12919 21076 -12801
rect 21194 -12919 21270 -12801
rect 21000 -12961 21270 -12919
rect 21000 -13079 21076 -12961
rect 21194 -13079 21270 -12961
rect 21000 -13121 21270 -13079
rect 21000 -13239 21076 -13121
rect 21194 -13239 21270 -13121
rect 21000 -13281 21270 -13239
rect 21000 -13399 21076 -13281
rect 21194 -13399 21270 -13281
rect 21000 -13441 21270 -13399
rect 21000 -13559 21076 -13441
rect 21194 -13559 21270 -13441
rect 21000 -13601 21270 -13559
rect 21000 -13719 21076 -13601
rect 21194 -13719 21270 -13601
rect 21000 -13761 21270 -13719
rect 21000 -13879 21076 -13761
rect 21194 -13879 21270 -13761
rect 21000 -13921 21270 -13879
rect 21000 -14039 21076 -13921
rect 21194 -14039 21270 -13921
rect 21000 -14081 21270 -14039
rect 21000 -14199 21076 -14081
rect 21194 -14199 21270 -14081
rect 21000 -14241 21270 -14199
rect 21000 -14359 21076 -14241
rect 21194 -14359 21270 -14241
rect 21000 -14401 21270 -14359
rect 21000 -14519 21076 -14401
rect 21194 -14519 21270 -14401
rect 21000 -14561 21270 -14519
rect 21000 -14679 21076 -14561
rect 21194 -14679 21270 -14561
rect 21000 -14721 21270 -14679
rect 21000 -14839 21076 -14721
rect 21194 -14839 21270 -14721
rect 21000 -14881 21270 -14839
rect 21000 -14999 21076 -14881
rect 21194 -14999 21270 -14881
rect 21000 -15041 21270 -14999
rect 21000 -15159 21076 -15041
rect 21194 -15159 21270 -15041
rect 21000 -15201 21270 -15159
rect 21000 -15319 21076 -15201
rect 21194 -15230 21270 -15201
rect 24730 -11799 24809 -11770
rect 24927 -11799 25000 -11681
rect 24730 -11841 25000 -11799
rect 24730 -11959 24809 -11841
rect 24927 -11959 25000 -11841
rect 24730 -12001 25000 -11959
rect 24730 -12119 24809 -12001
rect 24927 -12119 25000 -12001
rect 24730 -12161 25000 -12119
rect 24730 -12279 24809 -12161
rect 24927 -12279 25000 -12161
rect 24730 -12321 25000 -12279
rect 24730 -12439 24809 -12321
rect 24927 -12439 25000 -12321
rect 24730 -12481 25000 -12439
rect 24730 -12599 24809 -12481
rect 24927 -12599 25000 -12481
rect 24730 -12641 25000 -12599
rect 24730 -12759 24809 -12641
rect 24927 -12759 25000 -12641
rect 24730 -12801 25000 -12759
rect 24730 -12919 24809 -12801
rect 24927 -12919 25000 -12801
rect 24730 -12961 25000 -12919
rect 24730 -13079 24809 -12961
rect 24927 -13079 25000 -12961
rect 24730 -13121 25000 -13079
rect 24730 -13239 24809 -13121
rect 24927 -13239 25000 -13121
rect 24730 -13281 25000 -13239
rect 24730 -13399 24809 -13281
rect 24927 -13399 25000 -13281
rect 24730 -13441 25000 -13399
rect 24730 -13559 24809 -13441
rect 24927 -13559 25000 -13441
rect 24730 -13601 25000 -13559
rect 24730 -13719 24809 -13601
rect 24927 -13719 25000 -13601
rect 24730 -13761 25000 -13719
rect 24730 -13879 24809 -13761
rect 24927 -13879 25000 -13761
rect 24730 -13921 25000 -13879
rect 24730 -14039 24809 -13921
rect 24927 -14039 25000 -13921
rect 24730 -14081 25000 -14039
rect 24730 -14199 24809 -14081
rect 24927 -14199 25000 -14081
rect 24730 -14241 25000 -14199
rect 24730 -14359 24809 -14241
rect 24927 -14359 25000 -14241
rect 24730 -14401 25000 -14359
rect 24730 -14519 24809 -14401
rect 24927 -14519 25000 -14401
rect 24730 -14561 25000 -14519
rect 24730 -14679 24809 -14561
rect 24927 -14679 25000 -14561
rect 24730 -14721 25000 -14679
rect 24730 -14839 24809 -14721
rect 24927 -14839 25000 -14721
rect 24730 -14881 25000 -14839
rect 24730 -14999 24809 -14881
rect 24927 -14999 25000 -14881
rect 24730 -15041 25000 -14999
rect 24730 -15159 24809 -15041
rect 24927 -15159 25000 -15041
rect 24730 -15201 25000 -15159
rect 24730 -15230 24809 -15201
rect 21194 -15306 24809 -15230
rect 21194 -15319 21261 -15306
rect 21000 -15424 21261 -15319
rect 21379 -15424 21421 -15306
rect 21539 -15424 21581 -15306
rect 21699 -15424 21741 -15306
rect 21859 -15424 21901 -15306
rect 22019 -15424 22061 -15306
rect 22179 -15424 22221 -15306
rect 22339 -15424 22381 -15306
rect 22499 -15424 22541 -15306
rect 22659 -15424 22701 -15306
rect 22819 -15424 22861 -15306
rect 22979 -15424 23021 -15306
rect 23139 -15424 23181 -15306
rect 23299 -15424 23341 -15306
rect 23459 -15424 23501 -15306
rect 23619 -15424 23661 -15306
rect 23779 -15424 23821 -15306
rect 23939 -15424 23981 -15306
rect 24099 -15424 24141 -15306
rect 24259 -15424 24301 -15306
rect 24419 -15424 24461 -15306
rect 24579 -15424 24621 -15306
rect 24739 -15319 24809 -15306
rect 24927 -15319 25000 -15201
rect 24739 -15424 25000 -15319
rect 21000 -15500 25000 -15424
<< via4 >>
rect 3261 9381 3379 9424
rect 3261 9349 3304 9381
rect 3304 9349 3336 9381
rect 3336 9349 3379 9381
rect 3073 9276 3191 9319
rect 3261 9306 3379 9349
rect 3421 9381 3539 9424
rect 3421 9349 3464 9381
rect 3464 9349 3496 9381
rect 3496 9349 3539 9381
rect 3421 9306 3539 9349
rect 3581 9381 3699 9424
rect 3581 9349 3624 9381
rect 3624 9349 3656 9381
rect 3656 9349 3699 9381
rect 3581 9306 3699 9349
rect 3741 9381 3859 9424
rect 3741 9349 3784 9381
rect 3784 9349 3816 9381
rect 3816 9349 3859 9381
rect 3741 9306 3859 9349
rect 3901 9381 4019 9424
rect 3901 9349 3944 9381
rect 3944 9349 3976 9381
rect 3976 9349 4019 9381
rect 3901 9306 4019 9349
rect 4061 9381 4179 9424
rect 4061 9349 4104 9381
rect 4104 9349 4136 9381
rect 4136 9349 4179 9381
rect 4061 9306 4179 9349
rect 4221 9381 4339 9424
rect 4221 9349 4264 9381
rect 4264 9349 4296 9381
rect 4296 9349 4339 9381
rect 4221 9306 4339 9349
rect 4381 9381 4499 9424
rect 4381 9349 4424 9381
rect 4424 9349 4456 9381
rect 4456 9349 4499 9381
rect 4381 9306 4499 9349
rect 4541 9381 4659 9424
rect 4541 9349 4584 9381
rect 4584 9349 4616 9381
rect 4616 9349 4659 9381
rect 4541 9306 4659 9349
rect 4701 9381 4819 9424
rect 4701 9349 4744 9381
rect 4744 9349 4776 9381
rect 4776 9349 4819 9381
rect 4701 9306 4819 9349
rect 4861 9381 4979 9424
rect 4861 9349 4904 9381
rect 4904 9349 4936 9381
rect 4936 9349 4979 9381
rect 4861 9306 4979 9349
rect 5021 9381 5139 9424
rect 5021 9349 5064 9381
rect 5064 9349 5096 9381
rect 5096 9349 5139 9381
rect 5021 9306 5139 9349
rect 5181 9381 5299 9424
rect 5181 9349 5224 9381
rect 5224 9349 5256 9381
rect 5256 9349 5299 9381
rect 5181 9306 5299 9349
rect 5341 9381 5459 9424
rect 5341 9349 5384 9381
rect 5384 9349 5416 9381
rect 5416 9349 5459 9381
rect 5341 9306 5459 9349
rect 5501 9381 5619 9424
rect 5501 9349 5544 9381
rect 5544 9349 5576 9381
rect 5576 9349 5619 9381
rect 5501 9306 5619 9349
rect 5661 9381 5779 9424
rect 5661 9349 5704 9381
rect 5704 9349 5736 9381
rect 5736 9349 5779 9381
rect 5661 9306 5779 9349
rect 5821 9381 5939 9424
rect 5821 9349 5864 9381
rect 5864 9349 5896 9381
rect 5896 9349 5939 9381
rect 5821 9306 5939 9349
rect 5981 9381 6099 9424
rect 5981 9349 6024 9381
rect 6024 9349 6056 9381
rect 6056 9349 6099 9381
rect 5981 9306 6099 9349
rect 6141 9381 6259 9424
rect 6141 9349 6184 9381
rect 6184 9349 6216 9381
rect 6216 9349 6259 9381
rect 6141 9306 6259 9349
rect 6301 9381 6419 9424
rect 6301 9349 6344 9381
rect 6344 9349 6376 9381
rect 6376 9349 6419 9381
rect 6301 9306 6419 9349
rect 6461 9381 6579 9424
rect 6461 9349 6504 9381
rect 6504 9349 6536 9381
rect 6536 9349 6579 9381
rect 6461 9306 6579 9349
rect 6621 9381 6739 9424
rect 6621 9349 6664 9381
rect 6664 9349 6696 9381
rect 6696 9349 6739 9381
rect 6621 9306 6739 9349
rect 3073 9244 3116 9276
rect 3116 9244 3148 9276
rect 3148 9244 3191 9276
rect 3073 9201 3191 9244
rect 6806 9276 6924 9319
rect 6806 9244 6849 9276
rect 6849 9244 6881 9276
rect 6881 9244 6924 9276
rect 3073 9116 3191 9159
rect 3073 9084 3116 9116
rect 3116 9084 3148 9116
rect 3148 9084 3191 9116
rect 3073 9041 3191 9084
rect 3073 8956 3191 8999
rect 3073 8924 3116 8956
rect 3116 8924 3148 8956
rect 3148 8924 3191 8956
rect 3073 8881 3191 8924
rect 3073 8796 3191 8839
rect 3073 8764 3116 8796
rect 3116 8764 3148 8796
rect 3148 8764 3191 8796
rect 3073 8721 3191 8764
rect 3073 8636 3191 8679
rect 3073 8604 3116 8636
rect 3116 8604 3148 8636
rect 3148 8604 3191 8636
rect 3073 8561 3191 8604
rect 3073 8476 3191 8519
rect 3073 8444 3116 8476
rect 3116 8444 3148 8476
rect 3148 8444 3191 8476
rect 3073 8401 3191 8444
rect 3073 8316 3191 8359
rect 3073 8284 3116 8316
rect 3116 8284 3148 8316
rect 3148 8284 3191 8316
rect 3073 8241 3191 8284
rect 3073 8156 3191 8199
rect 3073 8124 3116 8156
rect 3116 8124 3148 8156
rect 3148 8124 3191 8156
rect 3073 8081 3191 8124
rect 3073 7996 3191 8039
rect 3073 7964 3116 7996
rect 3116 7964 3148 7996
rect 3148 7964 3191 7996
rect 3073 7921 3191 7964
rect 3073 7836 3191 7879
rect 3073 7804 3116 7836
rect 3116 7804 3148 7836
rect 3148 7804 3191 7836
rect 3073 7761 3191 7804
rect 3073 7676 3191 7719
rect 3073 7644 3116 7676
rect 3116 7644 3148 7676
rect 3148 7644 3191 7676
rect 3073 7601 3191 7644
rect 3073 7516 3191 7559
rect 3073 7484 3116 7516
rect 3116 7484 3148 7516
rect 3148 7484 3191 7516
rect 3073 7441 3191 7484
rect 3073 7356 3191 7399
rect 3073 7324 3116 7356
rect 3116 7324 3148 7356
rect 3148 7324 3191 7356
rect 3073 7281 3191 7324
rect 3073 7196 3191 7239
rect 3073 7164 3116 7196
rect 3116 7164 3148 7196
rect 3148 7164 3191 7196
rect 3073 7121 3191 7164
rect 3073 7036 3191 7079
rect 3073 7004 3116 7036
rect 3116 7004 3148 7036
rect 3148 7004 3191 7036
rect 3073 6961 3191 7004
rect 3073 6876 3191 6919
rect 3073 6844 3116 6876
rect 3116 6844 3148 6876
rect 3148 6844 3191 6876
rect 3073 6801 3191 6844
rect 3073 6716 3191 6759
rect 3073 6684 3116 6716
rect 3116 6684 3148 6716
rect 3148 6684 3191 6716
rect 3073 6641 3191 6684
rect 3073 6556 3191 6599
rect 3073 6524 3116 6556
rect 3116 6524 3148 6556
rect 3148 6524 3191 6556
rect 3073 6481 3191 6524
rect 3073 6396 3191 6439
rect 3073 6364 3116 6396
rect 3116 6364 3148 6396
rect 3148 6364 3191 6396
rect 3073 6321 3191 6364
rect 3073 6236 3191 6279
rect 3073 6204 3116 6236
rect 3116 6204 3148 6236
rect 3148 6204 3191 6236
rect 3073 6161 3191 6204
rect 3073 6076 3191 6119
rect 3073 6044 3116 6076
rect 3116 6044 3148 6076
rect 3148 6044 3191 6076
rect 3073 6001 3191 6044
rect 3073 5916 3191 5959
rect 3073 5884 3116 5916
rect 3116 5884 3148 5916
rect 3148 5884 3191 5916
rect 3073 5841 3191 5884
rect 3073 5756 3191 5799
rect 6806 9201 6924 9244
rect 6806 9116 6924 9159
rect 6806 9084 6849 9116
rect 6849 9084 6881 9116
rect 6881 9084 6924 9116
rect 6806 9041 6924 9084
rect 6806 8956 6924 8999
rect 6806 8924 6849 8956
rect 6849 8924 6881 8956
rect 6881 8924 6924 8956
rect 6806 8881 6924 8924
rect 6806 8796 6924 8839
rect 6806 8764 6849 8796
rect 6849 8764 6881 8796
rect 6881 8764 6924 8796
rect 6806 8721 6924 8764
rect 6806 8636 6924 8679
rect 6806 8604 6849 8636
rect 6849 8604 6881 8636
rect 6881 8604 6924 8636
rect 6806 8561 6924 8604
rect 6806 8476 6924 8519
rect 6806 8444 6849 8476
rect 6849 8444 6881 8476
rect 6881 8444 6924 8476
rect 6806 8401 6924 8444
rect 6806 8316 6924 8359
rect 6806 8284 6849 8316
rect 6849 8284 6881 8316
rect 6881 8284 6924 8316
rect 6806 8241 6924 8284
rect 6806 8156 6924 8199
rect 6806 8124 6849 8156
rect 6849 8124 6881 8156
rect 6881 8124 6924 8156
rect 6806 8081 6924 8124
rect 6806 7996 6924 8039
rect 6806 7964 6849 7996
rect 6849 7964 6881 7996
rect 6881 7964 6924 7996
rect 6806 7921 6924 7964
rect 6806 7836 6924 7879
rect 6806 7804 6849 7836
rect 6849 7804 6881 7836
rect 6881 7804 6924 7836
rect 6806 7761 6924 7804
rect 6806 7676 6924 7719
rect 6806 7644 6849 7676
rect 6849 7644 6881 7676
rect 6881 7644 6924 7676
rect 6806 7601 6924 7644
rect 6806 7516 6924 7559
rect 6806 7484 6849 7516
rect 6849 7484 6881 7516
rect 6881 7484 6924 7516
rect 6806 7441 6924 7484
rect 6806 7356 6924 7399
rect 6806 7324 6849 7356
rect 6849 7324 6881 7356
rect 6881 7324 6924 7356
rect 6806 7281 6924 7324
rect 6806 7196 6924 7239
rect 6806 7164 6849 7196
rect 6849 7164 6881 7196
rect 6881 7164 6924 7196
rect 6806 7121 6924 7164
rect 6806 7036 6924 7079
rect 6806 7004 6849 7036
rect 6849 7004 6881 7036
rect 6881 7004 6924 7036
rect 6806 6961 6924 7004
rect 6806 6876 6924 6919
rect 6806 6844 6849 6876
rect 6849 6844 6881 6876
rect 6881 6844 6924 6876
rect 6806 6801 6924 6844
rect 6806 6716 6924 6759
rect 6806 6684 6849 6716
rect 6849 6684 6881 6716
rect 6881 6684 6924 6716
rect 6806 6641 6924 6684
rect 6806 6556 6924 6599
rect 6806 6524 6849 6556
rect 6849 6524 6881 6556
rect 6881 6524 6924 6556
rect 6806 6481 6924 6524
rect 6806 6396 6924 6439
rect 6806 6364 6849 6396
rect 6849 6364 6881 6396
rect 6881 6364 6924 6396
rect 6806 6321 6924 6364
rect 6806 6236 6924 6279
rect 6806 6204 6849 6236
rect 6849 6204 6881 6236
rect 6881 6204 6924 6236
rect 6806 6161 6924 6204
rect 6806 6076 6924 6119
rect 6806 6044 6849 6076
rect 6849 6044 6881 6076
rect 6881 6044 6924 6076
rect 6806 6001 6924 6044
rect 6806 5916 6924 5959
rect 6806 5884 6849 5916
rect 6849 5884 6881 5916
rect 6881 5884 6924 5916
rect 6806 5841 6924 5884
rect 3073 5724 3116 5756
rect 3116 5724 3148 5756
rect 3148 5724 3191 5756
rect 3073 5681 3191 5724
rect 6806 5756 6924 5799
rect 6806 5724 6849 5756
rect 6849 5724 6881 5756
rect 6881 5724 6924 5756
rect 3261 5653 3379 5696
rect 3261 5621 3304 5653
rect 3304 5621 3336 5653
rect 3336 5621 3379 5653
rect 3261 5578 3379 5621
rect 3421 5653 3539 5696
rect 3421 5621 3464 5653
rect 3464 5621 3496 5653
rect 3496 5621 3539 5653
rect 3421 5578 3539 5621
rect 3581 5653 3699 5696
rect 3581 5621 3624 5653
rect 3624 5621 3656 5653
rect 3656 5621 3699 5653
rect 3581 5578 3699 5621
rect 3741 5653 3859 5696
rect 3741 5621 3784 5653
rect 3784 5621 3816 5653
rect 3816 5621 3859 5653
rect 3741 5578 3859 5621
rect 3901 5653 4019 5696
rect 3901 5621 3944 5653
rect 3944 5621 3976 5653
rect 3976 5621 4019 5653
rect 3901 5578 4019 5621
rect 4061 5653 4179 5696
rect 4061 5621 4104 5653
rect 4104 5621 4136 5653
rect 4136 5621 4179 5653
rect 4061 5578 4179 5621
rect 4221 5653 4339 5696
rect 4221 5621 4264 5653
rect 4264 5621 4296 5653
rect 4296 5621 4339 5653
rect 4221 5578 4339 5621
rect 4381 5653 4499 5696
rect 4381 5621 4424 5653
rect 4424 5621 4456 5653
rect 4456 5621 4499 5653
rect 4381 5578 4499 5621
rect 4541 5653 4659 5696
rect 4541 5621 4584 5653
rect 4584 5621 4616 5653
rect 4616 5621 4659 5653
rect 4541 5578 4659 5621
rect 4701 5653 4819 5696
rect 4701 5621 4744 5653
rect 4744 5621 4776 5653
rect 4776 5621 4819 5653
rect 4701 5578 4819 5621
rect 4861 5653 4979 5696
rect 4861 5621 4904 5653
rect 4904 5621 4936 5653
rect 4936 5621 4979 5653
rect 4861 5578 4979 5621
rect 5021 5653 5139 5696
rect 5021 5621 5064 5653
rect 5064 5621 5096 5653
rect 5096 5621 5139 5653
rect 5021 5578 5139 5621
rect 5181 5653 5299 5696
rect 5181 5621 5224 5653
rect 5224 5621 5256 5653
rect 5256 5621 5299 5653
rect 5181 5578 5299 5621
rect 5341 5653 5459 5696
rect 5341 5621 5384 5653
rect 5384 5621 5416 5653
rect 5416 5621 5459 5653
rect 5341 5578 5459 5621
rect 5501 5653 5619 5696
rect 5501 5621 5544 5653
rect 5544 5621 5576 5653
rect 5576 5621 5619 5653
rect 5501 5578 5619 5621
rect 5661 5653 5779 5696
rect 5661 5621 5704 5653
rect 5704 5621 5736 5653
rect 5736 5621 5779 5653
rect 5661 5578 5779 5621
rect 5821 5653 5939 5696
rect 5821 5621 5864 5653
rect 5864 5621 5896 5653
rect 5896 5621 5939 5653
rect 5821 5578 5939 5621
rect 5981 5653 6099 5696
rect 5981 5621 6024 5653
rect 6024 5621 6056 5653
rect 6056 5621 6099 5653
rect 5981 5578 6099 5621
rect 6141 5653 6259 5696
rect 6141 5621 6184 5653
rect 6184 5621 6216 5653
rect 6216 5621 6259 5653
rect 6141 5578 6259 5621
rect 6301 5653 6419 5696
rect 6301 5621 6344 5653
rect 6344 5621 6376 5653
rect 6376 5621 6419 5653
rect 6301 5578 6419 5621
rect 6461 5653 6579 5696
rect 6461 5621 6504 5653
rect 6504 5621 6536 5653
rect 6536 5621 6579 5653
rect 6461 5578 6579 5621
rect 6621 5653 6739 5696
rect 6806 5681 6924 5724
rect 6621 5621 6664 5653
rect 6664 5621 6696 5653
rect 6696 5621 6739 5653
rect 6621 5578 6739 5621
rect 9261 9381 9379 9424
rect 9261 9349 9304 9381
rect 9304 9349 9336 9381
rect 9336 9349 9379 9381
rect 9073 9276 9191 9319
rect 9261 9306 9379 9349
rect 9421 9381 9539 9424
rect 9421 9349 9464 9381
rect 9464 9349 9496 9381
rect 9496 9349 9539 9381
rect 9421 9306 9539 9349
rect 9581 9381 9699 9424
rect 9581 9349 9624 9381
rect 9624 9349 9656 9381
rect 9656 9349 9699 9381
rect 9581 9306 9699 9349
rect 9741 9381 9859 9424
rect 9741 9349 9784 9381
rect 9784 9349 9816 9381
rect 9816 9349 9859 9381
rect 9741 9306 9859 9349
rect 9901 9381 10019 9424
rect 9901 9349 9944 9381
rect 9944 9349 9976 9381
rect 9976 9349 10019 9381
rect 9901 9306 10019 9349
rect 10061 9381 10179 9424
rect 10061 9349 10104 9381
rect 10104 9349 10136 9381
rect 10136 9349 10179 9381
rect 10061 9306 10179 9349
rect 10221 9381 10339 9424
rect 10221 9349 10264 9381
rect 10264 9349 10296 9381
rect 10296 9349 10339 9381
rect 10221 9306 10339 9349
rect 10381 9381 10499 9424
rect 10381 9349 10424 9381
rect 10424 9349 10456 9381
rect 10456 9349 10499 9381
rect 10381 9306 10499 9349
rect 10541 9381 10659 9424
rect 10541 9349 10584 9381
rect 10584 9349 10616 9381
rect 10616 9349 10659 9381
rect 10541 9306 10659 9349
rect 10701 9381 10819 9424
rect 10701 9349 10744 9381
rect 10744 9349 10776 9381
rect 10776 9349 10819 9381
rect 10701 9306 10819 9349
rect 10861 9381 10979 9424
rect 10861 9349 10904 9381
rect 10904 9349 10936 9381
rect 10936 9349 10979 9381
rect 10861 9306 10979 9349
rect 11021 9381 11139 9424
rect 11021 9349 11064 9381
rect 11064 9349 11096 9381
rect 11096 9349 11139 9381
rect 11021 9306 11139 9349
rect 11181 9381 11299 9424
rect 11181 9349 11224 9381
rect 11224 9349 11256 9381
rect 11256 9349 11299 9381
rect 11181 9306 11299 9349
rect 11341 9381 11459 9424
rect 11341 9349 11384 9381
rect 11384 9349 11416 9381
rect 11416 9349 11459 9381
rect 11341 9306 11459 9349
rect 11501 9381 11619 9424
rect 11501 9349 11544 9381
rect 11544 9349 11576 9381
rect 11576 9349 11619 9381
rect 11501 9306 11619 9349
rect 11661 9381 11779 9424
rect 11661 9349 11704 9381
rect 11704 9349 11736 9381
rect 11736 9349 11779 9381
rect 11661 9306 11779 9349
rect 11821 9381 11939 9424
rect 11821 9349 11864 9381
rect 11864 9349 11896 9381
rect 11896 9349 11939 9381
rect 11821 9306 11939 9349
rect 11981 9381 12099 9424
rect 11981 9349 12024 9381
rect 12024 9349 12056 9381
rect 12056 9349 12099 9381
rect 11981 9306 12099 9349
rect 12141 9381 12259 9424
rect 12141 9349 12184 9381
rect 12184 9349 12216 9381
rect 12216 9349 12259 9381
rect 12141 9306 12259 9349
rect 12301 9381 12419 9424
rect 12301 9349 12344 9381
rect 12344 9349 12376 9381
rect 12376 9349 12419 9381
rect 12301 9306 12419 9349
rect 12461 9381 12579 9424
rect 12461 9349 12504 9381
rect 12504 9349 12536 9381
rect 12536 9349 12579 9381
rect 12461 9306 12579 9349
rect 12621 9381 12739 9424
rect 12621 9349 12664 9381
rect 12664 9349 12696 9381
rect 12696 9349 12739 9381
rect 12621 9306 12739 9349
rect 9073 9244 9116 9276
rect 9116 9244 9148 9276
rect 9148 9244 9191 9276
rect 9073 9201 9191 9244
rect 12806 9276 12924 9319
rect 12806 9244 12849 9276
rect 12849 9244 12881 9276
rect 12881 9244 12924 9276
rect 9073 9116 9191 9159
rect 9073 9084 9116 9116
rect 9116 9084 9148 9116
rect 9148 9084 9191 9116
rect 9073 9041 9191 9084
rect 9073 8956 9191 8999
rect 9073 8924 9116 8956
rect 9116 8924 9148 8956
rect 9148 8924 9191 8956
rect 9073 8881 9191 8924
rect 9073 8796 9191 8839
rect 9073 8764 9116 8796
rect 9116 8764 9148 8796
rect 9148 8764 9191 8796
rect 9073 8721 9191 8764
rect 9073 8636 9191 8679
rect 9073 8604 9116 8636
rect 9116 8604 9148 8636
rect 9148 8604 9191 8636
rect 9073 8561 9191 8604
rect 9073 8476 9191 8519
rect 9073 8444 9116 8476
rect 9116 8444 9148 8476
rect 9148 8444 9191 8476
rect 9073 8401 9191 8444
rect 9073 8316 9191 8359
rect 9073 8284 9116 8316
rect 9116 8284 9148 8316
rect 9148 8284 9191 8316
rect 9073 8241 9191 8284
rect 9073 8156 9191 8199
rect 9073 8124 9116 8156
rect 9116 8124 9148 8156
rect 9148 8124 9191 8156
rect 9073 8081 9191 8124
rect 9073 7996 9191 8039
rect 9073 7964 9116 7996
rect 9116 7964 9148 7996
rect 9148 7964 9191 7996
rect 9073 7921 9191 7964
rect 9073 7836 9191 7879
rect 9073 7804 9116 7836
rect 9116 7804 9148 7836
rect 9148 7804 9191 7836
rect 9073 7761 9191 7804
rect 9073 7676 9191 7719
rect 9073 7644 9116 7676
rect 9116 7644 9148 7676
rect 9148 7644 9191 7676
rect 9073 7601 9191 7644
rect 9073 7516 9191 7559
rect 9073 7484 9116 7516
rect 9116 7484 9148 7516
rect 9148 7484 9191 7516
rect 9073 7441 9191 7484
rect 9073 7356 9191 7399
rect 9073 7324 9116 7356
rect 9116 7324 9148 7356
rect 9148 7324 9191 7356
rect 9073 7281 9191 7324
rect 9073 7196 9191 7239
rect 9073 7164 9116 7196
rect 9116 7164 9148 7196
rect 9148 7164 9191 7196
rect 9073 7121 9191 7164
rect 9073 7036 9191 7079
rect 9073 7004 9116 7036
rect 9116 7004 9148 7036
rect 9148 7004 9191 7036
rect 9073 6961 9191 7004
rect 9073 6876 9191 6919
rect 9073 6844 9116 6876
rect 9116 6844 9148 6876
rect 9148 6844 9191 6876
rect 9073 6801 9191 6844
rect 9073 6716 9191 6759
rect 9073 6684 9116 6716
rect 9116 6684 9148 6716
rect 9148 6684 9191 6716
rect 9073 6641 9191 6684
rect 9073 6556 9191 6599
rect 9073 6524 9116 6556
rect 9116 6524 9148 6556
rect 9148 6524 9191 6556
rect 9073 6481 9191 6524
rect 9073 6396 9191 6439
rect 9073 6364 9116 6396
rect 9116 6364 9148 6396
rect 9148 6364 9191 6396
rect 9073 6321 9191 6364
rect 9073 6236 9191 6279
rect 9073 6204 9116 6236
rect 9116 6204 9148 6236
rect 9148 6204 9191 6236
rect 9073 6161 9191 6204
rect 9073 6076 9191 6119
rect 9073 6044 9116 6076
rect 9116 6044 9148 6076
rect 9148 6044 9191 6076
rect 9073 6001 9191 6044
rect 9073 5916 9191 5959
rect 9073 5884 9116 5916
rect 9116 5884 9148 5916
rect 9148 5884 9191 5916
rect 9073 5841 9191 5884
rect 9073 5756 9191 5799
rect 12806 9201 12924 9244
rect 12806 9116 12924 9159
rect 12806 9084 12849 9116
rect 12849 9084 12881 9116
rect 12881 9084 12924 9116
rect 12806 9041 12924 9084
rect 12806 8956 12924 8999
rect 12806 8924 12849 8956
rect 12849 8924 12881 8956
rect 12881 8924 12924 8956
rect 12806 8881 12924 8924
rect 12806 8796 12924 8839
rect 12806 8764 12849 8796
rect 12849 8764 12881 8796
rect 12881 8764 12924 8796
rect 12806 8721 12924 8764
rect 12806 8636 12924 8679
rect 12806 8604 12849 8636
rect 12849 8604 12881 8636
rect 12881 8604 12924 8636
rect 12806 8561 12924 8604
rect 12806 8476 12924 8519
rect 12806 8444 12849 8476
rect 12849 8444 12881 8476
rect 12881 8444 12924 8476
rect 12806 8401 12924 8444
rect 12806 8316 12924 8359
rect 12806 8284 12849 8316
rect 12849 8284 12881 8316
rect 12881 8284 12924 8316
rect 12806 8241 12924 8284
rect 12806 8156 12924 8199
rect 12806 8124 12849 8156
rect 12849 8124 12881 8156
rect 12881 8124 12924 8156
rect 12806 8081 12924 8124
rect 12806 7996 12924 8039
rect 12806 7964 12849 7996
rect 12849 7964 12881 7996
rect 12881 7964 12924 7996
rect 12806 7921 12924 7964
rect 12806 7836 12924 7879
rect 12806 7804 12849 7836
rect 12849 7804 12881 7836
rect 12881 7804 12924 7836
rect 12806 7761 12924 7804
rect 12806 7676 12924 7719
rect 12806 7644 12849 7676
rect 12849 7644 12881 7676
rect 12881 7644 12924 7676
rect 12806 7601 12924 7644
rect 12806 7516 12924 7559
rect 12806 7484 12849 7516
rect 12849 7484 12881 7516
rect 12881 7484 12924 7516
rect 12806 7441 12924 7484
rect 12806 7356 12924 7399
rect 12806 7324 12849 7356
rect 12849 7324 12881 7356
rect 12881 7324 12924 7356
rect 12806 7281 12924 7324
rect 12806 7196 12924 7239
rect 12806 7164 12849 7196
rect 12849 7164 12881 7196
rect 12881 7164 12924 7196
rect 12806 7121 12924 7164
rect 12806 7036 12924 7079
rect 12806 7004 12849 7036
rect 12849 7004 12881 7036
rect 12881 7004 12924 7036
rect 12806 6961 12924 7004
rect 12806 6876 12924 6919
rect 12806 6844 12849 6876
rect 12849 6844 12881 6876
rect 12881 6844 12924 6876
rect 12806 6801 12924 6844
rect 12806 6716 12924 6759
rect 12806 6684 12849 6716
rect 12849 6684 12881 6716
rect 12881 6684 12924 6716
rect 12806 6641 12924 6684
rect 12806 6556 12924 6599
rect 12806 6524 12849 6556
rect 12849 6524 12881 6556
rect 12881 6524 12924 6556
rect 12806 6481 12924 6524
rect 12806 6396 12924 6439
rect 12806 6364 12849 6396
rect 12849 6364 12881 6396
rect 12881 6364 12924 6396
rect 12806 6321 12924 6364
rect 12806 6236 12924 6279
rect 12806 6204 12849 6236
rect 12849 6204 12881 6236
rect 12881 6204 12924 6236
rect 12806 6161 12924 6204
rect 12806 6076 12924 6119
rect 12806 6044 12849 6076
rect 12849 6044 12881 6076
rect 12881 6044 12924 6076
rect 12806 6001 12924 6044
rect 12806 5916 12924 5959
rect 12806 5884 12849 5916
rect 12849 5884 12881 5916
rect 12881 5884 12924 5916
rect 12806 5841 12924 5884
rect 9073 5724 9116 5756
rect 9116 5724 9148 5756
rect 9148 5724 9191 5756
rect 9073 5681 9191 5724
rect 12806 5756 12924 5799
rect 12806 5724 12849 5756
rect 12849 5724 12881 5756
rect 12881 5724 12924 5756
rect 9261 5653 9379 5696
rect 9261 5621 9304 5653
rect 9304 5621 9336 5653
rect 9336 5621 9379 5653
rect 9261 5578 9379 5621
rect 9421 5653 9539 5696
rect 9421 5621 9464 5653
rect 9464 5621 9496 5653
rect 9496 5621 9539 5653
rect 9421 5578 9539 5621
rect 9581 5653 9699 5696
rect 9581 5621 9624 5653
rect 9624 5621 9656 5653
rect 9656 5621 9699 5653
rect 9581 5578 9699 5621
rect 9741 5653 9859 5696
rect 9741 5621 9784 5653
rect 9784 5621 9816 5653
rect 9816 5621 9859 5653
rect 9741 5578 9859 5621
rect 9901 5653 10019 5696
rect 9901 5621 9944 5653
rect 9944 5621 9976 5653
rect 9976 5621 10019 5653
rect 9901 5578 10019 5621
rect 10061 5653 10179 5696
rect 10061 5621 10104 5653
rect 10104 5621 10136 5653
rect 10136 5621 10179 5653
rect 10061 5578 10179 5621
rect 10221 5653 10339 5696
rect 10221 5621 10264 5653
rect 10264 5621 10296 5653
rect 10296 5621 10339 5653
rect 10221 5578 10339 5621
rect 10381 5653 10499 5696
rect 10381 5621 10424 5653
rect 10424 5621 10456 5653
rect 10456 5621 10499 5653
rect 10381 5578 10499 5621
rect 10541 5653 10659 5696
rect 10541 5621 10584 5653
rect 10584 5621 10616 5653
rect 10616 5621 10659 5653
rect 10541 5578 10659 5621
rect 10701 5653 10819 5696
rect 10701 5621 10744 5653
rect 10744 5621 10776 5653
rect 10776 5621 10819 5653
rect 10701 5578 10819 5621
rect 10861 5653 10979 5696
rect 10861 5621 10904 5653
rect 10904 5621 10936 5653
rect 10936 5621 10979 5653
rect 10861 5578 10979 5621
rect 11021 5653 11139 5696
rect 11021 5621 11064 5653
rect 11064 5621 11096 5653
rect 11096 5621 11139 5653
rect 11021 5578 11139 5621
rect 11181 5653 11299 5696
rect 11181 5621 11224 5653
rect 11224 5621 11256 5653
rect 11256 5621 11299 5653
rect 11181 5578 11299 5621
rect 11341 5653 11459 5696
rect 11341 5621 11384 5653
rect 11384 5621 11416 5653
rect 11416 5621 11459 5653
rect 11341 5578 11459 5621
rect 11501 5653 11619 5696
rect 11501 5621 11544 5653
rect 11544 5621 11576 5653
rect 11576 5621 11619 5653
rect 11501 5578 11619 5621
rect 11661 5653 11779 5696
rect 11661 5621 11704 5653
rect 11704 5621 11736 5653
rect 11736 5621 11779 5653
rect 11661 5578 11779 5621
rect 11821 5653 11939 5696
rect 11821 5621 11864 5653
rect 11864 5621 11896 5653
rect 11896 5621 11939 5653
rect 11821 5578 11939 5621
rect 11981 5653 12099 5696
rect 11981 5621 12024 5653
rect 12024 5621 12056 5653
rect 12056 5621 12099 5653
rect 11981 5578 12099 5621
rect 12141 5653 12259 5696
rect 12141 5621 12184 5653
rect 12184 5621 12216 5653
rect 12216 5621 12259 5653
rect 12141 5578 12259 5621
rect 12301 5653 12419 5696
rect 12301 5621 12344 5653
rect 12344 5621 12376 5653
rect 12376 5621 12419 5653
rect 12301 5578 12419 5621
rect 12461 5653 12579 5696
rect 12461 5621 12504 5653
rect 12504 5621 12536 5653
rect 12536 5621 12579 5653
rect 12461 5578 12579 5621
rect 12621 5653 12739 5696
rect 12806 5681 12924 5724
rect 12621 5621 12664 5653
rect 12664 5621 12696 5653
rect 12696 5621 12739 5653
rect 12621 5578 12739 5621
rect 15261 9381 15379 9424
rect 15261 9349 15304 9381
rect 15304 9349 15336 9381
rect 15336 9349 15379 9381
rect 15073 9276 15191 9319
rect 15261 9306 15379 9349
rect 15421 9381 15539 9424
rect 15421 9349 15464 9381
rect 15464 9349 15496 9381
rect 15496 9349 15539 9381
rect 15421 9306 15539 9349
rect 15581 9381 15699 9424
rect 15581 9349 15624 9381
rect 15624 9349 15656 9381
rect 15656 9349 15699 9381
rect 15581 9306 15699 9349
rect 15741 9381 15859 9424
rect 15741 9349 15784 9381
rect 15784 9349 15816 9381
rect 15816 9349 15859 9381
rect 15741 9306 15859 9349
rect 15901 9381 16019 9424
rect 15901 9349 15944 9381
rect 15944 9349 15976 9381
rect 15976 9349 16019 9381
rect 15901 9306 16019 9349
rect 16061 9381 16179 9424
rect 16061 9349 16104 9381
rect 16104 9349 16136 9381
rect 16136 9349 16179 9381
rect 16061 9306 16179 9349
rect 16221 9381 16339 9424
rect 16221 9349 16264 9381
rect 16264 9349 16296 9381
rect 16296 9349 16339 9381
rect 16221 9306 16339 9349
rect 16381 9381 16499 9424
rect 16381 9349 16424 9381
rect 16424 9349 16456 9381
rect 16456 9349 16499 9381
rect 16381 9306 16499 9349
rect 16541 9381 16659 9424
rect 16541 9349 16584 9381
rect 16584 9349 16616 9381
rect 16616 9349 16659 9381
rect 16541 9306 16659 9349
rect 16701 9381 16819 9424
rect 16701 9349 16744 9381
rect 16744 9349 16776 9381
rect 16776 9349 16819 9381
rect 16701 9306 16819 9349
rect 16861 9381 16979 9424
rect 16861 9349 16904 9381
rect 16904 9349 16936 9381
rect 16936 9349 16979 9381
rect 16861 9306 16979 9349
rect 17021 9381 17139 9424
rect 17021 9349 17064 9381
rect 17064 9349 17096 9381
rect 17096 9349 17139 9381
rect 17021 9306 17139 9349
rect 17181 9381 17299 9424
rect 17181 9349 17224 9381
rect 17224 9349 17256 9381
rect 17256 9349 17299 9381
rect 17181 9306 17299 9349
rect 17341 9381 17459 9424
rect 17341 9349 17384 9381
rect 17384 9349 17416 9381
rect 17416 9349 17459 9381
rect 17341 9306 17459 9349
rect 17501 9381 17619 9424
rect 17501 9349 17544 9381
rect 17544 9349 17576 9381
rect 17576 9349 17619 9381
rect 17501 9306 17619 9349
rect 17661 9381 17779 9424
rect 17661 9349 17704 9381
rect 17704 9349 17736 9381
rect 17736 9349 17779 9381
rect 17661 9306 17779 9349
rect 17821 9381 17939 9424
rect 17821 9349 17864 9381
rect 17864 9349 17896 9381
rect 17896 9349 17939 9381
rect 17821 9306 17939 9349
rect 17981 9381 18099 9424
rect 17981 9349 18024 9381
rect 18024 9349 18056 9381
rect 18056 9349 18099 9381
rect 17981 9306 18099 9349
rect 18141 9381 18259 9424
rect 18141 9349 18184 9381
rect 18184 9349 18216 9381
rect 18216 9349 18259 9381
rect 18141 9306 18259 9349
rect 18301 9381 18419 9424
rect 18301 9349 18344 9381
rect 18344 9349 18376 9381
rect 18376 9349 18419 9381
rect 18301 9306 18419 9349
rect 18461 9381 18579 9424
rect 18461 9349 18504 9381
rect 18504 9349 18536 9381
rect 18536 9349 18579 9381
rect 18461 9306 18579 9349
rect 18621 9381 18739 9424
rect 18621 9349 18664 9381
rect 18664 9349 18696 9381
rect 18696 9349 18739 9381
rect 18621 9306 18739 9349
rect 15073 9244 15116 9276
rect 15116 9244 15148 9276
rect 15148 9244 15191 9276
rect 15073 9201 15191 9244
rect 18806 9276 18924 9319
rect 18806 9244 18849 9276
rect 18849 9244 18881 9276
rect 18881 9244 18924 9276
rect 15073 9116 15191 9159
rect 15073 9084 15116 9116
rect 15116 9084 15148 9116
rect 15148 9084 15191 9116
rect 15073 9041 15191 9084
rect 15073 8956 15191 8999
rect 15073 8924 15116 8956
rect 15116 8924 15148 8956
rect 15148 8924 15191 8956
rect 15073 8881 15191 8924
rect 15073 8796 15191 8839
rect 15073 8764 15116 8796
rect 15116 8764 15148 8796
rect 15148 8764 15191 8796
rect 15073 8721 15191 8764
rect 15073 8636 15191 8679
rect 15073 8604 15116 8636
rect 15116 8604 15148 8636
rect 15148 8604 15191 8636
rect 15073 8561 15191 8604
rect 15073 8476 15191 8519
rect 15073 8444 15116 8476
rect 15116 8444 15148 8476
rect 15148 8444 15191 8476
rect 15073 8401 15191 8444
rect 15073 8316 15191 8359
rect 15073 8284 15116 8316
rect 15116 8284 15148 8316
rect 15148 8284 15191 8316
rect 15073 8241 15191 8284
rect 15073 8156 15191 8199
rect 15073 8124 15116 8156
rect 15116 8124 15148 8156
rect 15148 8124 15191 8156
rect 15073 8081 15191 8124
rect 15073 7996 15191 8039
rect 15073 7964 15116 7996
rect 15116 7964 15148 7996
rect 15148 7964 15191 7996
rect 15073 7921 15191 7964
rect 15073 7836 15191 7879
rect 15073 7804 15116 7836
rect 15116 7804 15148 7836
rect 15148 7804 15191 7836
rect 15073 7761 15191 7804
rect 15073 7676 15191 7719
rect 15073 7644 15116 7676
rect 15116 7644 15148 7676
rect 15148 7644 15191 7676
rect 15073 7601 15191 7644
rect 15073 7516 15191 7559
rect 15073 7484 15116 7516
rect 15116 7484 15148 7516
rect 15148 7484 15191 7516
rect 15073 7441 15191 7484
rect 15073 7356 15191 7399
rect 15073 7324 15116 7356
rect 15116 7324 15148 7356
rect 15148 7324 15191 7356
rect 15073 7281 15191 7324
rect 15073 7196 15191 7239
rect 15073 7164 15116 7196
rect 15116 7164 15148 7196
rect 15148 7164 15191 7196
rect 15073 7121 15191 7164
rect 15073 7036 15191 7079
rect 15073 7004 15116 7036
rect 15116 7004 15148 7036
rect 15148 7004 15191 7036
rect 15073 6961 15191 7004
rect 15073 6876 15191 6919
rect 15073 6844 15116 6876
rect 15116 6844 15148 6876
rect 15148 6844 15191 6876
rect 15073 6801 15191 6844
rect 15073 6716 15191 6759
rect 15073 6684 15116 6716
rect 15116 6684 15148 6716
rect 15148 6684 15191 6716
rect 15073 6641 15191 6684
rect 15073 6556 15191 6599
rect 15073 6524 15116 6556
rect 15116 6524 15148 6556
rect 15148 6524 15191 6556
rect 15073 6481 15191 6524
rect 15073 6396 15191 6439
rect 15073 6364 15116 6396
rect 15116 6364 15148 6396
rect 15148 6364 15191 6396
rect 15073 6321 15191 6364
rect 15073 6236 15191 6279
rect 15073 6204 15116 6236
rect 15116 6204 15148 6236
rect 15148 6204 15191 6236
rect 15073 6161 15191 6204
rect 15073 6076 15191 6119
rect 15073 6044 15116 6076
rect 15116 6044 15148 6076
rect 15148 6044 15191 6076
rect 15073 6001 15191 6044
rect 15073 5916 15191 5959
rect 15073 5884 15116 5916
rect 15116 5884 15148 5916
rect 15148 5884 15191 5916
rect 15073 5841 15191 5884
rect 15073 5756 15191 5799
rect 18806 9201 18924 9244
rect 18806 9116 18924 9159
rect 18806 9084 18849 9116
rect 18849 9084 18881 9116
rect 18881 9084 18924 9116
rect 18806 9041 18924 9084
rect 18806 8956 18924 8999
rect 18806 8924 18849 8956
rect 18849 8924 18881 8956
rect 18881 8924 18924 8956
rect 18806 8881 18924 8924
rect 18806 8796 18924 8839
rect 18806 8764 18849 8796
rect 18849 8764 18881 8796
rect 18881 8764 18924 8796
rect 18806 8721 18924 8764
rect 18806 8636 18924 8679
rect 18806 8604 18849 8636
rect 18849 8604 18881 8636
rect 18881 8604 18924 8636
rect 18806 8561 18924 8604
rect 18806 8476 18924 8519
rect 18806 8444 18849 8476
rect 18849 8444 18881 8476
rect 18881 8444 18924 8476
rect 18806 8401 18924 8444
rect 18806 8316 18924 8359
rect 18806 8284 18849 8316
rect 18849 8284 18881 8316
rect 18881 8284 18924 8316
rect 18806 8241 18924 8284
rect 18806 8156 18924 8199
rect 18806 8124 18849 8156
rect 18849 8124 18881 8156
rect 18881 8124 18924 8156
rect 18806 8081 18924 8124
rect 18806 7996 18924 8039
rect 18806 7964 18849 7996
rect 18849 7964 18881 7996
rect 18881 7964 18924 7996
rect 18806 7921 18924 7964
rect 18806 7836 18924 7879
rect 18806 7804 18849 7836
rect 18849 7804 18881 7836
rect 18881 7804 18924 7836
rect 18806 7761 18924 7804
rect 18806 7676 18924 7719
rect 18806 7644 18849 7676
rect 18849 7644 18881 7676
rect 18881 7644 18924 7676
rect 18806 7601 18924 7644
rect 18806 7516 18924 7559
rect 18806 7484 18849 7516
rect 18849 7484 18881 7516
rect 18881 7484 18924 7516
rect 18806 7441 18924 7484
rect 18806 7356 18924 7399
rect 18806 7324 18849 7356
rect 18849 7324 18881 7356
rect 18881 7324 18924 7356
rect 18806 7281 18924 7324
rect 18806 7196 18924 7239
rect 18806 7164 18849 7196
rect 18849 7164 18881 7196
rect 18881 7164 18924 7196
rect 18806 7121 18924 7164
rect 18806 7036 18924 7079
rect 18806 7004 18849 7036
rect 18849 7004 18881 7036
rect 18881 7004 18924 7036
rect 18806 6961 18924 7004
rect 18806 6876 18924 6919
rect 18806 6844 18849 6876
rect 18849 6844 18881 6876
rect 18881 6844 18924 6876
rect 18806 6801 18924 6844
rect 18806 6716 18924 6759
rect 18806 6684 18849 6716
rect 18849 6684 18881 6716
rect 18881 6684 18924 6716
rect 18806 6641 18924 6684
rect 18806 6556 18924 6599
rect 18806 6524 18849 6556
rect 18849 6524 18881 6556
rect 18881 6524 18924 6556
rect 18806 6481 18924 6524
rect 18806 6396 18924 6439
rect 18806 6364 18849 6396
rect 18849 6364 18881 6396
rect 18881 6364 18924 6396
rect 18806 6321 18924 6364
rect 18806 6236 18924 6279
rect 18806 6204 18849 6236
rect 18849 6204 18881 6236
rect 18881 6204 18924 6236
rect 18806 6161 18924 6204
rect 18806 6076 18924 6119
rect 18806 6044 18849 6076
rect 18849 6044 18881 6076
rect 18881 6044 18924 6076
rect 18806 6001 18924 6044
rect 18806 5916 18924 5959
rect 18806 5884 18849 5916
rect 18849 5884 18881 5916
rect 18881 5884 18924 5916
rect 18806 5841 18924 5884
rect 15073 5724 15116 5756
rect 15116 5724 15148 5756
rect 15148 5724 15191 5756
rect 15073 5681 15191 5724
rect 18806 5756 18924 5799
rect 18806 5724 18849 5756
rect 18849 5724 18881 5756
rect 18881 5724 18924 5756
rect 15261 5653 15379 5696
rect 15261 5621 15304 5653
rect 15304 5621 15336 5653
rect 15336 5621 15379 5653
rect 15261 5578 15379 5621
rect 15421 5653 15539 5696
rect 15421 5621 15464 5653
rect 15464 5621 15496 5653
rect 15496 5621 15539 5653
rect 15421 5578 15539 5621
rect 15581 5653 15699 5696
rect 15581 5621 15624 5653
rect 15624 5621 15656 5653
rect 15656 5621 15699 5653
rect 15581 5578 15699 5621
rect 15741 5653 15859 5696
rect 15741 5621 15784 5653
rect 15784 5621 15816 5653
rect 15816 5621 15859 5653
rect 15741 5578 15859 5621
rect 15901 5653 16019 5696
rect 15901 5621 15944 5653
rect 15944 5621 15976 5653
rect 15976 5621 16019 5653
rect 15901 5578 16019 5621
rect 16061 5653 16179 5696
rect 16061 5621 16104 5653
rect 16104 5621 16136 5653
rect 16136 5621 16179 5653
rect 16061 5578 16179 5621
rect 16221 5653 16339 5696
rect 16221 5621 16264 5653
rect 16264 5621 16296 5653
rect 16296 5621 16339 5653
rect 16221 5578 16339 5621
rect 16381 5653 16499 5696
rect 16381 5621 16424 5653
rect 16424 5621 16456 5653
rect 16456 5621 16499 5653
rect 16381 5578 16499 5621
rect 16541 5653 16659 5696
rect 16541 5621 16584 5653
rect 16584 5621 16616 5653
rect 16616 5621 16659 5653
rect 16541 5578 16659 5621
rect 16701 5653 16819 5696
rect 16701 5621 16744 5653
rect 16744 5621 16776 5653
rect 16776 5621 16819 5653
rect 16701 5578 16819 5621
rect 16861 5653 16979 5696
rect 16861 5621 16904 5653
rect 16904 5621 16936 5653
rect 16936 5621 16979 5653
rect 16861 5578 16979 5621
rect 17021 5653 17139 5696
rect 17021 5621 17064 5653
rect 17064 5621 17096 5653
rect 17096 5621 17139 5653
rect 17021 5578 17139 5621
rect 17181 5653 17299 5696
rect 17181 5621 17224 5653
rect 17224 5621 17256 5653
rect 17256 5621 17299 5653
rect 17181 5578 17299 5621
rect 17341 5653 17459 5696
rect 17341 5621 17384 5653
rect 17384 5621 17416 5653
rect 17416 5621 17459 5653
rect 17341 5578 17459 5621
rect 17501 5653 17619 5696
rect 17501 5621 17544 5653
rect 17544 5621 17576 5653
rect 17576 5621 17619 5653
rect 17501 5578 17619 5621
rect 17661 5653 17779 5696
rect 17661 5621 17704 5653
rect 17704 5621 17736 5653
rect 17736 5621 17779 5653
rect 17661 5578 17779 5621
rect 17821 5653 17939 5696
rect 17821 5621 17864 5653
rect 17864 5621 17896 5653
rect 17896 5621 17939 5653
rect 17821 5578 17939 5621
rect 17981 5653 18099 5696
rect 17981 5621 18024 5653
rect 18024 5621 18056 5653
rect 18056 5621 18099 5653
rect 17981 5578 18099 5621
rect 18141 5653 18259 5696
rect 18141 5621 18184 5653
rect 18184 5621 18216 5653
rect 18216 5621 18259 5653
rect 18141 5578 18259 5621
rect 18301 5653 18419 5696
rect 18301 5621 18344 5653
rect 18344 5621 18376 5653
rect 18376 5621 18419 5653
rect 18301 5578 18419 5621
rect 18461 5653 18579 5696
rect 18461 5621 18504 5653
rect 18504 5621 18536 5653
rect 18536 5621 18579 5653
rect 18461 5578 18579 5621
rect 18621 5653 18739 5696
rect 18806 5681 18924 5724
rect 18621 5621 18664 5653
rect 18664 5621 18696 5653
rect 18696 5621 18739 5653
rect 18621 5578 18739 5621
rect 21261 9381 21379 9424
rect 21261 9349 21304 9381
rect 21304 9349 21336 9381
rect 21336 9349 21379 9381
rect 21073 9276 21191 9319
rect 21261 9306 21379 9349
rect 21421 9381 21539 9424
rect 21421 9349 21464 9381
rect 21464 9349 21496 9381
rect 21496 9349 21539 9381
rect 21421 9306 21539 9349
rect 21581 9381 21699 9424
rect 21581 9349 21624 9381
rect 21624 9349 21656 9381
rect 21656 9349 21699 9381
rect 21581 9306 21699 9349
rect 21741 9381 21859 9424
rect 21741 9349 21784 9381
rect 21784 9349 21816 9381
rect 21816 9349 21859 9381
rect 21741 9306 21859 9349
rect 21901 9381 22019 9424
rect 21901 9349 21944 9381
rect 21944 9349 21976 9381
rect 21976 9349 22019 9381
rect 21901 9306 22019 9349
rect 22061 9381 22179 9424
rect 22061 9349 22104 9381
rect 22104 9349 22136 9381
rect 22136 9349 22179 9381
rect 22061 9306 22179 9349
rect 22221 9381 22339 9424
rect 22221 9349 22264 9381
rect 22264 9349 22296 9381
rect 22296 9349 22339 9381
rect 22221 9306 22339 9349
rect 22381 9381 22499 9424
rect 22381 9349 22424 9381
rect 22424 9349 22456 9381
rect 22456 9349 22499 9381
rect 22381 9306 22499 9349
rect 22541 9381 22659 9424
rect 22541 9349 22584 9381
rect 22584 9349 22616 9381
rect 22616 9349 22659 9381
rect 22541 9306 22659 9349
rect 22701 9381 22819 9424
rect 22701 9349 22744 9381
rect 22744 9349 22776 9381
rect 22776 9349 22819 9381
rect 22701 9306 22819 9349
rect 22861 9381 22979 9424
rect 22861 9349 22904 9381
rect 22904 9349 22936 9381
rect 22936 9349 22979 9381
rect 22861 9306 22979 9349
rect 23021 9381 23139 9424
rect 23021 9349 23064 9381
rect 23064 9349 23096 9381
rect 23096 9349 23139 9381
rect 23021 9306 23139 9349
rect 23181 9381 23299 9424
rect 23181 9349 23224 9381
rect 23224 9349 23256 9381
rect 23256 9349 23299 9381
rect 23181 9306 23299 9349
rect 23341 9381 23459 9424
rect 23341 9349 23384 9381
rect 23384 9349 23416 9381
rect 23416 9349 23459 9381
rect 23341 9306 23459 9349
rect 23501 9381 23619 9424
rect 23501 9349 23544 9381
rect 23544 9349 23576 9381
rect 23576 9349 23619 9381
rect 23501 9306 23619 9349
rect 23661 9381 23779 9424
rect 23661 9349 23704 9381
rect 23704 9349 23736 9381
rect 23736 9349 23779 9381
rect 23661 9306 23779 9349
rect 23821 9381 23939 9424
rect 23821 9349 23864 9381
rect 23864 9349 23896 9381
rect 23896 9349 23939 9381
rect 23821 9306 23939 9349
rect 23981 9381 24099 9424
rect 23981 9349 24024 9381
rect 24024 9349 24056 9381
rect 24056 9349 24099 9381
rect 23981 9306 24099 9349
rect 24141 9381 24259 9424
rect 24141 9349 24184 9381
rect 24184 9349 24216 9381
rect 24216 9349 24259 9381
rect 24141 9306 24259 9349
rect 24301 9381 24419 9424
rect 24301 9349 24344 9381
rect 24344 9349 24376 9381
rect 24376 9349 24419 9381
rect 24301 9306 24419 9349
rect 24461 9381 24579 9424
rect 24461 9349 24504 9381
rect 24504 9349 24536 9381
rect 24536 9349 24579 9381
rect 24461 9306 24579 9349
rect 24621 9381 24739 9424
rect 24621 9349 24664 9381
rect 24664 9349 24696 9381
rect 24696 9349 24739 9381
rect 24621 9306 24739 9349
rect 21073 9244 21116 9276
rect 21116 9244 21148 9276
rect 21148 9244 21191 9276
rect 21073 9201 21191 9244
rect 24806 9276 24924 9319
rect 24806 9244 24849 9276
rect 24849 9244 24881 9276
rect 24881 9244 24924 9276
rect 21073 9116 21191 9159
rect 21073 9084 21116 9116
rect 21116 9084 21148 9116
rect 21148 9084 21191 9116
rect 21073 9041 21191 9084
rect 21073 8956 21191 8999
rect 21073 8924 21116 8956
rect 21116 8924 21148 8956
rect 21148 8924 21191 8956
rect 21073 8881 21191 8924
rect 21073 8796 21191 8839
rect 21073 8764 21116 8796
rect 21116 8764 21148 8796
rect 21148 8764 21191 8796
rect 21073 8721 21191 8764
rect 21073 8636 21191 8679
rect 21073 8604 21116 8636
rect 21116 8604 21148 8636
rect 21148 8604 21191 8636
rect 21073 8561 21191 8604
rect 21073 8476 21191 8519
rect 21073 8444 21116 8476
rect 21116 8444 21148 8476
rect 21148 8444 21191 8476
rect 21073 8401 21191 8444
rect 21073 8316 21191 8359
rect 21073 8284 21116 8316
rect 21116 8284 21148 8316
rect 21148 8284 21191 8316
rect 21073 8241 21191 8284
rect 21073 8156 21191 8199
rect 21073 8124 21116 8156
rect 21116 8124 21148 8156
rect 21148 8124 21191 8156
rect 21073 8081 21191 8124
rect 21073 7996 21191 8039
rect 21073 7964 21116 7996
rect 21116 7964 21148 7996
rect 21148 7964 21191 7996
rect 21073 7921 21191 7964
rect 21073 7836 21191 7879
rect 21073 7804 21116 7836
rect 21116 7804 21148 7836
rect 21148 7804 21191 7836
rect 21073 7761 21191 7804
rect 21073 7676 21191 7719
rect 21073 7644 21116 7676
rect 21116 7644 21148 7676
rect 21148 7644 21191 7676
rect 21073 7601 21191 7644
rect 21073 7516 21191 7559
rect 21073 7484 21116 7516
rect 21116 7484 21148 7516
rect 21148 7484 21191 7516
rect 21073 7441 21191 7484
rect 21073 7356 21191 7399
rect 21073 7324 21116 7356
rect 21116 7324 21148 7356
rect 21148 7324 21191 7356
rect 21073 7281 21191 7324
rect 21073 7196 21191 7239
rect 21073 7164 21116 7196
rect 21116 7164 21148 7196
rect 21148 7164 21191 7196
rect 21073 7121 21191 7164
rect 21073 7036 21191 7079
rect 21073 7004 21116 7036
rect 21116 7004 21148 7036
rect 21148 7004 21191 7036
rect 21073 6961 21191 7004
rect 21073 6876 21191 6919
rect 21073 6844 21116 6876
rect 21116 6844 21148 6876
rect 21148 6844 21191 6876
rect 21073 6801 21191 6844
rect 21073 6716 21191 6759
rect 21073 6684 21116 6716
rect 21116 6684 21148 6716
rect 21148 6684 21191 6716
rect 21073 6641 21191 6684
rect 21073 6556 21191 6599
rect 21073 6524 21116 6556
rect 21116 6524 21148 6556
rect 21148 6524 21191 6556
rect 21073 6481 21191 6524
rect 21073 6396 21191 6439
rect 21073 6364 21116 6396
rect 21116 6364 21148 6396
rect 21148 6364 21191 6396
rect 21073 6321 21191 6364
rect 21073 6236 21191 6279
rect 21073 6204 21116 6236
rect 21116 6204 21148 6236
rect 21148 6204 21191 6236
rect 21073 6161 21191 6204
rect 21073 6076 21191 6119
rect 21073 6044 21116 6076
rect 21116 6044 21148 6076
rect 21148 6044 21191 6076
rect 21073 6001 21191 6044
rect 21073 5916 21191 5959
rect 21073 5884 21116 5916
rect 21116 5884 21148 5916
rect 21148 5884 21191 5916
rect 21073 5841 21191 5884
rect 21073 5756 21191 5799
rect 24806 9201 24924 9244
rect 24806 9116 24924 9159
rect 24806 9084 24849 9116
rect 24849 9084 24881 9116
rect 24881 9084 24924 9116
rect 24806 9041 24924 9084
rect 24806 8956 24924 8999
rect 24806 8924 24849 8956
rect 24849 8924 24881 8956
rect 24881 8924 24924 8956
rect 24806 8881 24924 8924
rect 24806 8796 24924 8839
rect 24806 8764 24849 8796
rect 24849 8764 24881 8796
rect 24881 8764 24924 8796
rect 24806 8721 24924 8764
rect 24806 8636 24924 8679
rect 24806 8604 24849 8636
rect 24849 8604 24881 8636
rect 24881 8604 24924 8636
rect 24806 8561 24924 8604
rect 24806 8476 24924 8519
rect 24806 8444 24849 8476
rect 24849 8444 24881 8476
rect 24881 8444 24924 8476
rect 24806 8401 24924 8444
rect 24806 8316 24924 8359
rect 24806 8284 24849 8316
rect 24849 8284 24881 8316
rect 24881 8284 24924 8316
rect 24806 8241 24924 8284
rect 24806 8156 24924 8199
rect 24806 8124 24849 8156
rect 24849 8124 24881 8156
rect 24881 8124 24924 8156
rect 24806 8081 24924 8124
rect 24806 7996 24924 8039
rect 24806 7964 24849 7996
rect 24849 7964 24881 7996
rect 24881 7964 24924 7996
rect 24806 7921 24924 7964
rect 24806 7836 24924 7879
rect 24806 7804 24849 7836
rect 24849 7804 24881 7836
rect 24881 7804 24924 7836
rect 24806 7761 24924 7804
rect 24806 7676 24924 7719
rect 24806 7644 24849 7676
rect 24849 7644 24881 7676
rect 24881 7644 24924 7676
rect 24806 7601 24924 7644
rect 24806 7516 24924 7559
rect 24806 7484 24849 7516
rect 24849 7484 24881 7516
rect 24881 7484 24924 7516
rect 24806 7441 24924 7484
rect 24806 7356 24924 7399
rect 24806 7324 24849 7356
rect 24849 7324 24881 7356
rect 24881 7324 24924 7356
rect 24806 7281 24924 7324
rect 24806 7196 24924 7239
rect 24806 7164 24849 7196
rect 24849 7164 24881 7196
rect 24881 7164 24924 7196
rect 24806 7121 24924 7164
rect 24806 7036 24924 7079
rect 24806 7004 24849 7036
rect 24849 7004 24881 7036
rect 24881 7004 24924 7036
rect 24806 6961 24924 7004
rect 24806 6876 24924 6919
rect 24806 6844 24849 6876
rect 24849 6844 24881 6876
rect 24881 6844 24924 6876
rect 24806 6801 24924 6844
rect 24806 6716 24924 6759
rect 24806 6684 24849 6716
rect 24849 6684 24881 6716
rect 24881 6684 24924 6716
rect 24806 6641 24924 6684
rect 24806 6556 24924 6599
rect 24806 6524 24849 6556
rect 24849 6524 24881 6556
rect 24881 6524 24924 6556
rect 24806 6481 24924 6524
rect 24806 6396 24924 6439
rect 24806 6364 24849 6396
rect 24849 6364 24881 6396
rect 24881 6364 24924 6396
rect 24806 6321 24924 6364
rect 24806 6236 24924 6279
rect 24806 6204 24849 6236
rect 24849 6204 24881 6236
rect 24881 6204 24924 6236
rect 24806 6161 24924 6204
rect 24806 6076 24924 6119
rect 24806 6044 24849 6076
rect 24849 6044 24881 6076
rect 24881 6044 24924 6076
rect 24806 6001 24924 6044
rect 24806 5916 24924 5959
rect 24806 5884 24849 5916
rect 24849 5884 24881 5916
rect 24881 5884 24924 5916
rect 24806 5841 24924 5884
rect 21073 5724 21116 5756
rect 21116 5724 21148 5756
rect 21148 5724 21191 5756
rect 21073 5681 21191 5724
rect 24806 5756 24924 5799
rect 24806 5724 24849 5756
rect 24849 5724 24881 5756
rect 24881 5724 24924 5756
rect 21261 5653 21379 5696
rect 21261 5621 21304 5653
rect 21304 5621 21336 5653
rect 21336 5621 21379 5653
rect 21261 5578 21379 5621
rect 21421 5653 21539 5696
rect 21421 5621 21464 5653
rect 21464 5621 21496 5653
rect 21496 5621 21539 5653
rect 21421 5578 21539 5621
rect 21581 5653 21699 5696
rect 21581 5621 21624 5653
rect 21624 5621 21656 5653
rect 21656 5621 21699 5653
rect 21581 5578 21699 5621
rect 21741 5653 21859 5696
rect 21741 5621 21784 5653
rect 21784 5621 21816 5653
rect 21816 5621 21859 5653
rect 21741 5578 21859 5621
rect 21901 5653 22019 5696
rect 21901 5621 21944 5653
rect 21944 5621 21976 5653
rect 21976 5621 22019 5653
rect 21901 5578 22019 5621
rect 22061 5653 22179 5696
rect 22061 5621 22104 5653
rect 22104 5621 22136 5653
rect 22136 5621 22179 5653
rect 22061 5578 22179 5621
rect 22221 5653 22339 5696
rect 22221 5621 22264 5653
rect 22264 5621 22296 5653
rect 22296 5621 22339 5653
rect 22221 5578 22339 5621
rect 22381 5653 22499 5696
rect 22381 5621 22424 5653
rect 22424 5621 22456 5653
rect 22456 5621 22499 5653
rect 22381 5578 22499 5621
rect 22541 5653 22659 5696
rect 22541 5621 22584 5653
rect 22584 5621 22616 5653
rect 22616 5621 22659 5653
rect 22541 5578 22659 5621
rect 22701 5653 22819 5696
rect 22701 5621 22744 5653
rect 22744 5621 22776 5653
rect 22776 5621 22819 5653
rect 22701 5578 22819 5621
rect 22861 5653 22979 5696
rect 22861 5621 22904 5653
rect 22904 5621 22936 5653
rect 22936 5621 22979 5653
rect 22861 5578 22979 5621
rect 23021 5653 23139 5696
rect 23021 5621 23064 5653
rect 23064 5621 23096 5653
rect 23096 5621 23139 5653
rect 23021 5578 23139 5621
rect 23181 5653 23299 5696
rect 23181 5621 23224 5653
rect 23224 5621 23256 5653
rect 23256 5621 23299 5653
rect 23181 5578 23299 5621
rect 23341 5653 23459 5696
rect 23341 5621 23384 5653
rect 23384 5621 23416 5653
rect 23416 5621 23459 5653
rect 23341 5578 23459 5621
rect 23501 5653 23619 5696
rect 23501 5621 23544 5653
rect 23544 5621 23576 5653
rect 23576 5621 23619 5653
rect 23501 5578 23619 5621
rect 23661 5653 23779 5696
rect 23661 5621 23704 5653
rect 23704 5621 23736 5653
rect 23736 5621 23779 5653
rect 23661 5578 23779 5621
rect 23821 5653 23939 5696
rect 23821 5621 23864 5653
rect 23864 5621 23896 5653
rect 23896 5621 23939 5653
rect 23821 5578 23939 5621
rect 23981 5653 24099 5696
rect 23981 5621 24024 5653
rect 24024 5621 24056 5653
rect 24056 5621 24099 5653
rect 23981 5578 24099 5621
rect 24141 5653 24259 5696
rect 24141 5621 24184 5653
rect 24184 5621 24216 5653
rect 24216 5621 24259 5653
rect 24141 5578 24259 5621
rect 24301 5653 24419 5696
rect 24301 5621 24344 5653
rect 24344 5621 24376 5653
rect 24376 5621 24419 5653
rect 24301 5578 24419 5621
rect 24461 5653 24579 5696
rect 24461 5621 24504 5653
rect 24504 5621 24536 5653
rect 24536 5621 24579 5653
rect 24461 5578 24579 5621
rect 24621 5653 24739 5696
rect 24806 5681 24924 5724
rect 24621 5621 24664 5653
rect 24664 5621 24696 5653
rect 24696 5621 24739 5653
rect 24621 5578 24739 5621
rect 3261 3381 3379 3424
rect 3261 3349 3304 3381
rect 3304 3349 3336 3381
rect 3336 3349 3379 3381
rect 3073 3276 3191 3319
rect 3261 3306 3379 3349
rect 3421 3381 3539 3424
rect 3421 3349 3464 3381
rect 3464 3349 3496 3381
rect 3496 3349 3539 3381
rect 3421 3306 3539 3349
rect 3581 3381 3699 3424
rect 3581 3349 3624 3381
rect 3624 3349 3656 3381
rect 3656 3349 3699 3381
rect 3581 3306 3699 3349
rect 3741 3381 3859 3424
rect 3741 3349 3784 3381
rect 3784 3349 3816 3381
rect 3816 3349 3859 3381
rect 3741 3306 3859 3349
rect 3901 3381 4019 3424
rect 3901 3349 3944 3381
rect 3944 3349 3976 3381
rect 3976 3349 4019 3381
rect 3901 3306 4019 3349
rect 4061 3381 4179 3424
rect 4061 3349 4104 3381
rect 4104 3349 4136 3381
rect 4136 3349 4179 3381
rect 4061 3306 4179 3349
rect 4221 3381 4339 3424
rect 4221 3349 4264 3381
rect 4264 3349 4296 3381
rect 4296 3349 4339 3381
rect 4221 3306 4339 3349
rect 4381 3381 4499 3424
rect 4381 3349 4424 3381
rect 4424 3349 4456 3381
rect 4456 3349 4499 3381
rect 4381 3306 4499 3349
rect 4541 3381 4659 3424
rect 4541 3349 4584 3381
rect 4584 3349 4616 3381
rect 4616 3349 4659 3381
rect 4541 3306 4659 3349
rect 4701 3381 4819 3424
rect 4701 3349 4744 3381
rect 4744 3349 4776 3381
rect 4776 3349 4819 3381
rect 4701 3306 4819 3349
rect 4861 3381 4979 3424
rect 4861 3349 4904 3381
rect 4904 3349 4936 3381
rect 4936 3349 4979 3381
rect 4861 3306 4979 3349
rect 5021 3381 5139 3424
rect 5021 3349 5064 3381
rect 5064 3349 5096 3381
rect 5096 3349 5139 3381
rect 5021 3306 5139 3349
rect 5181 3381 5299 3424
rect 5181 3349 5224 3381
rect 5224 3349 5256 3381
rect 5256 3349 5299 3381
rect 5181 3306 5299 3349
rect 5341 3381 5459 3424
rect 5341 3349 5384 3381
rect 5384 3349 5416 3381
rect 5416 3349 5459 3381
rect 5341 3306 5459 3349
rect 5501 3381 5619 3424
rect 5501 3349 5544 3381
rect 5544 3349 5576 3381
rect 5576 3349 5619 3381
rect 5501 3306 5619 3349
rect 5661 3381 5779 3424
rect 5661 3349 5704 3381
rect 5704 3349 5736 3381
rect 5736 3349 5779 3381
rect 5661 3306 5779 3349
rect 5821 3381 5939 3424
rect 5821 3349 5864 3381
rect 5864 3349 5896 3381
rect 5896 3349 5939 3381
rect 5821 3306 5939 3349
rect 5981 3381 6099 3424
rect 5981 3349 6024 3381
rect 6024 3349 6056 3381
rect 6056 3349 6099 3381
rect 5981 3306 6099 3349
rect 6141 3381 6259 3424
rect 6141 3349 6184 3381
rect 6184 3349 6216 3381
rect 6216 3349 6259 3381
rect 6141 3306 6259 3349
rect 6301 3381 6419 3424
rect 6301 3349 6344 3381
rect 6344 3349 6376 3381
rect 6376 3349 6419 3381
rect 6301 3306 6419 3349
rect 6461 3381 6579 3424
rect 6461 3349 6504 3381
rect 6504 3349 6536 3381
rect 6536 3349 6579 3381
rect 6461 3306 6579 3349
rect 6621 3381 6739 3424
rect 6621 3349 6664 3381
rect 6664 3349 6696 3381
rect 6696 3349 6739 3381
rect 6621 3306 6739 3349
rect 3073 3244 3116 3276
rect 3116 3244 3148 3276
rect 3148 3244 3191 3276
rect 3073 3201 3191 3244
rect 6806 3276 6924 3319
rect 6806 3244 6849 3276
rect 6849 3244 6881 3276
rect 6881 3244 6924 3276
rect 3073 3116 3191 3159
rect 3073 3084 3116 3116
rect 3116 3084 3148 3116
rect 3148 3084 3191 3116
rect 3073 3041 3191 3084
rect 3073 2956 3191 2999
rect 3073 2924 3116 2956
rect 3116 2924 3148 2956
rect 3148 2924 3191 2956
rect 3073 2881 3191 2924
rect 3073 2796 3191 2839
rect 3073 2764 3116 2796
rect 3116 2764 3148 2796
rect 3148 2764 3191 2796
rect 3073 2721 3191 2764
rect 3073 2636 3191 2679
rect 3073 2604 3116 2636
rect 3116 2604 3148 2636
rect 3148 2604 3191 2636
rect 3073 2561 3191 2604
rect 3073 2476 3191 2519
rect 3073 2444 3116 2476
rect 3116 2444 3148 2476
rect 3148 2444 3191 2476
rect 3073 2401 3191 2444
rect 3073 2316 3191 2359
rect 3073 2284 3116 2316
rect 3116 2284 3148 2316
rect 3148 2284 3191 2316
rect 3073 2241 3191 2284
rect 3073 2156 3191 2199
rect 3073 2124 3116 2156
rect 3116 2124 3148 2156
rect 3148 2124 3191 2156
rect 3073 2081 3191 2124
rect 3073 1996 3191 2039
rect 3073 1964 3116 1996
rect 3116 1964 3148 1996
rect 3148 1964 3191 1996
rect 3073 1921 3191 1964
rect 3073 1836 3191 1879
rect 3073 1804 3116 1836
rect 3116 1804 3148 1836
rect 3148 1804 3191 1836
rect 3073 1761 3191 1804
rect 3073 1676 3191 1719
rect 3073 1644 3116 1676
rect 3116 1644 3148 1676
rect 3148 1644 3191 1676
rect 3073 1601 3191 1644
rect 3073 1516 3191 1559
rect 3073 1484 3116 1516
rect 3116 1484 3148 1516
rect 3148 1484 3191 1516
rect 3073 1441 3191 1484
rect 3073 1356 3191 1399
rect 3073 1324 3116 1356
rect 3116 1324 3148 1356
rect 3148 1324 3191 1356
rect 3073 1281 3191 1324
rect 3073 1196 3191 1239
rect 3073 1164 3116 1196
rect 3116 1164 3148 1196
rect 3148 1164 3191 1196
rect 3073 1121 3191 1164
rect 3073 1036 3191 1079
rect 3073 1004 3116 1036
rect 3116 1004 3148 1036
rect 3148 1004 3191 1036
rect 3073 961 3191 1004
rect 3073 876 3191 919
rect 3073 844 3116 876
rect 3116 844 3148 876
rect 3148 844 3191 876
rect 3073 801 3191 844
rect 3073 716 3191 759
rect 3073 684 3116 716
rect 3116 684 3148 716
rect 3148 684 3191 716
rect 3073 641 3191 684
rect 3073 556 3191 599
rect 3073 524 3116 556
rect 3116 524 3148 556
rect 3148 524 3191 556
rect 3073 481 3191 524
rect 3073 396 3191 439
rect 3073 364 3116 396
rect 3116 364 3148 396
rect 3148 364 3191 396
rect 3073 321 3191 364
rect 3073 236 3191 279
rect 3073 204 3116 236
rect 3116 204 3148 236
rect 3148 204 3191 236
rect 3073 161 3191 204
rect 3073 76 3191 119
rect 3073 44 3116 76
rect 3116 44 3148 76
rect 3148 44 3191 76
rect 3073 1 3191 44
rect 3073 -84 3191 -41
rect 3073 -116 3116 -84
rect 3116 -116 3148 -84
rect 3148 -116 3191 -84
rect 3073 -159 3191 -116
rect 3073 -244 3191 -201
rect 6806 3201 6924 3244
rect 6806 3116 6924 3159
rect 6806 3084 6849 3116
rect 6849 3084 6881 3116
rect 6881 3084 6924 3116
rect 6806 3041 6924 3084
rect 6806 2956 6924 2999
rect 6806 2924 6849 2956
rect 6849 2924 6881 2956
rect 6881 2924 6924 2956
rect 6806 2881 6924 2924
rect 6806 2796 6924 2839
rect 6806 2764 6849 2796
rect 6849 2764 6881 2796
rect 6881 2764 6924 2796
rect 6806 2721 6924 2764
rect 6806 2636 6924 2679
rect 6806 2604 6849 2636
rect 6849 2604 6881 2636
rect 6881 2604 6924 2636
rect 6806 2561 6924 2604
rect 6806 2476 6924 2519
rect 6806 2444 6849 2476
rect 6849 2444 6881 2476
rect 6881 2444 6924 2476
rect 6806 2401 6924 2444
rect 6806 2316 6924 2359
rect 6806 2284 6849 2316
rect 6849 2284 6881 2316
rect 6881 2284 6924 2316
rect 6806 2241 6924 2284
rect 6806 2156 6924 2199
rect 6806 2124 6849 2156
rect 6849 2124 6881 2156
rect 6881 2124 6924 2156
rect 6806 2081 6924 2124
rect 6806 1996 6924 2039
rect 6806 1964 6849 1996
rect 6849 1964 6881 1996
rect 6881 1964 6924 1996
rect 6806 1921 6924 1964
rect 6806 1836 6924 1879
rect 6806 1804 6849 1836
rect 6849 1804 6881 1836
rect 6881 1804 6924 1836
rect 6806 1761 6924 1804
rect 6806 1676 6924 1719
rect 6806 1644 6849 1676
rect 6849 1644 6881 1676
rect 6881 1644 6924 1676
rect 6806 1601 6924 1644
rect 6806 1516 6924 1559
rect 6806 1484 6849 1516
rect 6849 1484 6881 1516
rect 6881 1484 6924 1516
rect 6806 1441 6924 1484
rect 6806 1356 6924 1399
rect 6806 1324 6849 1356
rect 6849 1324 6881 1356
rect 6881 1324 6924 1356
rect 6806 1281 6924 1324
rect 6806 1196 6924 1239
rect 6806 1164 6849 1196
rect 6849 1164 6881 1196
rect 6881 1164 6924 1196
rect 6806 1121 6924 1164
rect 6806 1036 6924 1079
rect 6806 1004 6849 1036
rect 6849 1004 6881 1036
rect 6881 1004 6924 1036
rect 6806 961 6924 1004
rect 6806 876 6924 919
rect 6806 844 6849 876
rect 6849 844 6881 876
rect 6881 844 6924 876
rect 6806 801 6924 844
rect 6806 716 6924 759
rect 6806 684 6849 716
rect 6849 684 6881 716
rect 6881 684 6924 716
rect 6806 641 6924 684
rect 6806 556 6924 599
rect 6806 524 6849 556
rect 6849 524 6881 556
rect 6881 524 6924 556
rect 6806 481 6924 524
rect 6806 396 6924 439
rect 6806 364 6849 396
rect 6849 364 6881 396
rect 6881 364 6924 396
rect 6806 321 6924 364
rect 6806 236 6924 279
rect 6806 204 6849 236
rect 6849 204 6881 236
rect 6881 204 6924 236
rect 6806 161 6924 204
rect 6806 76 6924 119
rect 6806 44 6849 76
rect 6849 44 6881 76
rect 6881 44 6924 76
rect 6806 1 6924 44
rect 6806 -84 6924 -41
rect 6806 -116 6849 -84
rect 6849 -116 6881 -84
rect 6881 -116 6924 -84
rect 6806 -159 6924 -116
rect 3073 -276 3116 -244
rect 3116 -276 3148 -244
rect 3148 -276 3191 -244
rect 3073 -319 3191 -276
rect 6806 -244 6924 -201
rect 6806 -276 6849 -244
rect 6849 -276 6881 -244
rect 6881 -276 6924 -244
rect 9261 3381 9379 3424
rect 9261 3349 9304 3381
rect 9304 3349 9336 3381
rect 9336 3349 9379 3381
rect 9073 3276 9191 3319
rect 9261 3306 9379 3349
rect 9421 3381 9539 3424
rect 9421 3349 9464 3381
rect 9464 3349 9496 3381
rect 9496 3349 9539 3381
rect 9421 3306 9539 3349
rect 9581 3381 9699 3424
rect 9581 3349 9624 3381
rect 9624 3349 9656 3381
rect 9656 3349 9699 3381
rect 9581 3306 9699 3349
rect 9741 3381 9859 3424
rect 9741 3349 9784 3381
rect 9784 3349 9816 3381
rect 9816 3349 9859 3381
rect 9741 3306 9859 3349
rect 9901 3381 10019 3424
rect 9901 3349 9944 3381
rect 9944 3349 9976 3381
rect 9976 3349 10019 3381
rect 9901 3306 10019 3349
rect 10061 3381 10179 3424
rect 10061 3349 10104 3381
rect 10104 3349 10136 3381
rect 10136 3349 10179 3381
rect 10061 3306 10179 3349
rect 10221 3381 10339 3424
rect 10221 3349 10264 3381
rect 10264 3349 10296 3381
rect 10296 3349 10339 3381
rect 10221 3306 10339 3349
rect 10381 3381 10499 3424
rect 10381 3349 10424 3381
rect 10424 3349 10456 3381
rect 10456 3349 10499 3381
rect 10381 3306 10499 3349
rect 10541 3381 10659 3424
rect 10541 3349 10584 3381
rect 10584 3349 10616 3381
rect 10616 3349 10659 3381
rect 10541 3306 10659 3349
rect 10701 3381 10819 3424
rect 10701 3349 10744 3381
rect 10744 3349 10776 3381
rect 10776 3349 10819 3381
rect 10701 3306 10819 3349
rect 10861 3381 10979 3424
rect 10861 3349 10904 3381
rect 10904 3349 10936 3381
rect 10936 3349 10979 3381
rect 10861 3306 10979 3349
rect 11021 3381 11139 3424
rect 11021 3349 11064 3381
rect 11064 3349 11096 3381
rect 11096 3349 11139 3381
rect 11021 3306 11139 3349
rect 11181 3381 11299 3424
rect 11181 3349 11224 3381
rect 11224 3349 11256 3381
rect 11256 3349 11299 3381
rect 11181 3306 11299 3349
rect 11341 3381 11459 3424
rect 11341 3349 11384 3381
rect 11384 3349 11416 3381
rect 11416 3349 11459 3381
rect 11341 3306 11459 3349
rect 11501 3381 11619 3424
rect 11501 3349 11544 3381
rect 11544 3349 11576 3381
rect 11576 3349 11619 3381
rect 11501 3306 11619 3349
rect 11661 3381 11779 3424
rect 11661 3349 11704 3381
rect 11704 3349 11736 3381
rect 11736 3349 11779 3381
rect 11661 3306 11779 3349
rect 11821 3381 11939 3424
rect 11821 3349 11864 3381
rect 11864 3349 11896 3381
rect 11896 3349 11939 3381
rect 11821 3306 11939 3349
rect 11981 3381 12099 3424
rect 11981 3349 12024 3381
rect 12024 3349 12056 3381
rect 12056 3349 12099 3381
rect 11981 3306 12099 3349
rect 12141 3381 12259 3424
rect 12141 3349 12184 3381
rect 12184 3349 12216 3381
rect 12216 3349 12259 3381
rect 12141 3306 12259 3349
rect 12301 3381 12419 3424
rect 12301 3349 12344 3381
rect 12344 3349 12376 3381
rect 12376 3349 12419 3381
rect 12301 3306 12419 3349
rect 12461 3381 12579 3424
rect 12461 3349 12504 3381
rect 12504 3349 12536 3381
rect 12536 3349 12579 3381
rect 12461 3306 12579 3349
rect 12621 3381 12739 3424
rect 12621 3349 12664 3381
rect 12664 3349 12696 3381
rect 12696 3349 12739 3381
rect 12621 3306 12739 3349
rect 9073 3244 9116 3276
rect 9116 3244 9148 3276
rect 9148 3244 9191 3276
rect 9073 3201 9191 3244
rect 12806 3276 12924 3319
rect 12806 3244 12849 3276
rect 12849 3244 12881 3276
rect 12881 3244 12924 3276
rect 9073 3116 9191 3159
rect 9073 3084 9116 3116
rect 9116 3084 9148 3116
rect 9148 3084 9191 3116
rect 9073 3041 9191 3084
rect 9073 2956 9191 2999
rect 9073 2924 9116 2956
rect 9116 2924 9148 2956
rect 9148 2924 9191 2956
rect 9073 2881 9191 2924
rect 9073 2796 9191 2839
rect 9073 2764 9116 2796
rect 9116 2764 9148 2796
rect 9148 2764 9191 2796
rect 9073 2721 9191 2764
rect 9073 2636 9191 2679
rect 9073 2604 9116 2636
rect 9116 2604 9148 2636
rect 9148 2604 9191 2636
rect 9073 2561 9191 2604
rect 9073 2476 9191 2519
rect 9073 2444 9116 2476
rect 9116 2444 9148 2476
rect 9148 2444 9191 2476
rect 9073 2401 9191 2444
rect 9073 2316 9191 2359
rect 9073 2284 9116 2316
rect 9116 2284 9148 2316
rect 9148 2284 9191 2316
rect 9073 2241 9191 2284
rect 9073 2156 9191 2199
rect 9073 2124 9116 2156
rect 9116 2124 9148 2156
rect 9148 2124 9191 2156
rect 9073 2081 9191 2124
rect 9073 1996 9191 2039
rect 9073 1964 9116 1996
rect 9116 1964 9148 1996
rect 9148 1964 9191 1996
rect 9073 1921 9191 1964
rect 9073 1836 9191 1879
rect 9073 1804 9116 1836
rect 9116 1804 9148 1836
rect 9148 1804 9191 1836
rect 9073 1761 9191 1804
rect 9073 1676 9191 1719
rect 9073 1644 9116 1676
rect 9116 1644 9148 1676
rect 9148 1644 9191 1676
rect 9073 1601 9191 1644
rect 9073 1516 9191 1559
rect 9073 1484 9116 1516
rect 9116 1484 9148 1516
rect 9148 1484 9191 1516
rect 9073 1441 9191 1484
rect 9073 1356 9191 1399
rect 9073 1324 9116 1356
rect 9116 1324 9148 1356
rect 9148 1324 9191 1356
rect 9073 1281 9191 1324
rect 9073 1196 9191 1239
rect 9073 1164 9116 1196
rect 9116 1164 9148 1196
rect 9148 1164 9191 1196
rect 9073 1121 9191 1164
rect 9073 1036 9191 1079
rect 9073 1004 9116 1036
rect 9116 1004 9148 1036
rect 9148 1004 9191 1036
rect 9073 961 9191 1004
rect 9073 876 9191 919
rect 9073 844 9116 876
rect 9116 844 9148 876
rect 9148 844 9191 876
rect 9073 801 9191 844
rect 9073 716 9191 759
rect 9073 684 9116 716
rect 9116 684 9148 716
rect 9148 684 9191 716
rect 9073 641 9191 684
rect 9073 556 9191 599
rect 9073 524 9116 556
rect 9116 524 9148 556
rect 9148 524 9191 556
rect 9073 481 9191 524
rect 9073 396 9191 439
rect 9073 364 9116 396
rect 9116 364 9148 396
rect 9148 364 9191 396
rect 9073 321 9191 364
rect 9073 236 9191 279
rect 9073 204 9116 236
rect 9116 204 9148 236
rect 9148 204 9191 236
rect 9073 161 9191 204
rect 9073 76 9191 119
rect 9073 44 9116 76
rect 9116 44 9148 76
rect 9148 44 9191 76
rect 9073 1 9191 44
rect 9073 -84 9191 -41
rect 9073 -116 9116 -84
rect 9116 -116 9148 -84
rect 9148 -116 9191 -84
rect 9073 -159 9191 -116
rect 3261 -347 3379 -304
rect 3261 -379 3304 -347
rect 3304 -379 3336 -347
rect 3336 -379 3379 -347
rect 3261 -422 3379 -379
rect 3421 -347 3539 -304
rect 3421 -379 3464 -347
rect 3464 -379 3496 -347
rect 3496 -379 3539 -347
rect 3421 -422 3539 -379
rect 3581 -347 3699 -304
rect 3581 -379 3624 -347
rect 3624 -379 3656 -347
rect 3656 -379 3699 -347
rect 3581 -422 3699 -379
rect 3741 -347 3859 -304
rect 3741 -379 3784 -347
rect 3784 -379 3816 -347
rect 3816 -379 3859 -347
rect 3741 -422 3859 -379
rect 3901 -347 4019 -304
rect 3901 -379 3944 -347
rect 3944 -379 3976 -347
rect 3976 -379 4019 -347
rect 3901 -422 4019 -379
rect 4061 -347 4179 -304
rect 4061 -379 4104 -347
rect 4104 -379 4136 -347
rect 4136 -379 4179 -347
rect 4061 -422 4179 -379
rect 4221 -347 4339 -304
rect 4221 -379 4264 -347
rect 4264 -379 4296 -347
rect 4296 -379 4339 -347
rect 4221 -422 4339 -379
rect 4381 -347 4499 -304
rect 4381 -379 4424 -347
rect 4424 -379 4456 -347
rect 4456 -379 4499 -347
rect 4381 -422 4499 -379
rect 4541 -347 4659 -304
rect 4541 -379 4584 -347
rect 4584 -379 4616 -347
rect 4616 -379 4659 -347
rect 4541 -422 4659 -379
rect 4701 -347 4819 -304
rect 4701 -379 4744 -347
rect 4744 -379 4776 -347
rect 4776 -379 4819 -347
rect 4701 -422 4819 -379
rect 4861 -347 4979 -304
rect 4861 -379 4904 -347
rect 4904 -379 4936 -347
rect 4936 -379 4979 -347
rect 4861 -422 4979 -379
rect 5021 -347 5139 -304
rect 5021 -379 5064 -347
rect 5064 -379 5096 -347
rect 5096 -379 5139 -347
rect 5021 -422 5139 -379
rect 5181 -347 5299 -304
rect 5181 -379 5224 -347
rect 5224 -379 5256 -347
rect 5256 -379 5299 -347
rect 5181 -422 5299 -379
rect 5341 -347 5459 -304
rect 5341 -379 5384 -347
rect 5384 -379 5416 -347
rect 5416 -379 5459 -347
rect 5341 -422 5459 -379
rect 5501 -347 5619 -304
rect 5501 -379 5544 -347
rect 5544 -379 5576 -347
rect 5576 -379 5619 -347
rect 5501 -422 5619 -379
rect 5661 -347 5779 -304
rect 5661 -379 5704 -347
rect 5704 -379 5736 -347
rect 5736 -379 5779 -347
rect 5661 -422 5779 -379
rect 5821 -347 5939 -304
rect 5821 -379 5864 -347
rect 5864 -379 5896 -347
rect 5896 -379 5939 -347
rect 5821 -422 5939 -379
rect 5981 -347 6099 -304
rect 5981 -379 6024 -347
rect 6024 -379 6056 -347
rect 6056 -379 6099 -347
rect 5981 -422 6099 -379
rect 6141 -347 6259 -304
rect 6141 -379 6184 -347
rect 6184 -379 6216 -347
rect 6216 -379 6259 -347
rect 6141 -422 6259 -379
rect 6301 -347 6419 -304
rect 6301 -379 6344 -347
rect 6344 -379 6376 -347
rect 6376 -379 6419 -347
rect 6301 -422 6419 -379
rect 6461 -347 6579 -304
rect 6461 -379 6504 -347
rect 6504 -379 6536 -347
rect 6536 -379 6579 -347
rect 6461 -422 6579 -379
rect 6621 -347 6739 -304
rect 6806 -319 6924 -276
rect 6621 -379 6664 -347
rect 6664 -379 6696 -347
rect 6696 -379 6739 -347
rect 6621 -422 6739 -379
rect 9073 -244 9191 -201
rect 12806 3201 12924 3244
rect 12806 3116 12924 3159
rect 12806 3084 12849 3116
rect 12849 3084 12881 3116
rect 12881 3084 12924 3116
rect 12806 3041 12924 3084
rect 12806 2956 12924 2999
rect 12806 2924 12849 2956
rect 12849 2924 12881 2956
rect 12881 2924 12924 2956
rect 12806 2881 12924 2924
rect 12806 2796 12924 2839
rect 12806 2764 12849 2796
rect 12849 2764 12881 2796
rect 12881 2764 12924 2796
rect 12806 2721 12924 2764
rect 12806 2636 12924 2679
rect 12806 2604 12849 2636
rect 12849 2604 12881 2636
rect 12881 2604 12924 2636
rect 12806 2561 12924 2604
rect 12806 2476 12924 2519
rect 12806 2444 12849 2476
rect 12849 2444 12881 2476
rect 12881 2444 12924 2476
rect 12806 2401 12924 2444
rect 12806 2316 12924 2359
rect 12806 2284 12849 2316
rect 12849 2284 12881 2316
rect 12881 2284 12924 2316
rect 12806 2241 12924 2284
rect 12806 2156 12924 2199
rect 12806 2124 12849 2156
rect 12849 2124 12881 2156
rect 12881 2124 12924 2156
rect 12806 2081 12924 2124
rect 12806 1996 12924 2039
rect 12806 1964 12849 1996
rect 12849 1964 12881 1996
rect 12881 1964 12924 1996
rect 12806 1921 12924 1964
rect 12806 1836 12924 1879
rect 12806 1804 12849 1836
rect 12849 1804 12881 1836
rect 12881 1804 12924 1836
rect 12806 1761 12924 1804
rect 12806 1676 12924 1719
rect 12806 1644 12849 1676
rect 12849 1644 12881 1676
rect 12881 1644 12924 1676
rect 12806 1601 12924 1644
rect 12806 1516 12924 1559
rect 12806 1484 12849 1516
rect 12849 1484 12881 1516
rect 12881 1484 12924 1516
rect 12806 1441 12924 1484
rect 12806 1356 12924 1399
rect 12806 1324 12849 1356
rect 12849 1324 12881 1356
rect 12881 1324 12924 1356
rect 12806 1281 12924 1324
rect 12806 1196 12924 1239
rect 12806 1164 12849 1196
rect 12849 1164 12881 1196
rect 12881 1164 12924 1196
rect 12806 1121 12924 1164
rect 12806 1036 12924 1079
rect 12806 1004 12849 1036
rect 12849 1004 12881 1036
rect 12881 1004 12924 1036
rect 12806 961 12924 1004
rect 12806 876 12924 919
rect 12806 844 12849 876
rect 12849 844 12881 876
rect 12881 844 12924 876
rect 12806 801 12924 844
rect 12806 716 12924 759
rect 12806 684 12849 716
rect 12849 684 12881 716
rect 12881 684 12924 716
rect 12806 641 12924 684
rect 12806 556 12924 599
rect 12806 524 12849 556
rect 12849 524 12881 556
rect 12881 524 12924 556
rect 12806 481 12924 524
rect 12806 396 12924 439
rect 12806 364 12849 396
rect 12849 364 12881 396
rect 12881 364 12924 396
rect 12806 321 12924 364
rect 12806 236 12924 279
rect 12806 204 12849 236
rect 12849 204 12881 236
rect 12881 204 12924 236
rect 12806 161 12924 204
rect 12806 76 12924 119
rect 12806 44 12849 76
rect 12849 44 12881 76
rect 12881 44 12924 76
rect 12806 1 12924 44
rect 12806 -84 12924 -41
rect 12806 -116 12849 -84
rect 12849 -116 12881 -84
rect 12881 -116 12924 -84
rect 12806 -159 12924 -116
rect 9073 -276 9116 -244
rect 9116 -276 9148 -244
rect 9148 -276 9191 -244
rect 9073 -319 9191 -276
rect 12806 -244 12924 -201
rect 12806 -276 12849 -244
rect 12849 -276 12881 -244
rect 12881 -276 12924 -244
rect 9261 -347 9379 -304
rect 9261 -379 9304 -347
rect 9304 -379 9336 -347
rect 9336 -379 9379 -347
rect 9261 -422 9379 -379
rect 9421 -347 9539 -304
rect 9421 -379 9464 -347
rect 9464 -379 9496 -347
rect 9496 -379 9539 -347
rect 9421 -422 9539 -379
rect 9581 -347 9699 -304
rect 9581 -379 9624 -347
rect 9624 -379 9656 -347
rect 9656 -379 9699 -347
rect 9581 -422 9699 -379
rect 9741 -347 9859 -304
rect 9741 -379 9784 -347
rect 9784 -379 9816 -347
rect 9816 -379 9859 -347
rect 9741 -422 9859 -379
rect 9901 -347 10019 -304
rect 9901 -379 9944 -347
rect 9944 -379 9976 -347
rect 9976 -379 10019 -347
rect 9901 -422 10019 -379
rect 10061 -347 10179 -304
rect 10061 -379 10104 -347
rect 10104 -379 10136 -347
rect 10136 -379 10179 -347
rect 10061 -422 10179 -379
rect 10221 -347 10339 -304
rect 10221 -379 10264 -347
rect 10264 -379 10296 -347
rect 10296 -379 10339 -347
rect 10221 -422 10339 -379
rect 10381 -347 10499 -304
rect 10381 -379 10424 -347
rect 10424 -379 10456 -347
rect 10456 -379 10499 -347
rect 10381 -422 10499 -379
rect 10541 -347 10659 -304
rect 10541 -379 10584 -347
rect 10584 -379 10616 -347
rect 10616 -379 10659 -347
rect 10541 -422 10659 -379
rect 10701 -347 10819 -304
rect 10701 -379 10744 -347
rect 10744 -379 10776 -347
rect 10776 -379 10819 -347
rect 10701 -422 10819 -379
rect 10861 -347 10979 -304
rect 10861 -379 10904 -347
rect 10904 -379 10936 -347
rect 10936 -379 10979 -347
rect 10861 -422 10979 -379
rect 11021 -347 11139 -304
rect 11021 -379 11064 -347
rect 11064 -379 11096 -347
rect 11096 -379 11139 -347
rect 11021 -422 11139 -379
rect 11181 -347 11299 -304
rect 11181 -379 11224 -347
rect 11224 -379 11256 -347
rect 11256 -379 11299 -347
rect 11181 -422 11299 -379
rect 11341 -347 11459 -304
rect 11341 -379 11384 -347
rect 11384 -379 11416 -347
rect 11416 -379 11459 -347
rect 11341 -422 11459 -379
rect 11501 -347 11619 -304
rect 11501 -379 11544 -347
rect 11544 -379 11576 -347
rect 11576 -379 11619 -347
rect 11501 -422 11619 -379
rect 11661 -347 11779 -304
rect 11661 -379 11704 -347
rect 11704 -379 11736 -347
rect 11736 -379 11779 -347
rect 11661 -422 11779 -379
rect 11821 -347 11939 -304
rect 11821 -379 11864 -347
rect 11864 -379 11896 -347
rect 11896 -379 11939 -347
rect 11821 -422 11939 -379
rect 11981 -347 12099 -304
rect 11981 -379 12024 -347
rect 12024 -379 12056 -347
rect 12056 -379 12099 -347
rect 11981 -422 12099 -379
rect 12141 -347 12259 -304
rect 12141 -379 12184 -347
rect 12184 -379 12216 -347
rect 12216 -379 12259 -347
rect 12141 -422 12259 -379
rect 12301 -347 12419 -304
rect 12301 -379 12344 -347
rect 12344 -379 12376 -347
rect 12376 -379 12419 -347
rect 12301 -422 12419 -379
rect 12461 -347 12579 -304
rect 12461 -379 12504 -347
rect 12504 -379 12536 -347
rect 12536 -379 12579 -347
rect 12461 -422 12579 -379
rect 12621 -347 12739 -304
rect 12806 -319 12924 -276
rect 12621 -379 12664 -347
rect 12664 -379 12696 -347
rect 12696 -379 12739 -347
rect 12621 -422 12739 -379
rect 15261 3381 15379 3424
rect 15261 3349 15304 3381
rect 15304 3349 15336 3381
rect 15336 3349 15379 3381
rect 15073 3276 15191 3319
rect 15261 3306 15379 3349
rect 15421 3381 15539 3424
rect 15421 3349 15464 3381
rect 15464 3349 15496 3381
rect 15496 3349 15539 3381
rect 15421 3306 15539 3349
rect 15581 3381 15699 3424
rect 15581 3349 15624 3381
rect 15624 3349 15656 3381
rect 15656 3349 15699 3381
rect 15581 3306 15699 3349
rect 15741 3381 15859 3424
rect 15741 3349 15784 3381
rect 15784 3349 15816 3381
rect 15816 3349 15859 3381
rect 15741 3306 15859 3349
rect 15901 3381 16019 3424
rect 15901 3349 15944 3381
rect 15944 3349 15976 3381
rect 15976 3349 16019 3381
rect 15901 3306 16019 3349
rect 16061 3381 16179 3424
rect 16061 3349 16104 3381
rect 16104 3349 16136 3381
rect 16136 3349 16179 3381
rect 16061 3306 16179 3349
rect 16221 3381 16339 3424
rect 16221 3349 16264 3381
rect 16264 3349 16296 3381
rect 16296 3349 16339 3381
rect 16221 3306 16339 3349
rect 16381 3381 16499 3424
rect 16381 3349 16424 3381
rect 16424 3349 16456 3381
rect 16456 3349 16499 3381
rect 16381 3306 16499 3349
rect 16541 3381 16659 3424
rect 16541 3349 16584 3381
rect 16584 3349 16616 3381
rect 16616 3349 16659 3381
rect 16541 3306 16659 3349
rect 16701 3381 16819 3424
rect 16701 3349 16744 3381
rect 16744 3349 16776 3381
rect 16776 3349 16819 3381
rect 16701 3306 16819 3349
rect 16861 3381 16979 3424
rect 16861 3349 16904 3381
rect 16904 3349 16936 3381
rect 16936 3349 16979 3381
rect 16861 3306 16979 3349
rect 17021 3381 17139 3424
rect 17021 3349 17064 3381
rect 17064 3349 17096 3381
rect 17096 3349 17139 3381
rect 17021 3306 17139 3349
rect 17181 3381 17299 3424
rect 17181 3349 17224 3381
rect 17224 3349 17256 3381
rect 17256 3349 17299 3381
rect 17181 3306 17299 3349
rect 17341 3381 17459 3424
rect 17341 3349 17384 3381
rect 17384 3349 17416 3381
rect 17416 3349 17459 3381
rect 17341 3306 17459 3349
rect 17501 3381 17619 3424
rect 17501 3349 17544 3381
rect 17544 3349 17576 3381
rect 17576 3349 17619 3381
rect 17501 3306 17619 3349
rect 17661 3381 17779 3424
rect 17661 3349 17704 3381
rect 17704 3349 17736 3381
rect 17736 3349 17779 3381
rect 17661 3306 17779 3349
rect 17821 3381 17939 3424
rect 17821 3349 17864 3381
rect 17864 3349 17896 3381
rect 17896 3349 17939 3381
rect 17821 3306 17939 3349
rect 17981 3381 18099 3424
rect 17981 3349 18024 3381
rect 18024 3349 18056 3381
rect 18056 3349 18099 3381
rect 17981 3306 18099 3349
rect 18141 3381 18259 3424
rect 18141 3349 18184 3381
rect 18184 3349 18216 3381
rect 18216 3349 18259 3381
rect 18141 3306 18259 3349
rect 18301 3381 18419 3424
rect 18301 3349 18344 3381
rect 18344 3349 18376 3381
rect 18376 3349 18419 3381
rect 18301 3306 18419 3349
rect 18461 3381 18579 3424
rect 18461 3349 18504 3381
rect 18504 3349 18536 3381
rect 18536 3349 18579 3381
rect 18461 3306 18579 3349
rect 18621 3381 18739 3424
rect 18621 3349 18664 3381
rect 18664 3349 18696 3381
rect 18696 3349 18739 3381
rect 18621 3306 18739 3349
rect 15073 3244 15116 3276
rect 15116 3244 15148 3276
rect 15148 3244 15191 3276
rect 15073 3201 15191 3244
rect 18806 3276 18924 3319
rect 18806 3244 18849 3276
rect 18849 3244 18881 3276
rect 18881 3244 18924 3276
rect 15073 3116 15191 3159
rect 15073 3084 15116 3116
rect 15116 3084 15148 3116
rect 15148 3084 15191 3116
rect 15073 3041 15191 3084
rect 15073 2956 15191 2999
rect 15073 2924 15116 2956
rect 15116 2924 15148 2956
rect 15148 2924 15191 2956
rect 15073 2881 15191 2924
rect 15073 2796 15191 2839
rect 15073 2764 15116 2796
rect 15116 2764 15148 2796
rect 15148 2764 15191 2796
rect 15073 2721 15191 2764
rect 15073 2636 15191 2679
rect 15073 2604 15116 2636
rect 15116 2604 15148 2636
rect 15148 2604 15191 2636
rect 15073 2561 15191 2604
rect 15073 2476 15191 2519
rect 15073 2444 15116 2476
rect 15116 2444 15148 2476
rect 15148 2444 15191 2476
rect 15073 2401 15191 2444
rect 15073 2316 15191 2359
rect 15073 2284 15116 2316
rect 15116 2284 15148 2316
rect 15148 2284 15191 2316
rect 15073 2241 15191 2284
rect 15073 2156 15191 2199
rect 15073 2124 15116 2156
rect 15116 2124 15148 2156
rect 15148 2124 15191 2156
rect 15073 2081 15191 2124
rect 15073 1996 15191 2039
rect 15073 1964 15116 1996
rect 15116 1964 15148 1996
rect 15148 1964 15191 1996
rect 15073 1921 15191 1964
rect 15073 1836 15191 1879
rect 15073 1804 15116 1836
rect 15116 1804 15148 1836
rect 15148 1804 15191 1836
rect 15073 1761 15191 1804
rect 15073 1676 15191 1719
rect 15073 1644 15116 1676
rect 15116 1644 15148 1676
rect 15148 1644 15191 1676
rect 15073 1601 15191 1644
rect 15073 1516 15191 1559
rect 15073 1484 15116 1516
rect 15116 1484 15148 1516
rect 15148 1484 15191 1516
rect 15073 1441 15191 1484
rect 15073 1356 15191 1399
rect 15073 1324 15116 1356
rect 15116 1324 15148 1356
rect 15148 1324 15191 1356
rect 15073 1281 15191 1324
rect 15073 1196 15191 1239
rect 15073 1164 15116 1196
rect 15116 1164 15148 1196
rect 15148 1164 15191 1196
rect 15073 1121 15191 1164
rect 15073 1036 15191 1079
rect 15073 1004 15116 1036
rect 15116 1004 15148 1036
rect 15148 1004 15191 1036
rect 15073 961 15191 1004
rect 15073 876 15191 919
rect 15073 844 15116 876
rect 15116 844 15148 876
rect 15148 844 15191 876
rect 15073 801 15191 844
rect 15073 716 15191 759
rect 15073 684 15116 716
rect 15116 684 15148 716
rect 15148 684 15191 716
rect 15073 641 15191 684
rect 15073 556 15191 599
rect 15073 524 15116 556
rect 15116 524 15148 556
rect 15148 524 15191 556
rect 15073 481 15191 524
rect 15073 396 15191 439
rect 15073 364 15116 396
rect 15116 364 15148 396
rect 15148 364 15191 396
rect 15073 321 15191 364
rect 15073 236 15191 279
rect 15073 204 15116 236
rect 15116 204 15148 236
rect 15148 204 15191 236
rect 15073 161 15191 204
rect 15073 76 15191 119
rect 15073 44 15116 76
rect 15116 44 15148 76
rect 15148 44 15191 76
rect 15073 1 15191 44
rect 15073 -84 15191 -41
rect 15073 -116 15116 -84
rect 15116 -116 15148 -84
rect 15148 -116 15191 -84
rect 15073 -159 15191 -116
rect 15073 -244 15191 -201
rect 18806 3201 18924 3244
rect 18806 3116 18924 3159
rect 18806 3084 18849 3116
rect 18849 3084 18881 3116
rect 18881 3084 18924 3116
rect 18806 3041 18924 3084
rect 18806 2956 18924 2999
rect 18806 2924 18849 2956
rect 18849 2924 18881 2956
rect 18881 2924 18924 2956
rect 18806 2881 18924 2924
rect 18806 2796 18924 2839
rect 18806 2764 18849 2796
rect 18849 2764 18881 2796
rect 18881 2764 18924 2796
rect 18806 2721 18924 2764
rect 18806 2636 18924 2679
rect 18806 2604 18849 2636
rect 18849 2604 18881 2636
rect 18881 2604 18924 2636
rect 18806 2561 18924 2604
rect 18806 2476 18924 2519
rect 18806 2444 18849 2476
rect 18849 2444 18881 2476
rect 18881 2444 18924 2476
rect 18806 2401 18924 2444
rect 18806 2316 18924 2359
rect 18806 2284 18849 2316
rect 18849 2284 18881 2316
rect 18881 2284 18924 2316
rect 18806 2241 18924 2284
rect 18806 2156 18924 2199
rect 18806 2124 18849 2156
rect 18849 2124 18881 2156
rect 18881 2124 18924 2156
rect 18806 2081 18924 2124
rect 18806 1996 18924 2039
rect 18806 1964 18849 1996
rect 18849 1964 18881 1996
rect 18881 1964 18924 1996
rect 18806 1921 18924 1964
rect 18806 1836 18924 1879
rect 18806 1804 18849 1836
rect 18849 1804 18881 1836
rect 18881 1804 18924 1836
rect 18806 1761 18924 1804
rect 18806 1676 18924 1719
rect 18806 1644 18849 1676
rect 18849 1644 18881 1676
rect 18881 1644 18924 1676
rect 18806 1601 18924 1644
rect 18806 1516 18924 1559
rect 18806 1484 18849 1516
rect 18849 1484 18881 1516
rect 18881 1484 18924 1516
rect 18806 1441 18924 1484
rect 18806 1356 18924 1399
rect 18806 1324 18849 1356
rect 18849 1324 18881 1356
rect 18881 1324 18924 1356
rect 18806 1281 18924 1324
rect 18806 1196 18924 1239
rect 18806 1164 18849 1196
rect 18849 1164 18881 1196
rect 18881 1164 18924 1196
rect 18806 1121 18924 1164
rect 18806 1036 18924 1079
rect 18806 1004 18849 1036
rect 18849 1004 18881 1036
rect 18881 1004 18924 1036
rect 18806 961 18924 1004
rect 18806 876 18924 919
rect 18806 844 18849 876
rect 18849 844 18881 876
rect 18881 844 18924 876
rect 18806 801 18924 844
rect 18806 716 18924 759
rect 18806 684 18849 716
rect 18849 684 18881 716
rect 18881 684 18924 716
rect 18806 641 18924 684
rect 18806 556 18924 599
rect 18806 524 18849 556
rect 18849 524 18881 556
rect 18881 524 18924 556
rect 18806 481 18924 524
rect 18806 396 18924 439
rect 18806 364 18849 396
rect 18849 364 18881 396
rect 18881 364 18924 396
rect 18806 321 18924 364
rect 18806 236 18924 279
rect 18806 204 18849 236
rect 18849 204 18881 236
rect 18881 204 18924 236
rect 18806 161 18924 204
rect 18806 76 18924 119
rect 18806 44 18849 76
rect 18849 44 18881 76
rect 18881 44 18924 76
rect 18806 1 18924 44
rect 18806 -84 18924 -41
rect 18806 -116 18849 -84
rect 18849 -116 18881 -84
rect 18881 -116 18924 -84
rect 18806 -159 18924 -116
rect 15073 -276 15116 -244
rect 15116 -276 15148 -244
rect 15148 -276 15191 -244
rect 15073 -319 15191 -276
rect 18806 -244 18924 -201
rect 18806 -276 18849 -244
rect 18849 -276 18881 -244
rect 18881 -276 18924 -244
rect 15261 -347 15379 -304
rect 15261 -379 15304 -347
rect 15304 -379 15336 -347
rect 15336 -379 15379 -347
rect 15261 -422 15379 -379
rect 15421 -347 15539 -304
rect 15421 -379 15464 -347
rect 15464 -379 15496 -347
rect 15496 -379 15539 -347
rect 15421 -422 15539 -379
rect 15581 -347 15699 -304
rect 15581 -379 15624 -347
rect 15624 -379 15656 -347
rect 15656 -379 15699 -347
rect 15581 -422 15699 -379
rect 15741 -347 15859 -304
rect 15741 -379 15784 -347
rect 15784 -379 15816 -347
rect 15816 -379 15859 -347
rect 15741 -422 15859 -379
rect 15901 -347 16019 -304
rect 15901 -379 15944 -347
rect 15944 -379 15976 -347
rect 15976 -379 16019 -347
rect 15901 -422 16019 -379
rect 16061 -347 16179 -304
rect 16061 -379 16104 -347
rect 16104 -379 16136 -347
rect 16136 -379 16179 -347
rect 16061 -422 16179 -379
rect 16221 -347 16339 -304
rect 16221 -379 16264 -347
rect 16264 -379 16296 -347
rect 16296 -379 16339 -347
rect 16221 -422 16339 -379
rect 16381 -347 16499 -304
rect 16381 -379 16424 -347
rect 16424 -379 16456 -347
rect 16456 -379 16499 -347
rect 16381 -422 16499 -379
rect 16541 -347 16659 -304
rect 16541 -379 16584 -347
rect 16584 -379 16616 -347
rect 16616 -379 16659 -347
rect 16541 -422 16659 -379
rect 16701 -347 16819 -304
rect 16701 -379 16744 -347
rect 16744 -379 16776 -347
rect 16776 -379 16819 -347
rect 16701 -422 16819 -379
rect 16861 -347 16979 -304
rect 16861 -379 16904 -347
rect 16904 -379 16936 -347
rect 16936 -379 16979 -347
rect 16861 -422 16979 -379
rect 17021 -347 17139 -304
rect 17021 -379 17064 -347
rect 17064 -379 17096 -347
rect 17096 -379 17139 -347
rect 17021 -422 17139 -379
rect 17181 -347 17299 -304
rect 17181 -379 17224 -347
rect 17224 -379 17256 -347
rect 17256 -379 17299 -347
rect 17181 -422 17299 -379
rect 17341 -347 17459 -304
rect 17341 -379 17384 -347
rect 17384 -379 17416 -347
rect 17416 -379 17459 -347
rect 17341 -422 17459 -379
rect 17501 -347 17619 -304
rect 17501 -379 17544 -347
rect 17544 -379 17576 -347
rect 17576 -379 17619 -347
rect 17501 -422 17619 -379
rect 17661 -347 17779 -304
rect 17661 -379 17704 -347
rect 17704 -379 17736 -347
rect 17736 -379 17779 -347
rect 17661 -422 17779 -379
rect 17821 -347 17939 -304
rect 17821 -379 17864 -347
rect 17864 -379 17896 -347
rect 17896 -379 17939 -347
rect 17821 -422 17939 -379
rect 17981 -347 18099 -304
rect 17981 -379 18024 -347
rect 18024 -379 18056 -347
rect 18056 -379 18099 -347
rect 17981 -422 18099 -379
rect 18141 -347 18259 -304
rect 18141 -379 18184 -347
rect 18184 -379 18216 -347
rect 18216 -379 18259 -347
rect 18141 -422 18259 -379
rect 18301 -347 18419 -304
rect 18301 -379 18344 -347
rect 18344 -379 18376 -347
rect 18376 -379 18419 -347
rect 18301 -422 18419 -379
rect 18461 -347 18579 -304
rect 18461 -379 18504 -347
rect 18504 -379 18536 -347
rect 18536 -379 18579 -347
rect 18461 -422 18579 -379
rect 18621 -347 18739 -304
rect 18806 -319 18924 -276
rect 18621 -379 18664 -347
rect 18664 -379 18696 -347
rect 18696 -379 18739 -347
rect 18621 -422 18739 -379
rect 21261 3381 21379 3424
rect 21261 3349 21304 3381
rect 21304 3349 21336 3381
rect 21336 3349 21379 3381
rect 21073 3276 21191 3319
rect 21261 3306 21379 3349
rect 21421 3381 21539 3424
rect 21421 3349 21464 3381
rect 21464 3349 21496 3381
rect 21496 3349 21539 3381
rect 21421 3306 21539 3349
rect 21581 3381 21699 3424
rect 21581 3349 21624 3381
rect 21624 3349 21656 3381
rect 21656 3349 21699 3381
rect 21581 3306 21699 3349
rect 21741 3381 21859 3424
rect 21741 3349 21784 3381
rect 21784 3349 21816 3381
rect 21816 3349 21859 3381
rect 21741 3306 21859 3349
rect 21901 3381 22019 3424
rect 21901 3349 21944 3381
rect 21944 3349 21976 3381
rect 21976 3349 22019 3381
rect 21901 3306 22019 3349
rect 22061 3381 22179 3424
rect 22061 3349 22104 3381
rect 22104 3349 22136 3381
rect 22136 3349 22179 3381
rect 22061 3306 22179 3349
rect 22221 3381 22339 3424
rect 22221 3349 22264 3381
rect 22264 3349 22296 3381
rect 22296 3349 22339 3381
rect 22221 3306 22339 3349
rect 22381 3381 22499 3424
rect 22381 3349 22424 3381
rect 22424 3349 22456 3381
rect 22456 3349 22499 3381
rect 22381 3306 22499 3349
rect 22541 3381 22659 3424
rect 22541 3349 22584 3381
rect 22584 3349 22616 3381
rect 22616 3349 22659 3381
rect 22541 3306 22659 3349
rect 22701 3381 22819 3424
rect 22701 3349 22744 3381
rect 22744 3349 22776 3381
rect 22776 3349 22819 3381
rect 22701 3306 22819 3349
rect 22861 3381 22979 3424
rect 22861 3349 22904 3381
rect 22904 3349 22936 3381
rect 22936 3349 22979 3381
rect 22861 3306 22979 3349
rect 23021 3381 23139 3424
rect 23021 3349 23064 3381
rect 23064 3349 23096 3381
rect 23096 3349 23139 3381
rect 23021 3306 23139 3349
rect 23181 3381 23299 3424
rect 23181 3349 23224 3381
rect 23224 3349 23256 3381
rect 23256 3349 23299 3381
rect 23181 3306 23299 3349
rect 23341 3381 23459 3424
rect 23341 3349 23384 3381
rect 23384 3349 23416 3381
rect 23416 3349 23459 3381
rect 23341 3306 23459 3349
rect 23501 3381 23619 3424
rect 23501 3349 23544 3381
rect 23544 3349 23576 3381
rect 23576 3349 23619 3381
rect 23501 3306 23619 3349
rect 23661 3381 23779 3424
rect 23661 3349 23704 3381
rect 23704 3349 23736 3381
rect 23736 3349 23779 3381
rect 23661 3306 23779 3349
rect 23821 3381 23939 3424
rect 23821 3349 23864 3381
rect 23864 3349 23896 3381
rect 23896 3349 23939 3381
rect 23821 3306 23939 3349
rect 23981 3381 24099 3424
rect 23981 3349 24024 3381
rect 24024 3349 24056 3381
rect 24056 3349 24099 3381
rect 23981 3306 24099 3349
rect 24141 3381 24259 3424
rect 24141 3349 24184 3381
rect 24184 3349 24216 3381
rect 24216 3349 24259 3381
rect 24141 3306 24259 3349
rect 24301 3381 24419 3424
rect 24301 3349 24344 3381
rect 24344 3349 24376 3381
rect 24376 3349 24419 3381
rect 24301 3306 24419 3349
rect 24461 3381 24579 3424
rect 24461 3349 24504 3381
rect 24504 3349 24536 3381
rect 24536 3349 24579 3381
rect 24461 3306 24579 3349
rect 24621 3381 24739 3424
rect 24621 3349 24664 3381
rect 24664 3349 24696 3381
rect 24696 3349 24739 3381
rect 24621 3306 24739 3349
rect 21073 3244 21116 3276
rect 21116 3244 21148 3276
rect 21148 3244 21191 3276
rect 21073 3201 21191 3244
rect 24806 3276 24924 3319
rect 24806 3244 24849 3276
rect 24849 3244 24881 3276
rect 24881 3244 24924 3276
rect 21073 3116 21191 3159
rect 21073 3084 21116 3116
rect 21116 3084 21148 3116
rect 21148 3084 21191 3116
rect 21073 3041 21191 3084
rect 21073 2956 21191 2999
rect 21073 2924 21116 2956
rect 21116 2924 21148 2956
rect 21148 2924 21191 2956
rect 21073 2881 21191 2924
rect 21073 2796 21191 2839
rect 21073 2764 21116 2796
rect 21116 2764 21148 2796
rect 21148 2764 21191 2796
rect 21073 2721 21191 2764
rect 21073 2636 21191 2679
rect 21073 2604 21116 2636
rect 21116 2604 21148 2636
rect 21148 2604 21191 2636
rect 21073 2561 21191 2604
rect 21073 2476 21191 2519
rect 21073 2444 21116 2476
rect 21116 2444 21148 2476
rect 21148 2444 21191 2476
rect 21073 2401 21191 2444
rect 21073 2316 21191 2359
rect 21073 2284 21116 2316
rect 21116 2284 21148 2316
rect 21148 2284 21191 2316
rect 21073 2241 21191 2284
rect 21073 2156 21191 2199
rect 21073 2124 21116 2156
rect 21116 2124 21148 2156
rect 21148 2124 21191 2156
rect 21073 2081 21191 2124
rect 21073 1996 21191 2039
rect 21073 1964 21116 1996
rect 21116 1964 21148 1996
rect 21148 1964 21191 1996
rect 21073 1921 21191 1964
rect 21073 1836 21191 1879
rect 21073 1804 21116 1836
rect 21116 1804 21148 1836
rect 21148 1804 21191 1836
rect 21073 1761 21191 1804
rect 21073 1676 21191 1719
rect 21073 1644 21116 1676
rect 21116 1644 21148 1676
rect 21148 1644 21191 1676
rect 21073 1601 21191 1644
rect 21073 1516 21191 1559
rect 21073 1484 21116 1516
rect 21116 1484 21148 1516
rect 21148 1484 21191 1516
rect 21073 1441 21191 1484
rect 21073 1356 21191 1399
rect 21073 1324 21116 1356
rect 21116 1324 21148 1356
rect 21148 1324 21191 1356
rect 21073 1281 21191 1324
rect 21073 1196 21191 1239
rect 21073 1164 21116 1196
rect 21116 1164 21148 1196
rect 21148 1164 21191 1196
rect 21073 1121 21191 1164
rect 21073 1036 21191 1079
rect 21073 1004 21116 1036
rect 21116 1004 21148 1036
rect 21148 1004 21191 1036
rect 21073 961 21191 1004
rect 21073 876 21191 919
rect 21073 844 21116 876
rect 21116 844 21148 876
rect 21148 844 21191 876
rect 21073 801 21191 844
rect 21073 716 21191 759
rect 21073 684 21116 716
rect 21116 684 21148 716
rect 21148 684 21191 716
rect 21073 641 21191 684
rect 21073 556 21191 599
rect 21073 524 21116 556
rect 21116 524 21148 556
rect 21148 524 21191 556
rect 21073 481 21191 524
rect 21073 396 21191 439
rect 21073 364 21116 396
rect 21116 364 21148 396
rect 21148 364 21191 396
rect 21073 321 21191 364
rect 21073 236 21191 279
rect 21073 204 21116 236
rect 21116 204 21148 236
rect 21148 204 21191 236
rect 21073 161 21191 204
rect 21073 76 21191 119
rect 21073 44 21116 76
rect 21116 44 21148 76
rect 21148 44 21191 76
rect 21073 1 21191 44
rect 21073 -84 21191 -41
rect 21073 -116 21116 -84
rect 21116 -116 21148 -84
rect 21148 -116 21191 -84
rect 21073 -159 21191 -116
rect 21073 -244 21191 -201
rect 24806 3201 24924 3244
rect 24806 3116 24924 3159
rect 24806 3084 24849 3116
rect 24849 3084 24881 3116
rect 24881 3084 24924 3116
rect 24806 3041 24924 3084
rect 24806 2956 24924 2999
rect 24806 2924 24849 2956
rect 24849 2924 24881 2956
rect 24881 2924 24924 2956
rect 24806 2881 24924 2924
rect 24806 2796 24924 2839
rect 24806 2764 24849 2796
rect 24849 2764 24881 2796
rect 24881 2764 24924 2796
rect 24806 2721 24924 2764
rect 24806 2636 24924 2679
rect 24806 2604 24849 2636
rect 24849 2604 24881 2636
rect 24881 2604 24924 2636
rect 24806 2561 24924 2604
rect 24806 2476 24924 2519
rect 24806 2444 24849 2476
rect 24849 2444 24881 2476
rect 24881 2444 24924 2476
rect 24806 2401 24924 2444
rect 24806 2316 24924 2359
rect 24806 2284 24849 2316
rect 24849 2284 24881 2316
rect 24881 2284 24924 2316
rect 24806 2241 24924 2284
rect 24806 2156 24924 2199
rect 24806 2124 24849 2156
rect 24849 2124 24881 2156
rect 24881 2124 24924 2156
rect 24806 2081 24924 2124
rect 24806 1996 24924 2039
rect 24806 1964 24849 1996
rect 24849 1964 24881 1996
rect 24881 1964 24924 1996
rect 24806 1921 24924 1964
rect 24806 1836 24924 1879
rect 24806 1804 24849 1836
rect 24849 1804 24881 1836
rect 24881 1804 24924 1836
rect 24806 1761 24924 1804
rect 24806 1676 24924 1719
rect 24806 1644 24849 1676
rect 24849 1644 24881 1676
rect 24881 1644 24924 1676
rect 24806 1601 24924 1644
rect 24806 1516 24924 1559
rect 24806 1484 24849 1516
rect 24849 1484 24881 1516
rect 24881 1484 24924 1516
rect 24806 1441 24924 1484
rect 24806 1356 24924 1399
rect 24806 1324 24849 1356
rect 24849 1324 24881 1356
rect 24881 1324 24924 1356
rect 24806 1281 24924 1324
rect 24806 1196 24924 1239
rect 24806 1164 24849 1196
rect 24849 1164 24881 1196
rect 24881 1164 24924 1196
rect 24806 1121 24924 1164
rect 24806 1036 24924 1079
rect 24806 1004 24849 1036
rect 24849 1004 24881 1036
rect 24881 1004 24924 1036
rect 24806 961 24924 1004
rect 24806 876 24924 919
rect 24806 844 24849 876
rect 24849 844 24881 876
rect 24881 844 24924 876
rect 24806 801 24924 844
rect 24806 716 24924 759
rect 24806 684 24849 716
rect 24849 684 24881 716
rect 24881 684 24924 716
rect 24806 641 24924 684
rect 24806 556 24924 599
rect 24806 524 24849 556
rect 24849 524 24881 556
rect 24881 524 24924 556
rect 24806 481 24924 524
rect 24806 396 24924 439
rect 24806 364 24849 396
rect 24849 364 24881 396
rect 24881 364 24924 396
rect 24806 321 24924 364
rect 24806 236 24924 279
rect 24806 204 24849 236
rect 24849 204 24881 236
rect 24881 204 24924 236
rect 24806 161 24924 204
rect 24806 76 24924 119
rect 24806 44 24849 76
rect 24849 44 24881 76
rect 24881 44 24924 76
rect 24806 1 24924 44
rect 24806 -84 24924 -41
rect 24806 -116 24849 -84
rect 24849 -116 24881 -84
rect 24881 -116 24924 -84
rect 24806 -159 24924 -116
rect 21073 -276 21116 -244
rect 21116 -276 21148 -244
rect 21148 -276 21191 -244
rect 21073 -319 21191 -276
rect 24806 -244 24924 -201
rect 24806 -276 24849 -244
rect 24849 -276 24881 -244
rect 24881 -276 24924 -244
rect 21261 -347 21379 -304
rect 21261 -379 21304 -347
rect 21304 -379 21336 -347
rect 21336 -379 21379 -347
rect 21261 -422 21379 -379
rect 21421 -347 21539 -304
rect 21421 -379 21464 -347
rect 21464 -379 21496 -347
rect 21496 -379 21539 -347
rect 21421 -422 21539 -379
rect 21581 -347 21699 -304
rect 21581 -379 21624 -347
rect 21624 -379 21656 -347
rect 21656 -379 21699 -347
rect 21581 -422 21699 -379
rect 21741 -347 21859 -304
rect 21741 -379 21784 -347
rect 21784 -379 21816 -347
rect 21816 -379 21859 -347
rect 21741 -422 21859 -379
rect 21901 -347 22019 -304
rect 21901 -379 21944 -347
rect 21944 -379 21976 -347
rect 21976 -379 22019 -347
rect 21901 -422 22019 -379
rect 22061 -347 22179 -304
rect 22061 -379 22104 -347
rect 22104 -379 22136 -347
rect 22136 -379 22179 -347
rect 22061 -422 22179 -379
rect 22221 -347 22339 -304
rect 22221 -379 22264 -347
rect 22264 -379 22296 -347
rect 22296 -379 22339 -347
rect 22221 -422 22339 -379
rect 22381 -347 22499 -304
rect 22381 -379 22424 -347
rect 22424 -379 22456 -347
rect 22456 -379 22499 -347
rect 22381 -422 22499 -379
rect 22541 -347 22659 -304
rect 22541 -379 22584 -347
rect 22584 -379 22616 -347
rect 22616 -379 22659 -347
rect 22541 -422 22659 -379
rect 22701 -347 22819 -304
rect 22701 -379 22744 -347
rect 22744 -379 22776 -347
rect 22776 -379 22819 -347
rect 22701 -422 22819 -379
rect 22861 -347 22979 -304
rect 22861 -379 22904 -347
rect 22904 -379 22936 -347
rect 22936 -379 22979 -347
rect 22861 -422 22979 -379
rect 23021 -347 23139 -304
rect 23021 -379 23064 -347
rect 23064 -379 23096 -347
rect 23096 -379 23139 -347
rect 23021 -422 23139 -379
rect 23181 -347 23299 -304
rect 23181 -379 23224 -347
rect 23224 -379 23256 -347
rect 23256 -379 23299 -347
rect 23181 -422 23299 -379
rect 23341 -347 23459 -304
rect 23341 -379 23384 -347
rect 23384 -379 23416 -347
rect 23416 -379 23459 -347
rect 23341 -422 23459 -379
rect 23501 -347 23619 -304
rect 23501 -379 23544 -347
rect 23544 -379 23576 -347
rect 23576 -379 23619 -347
rect 23501 -422 23619 -379
rect 23661 -347 23779 -304
rect 23661 -379 23704 -347
rect 23704 -379 23736 -347
rect 23736 -379 23779 -347
rect 23661 -422 23779 -379
rect 23821 -347 23939 -304
rect 23821 -379 23864 -347
rect 23864 -379 23896 -347
rect 23896 -379 23939 -347
rect 23821 -422 23939 -379
rect 23981 -347 24099 -304
rect 23981 -379 24024 -347
rect 24024 -379 24056 -347
rect 24056 -379 24099 -347
rect 23981 -422 24099 -379
rect 24141 -347 24259 -304
rect 24141 -379 24184 -347
rect 24184 -379 24216 -347
rect 24216 -379 24259 -347
rect 24141 -422 24259 -379
rect 24301 -347 24419 -304
rect 24301 -379 24344 -347
rect 24344 -379 24376 -347
rect 24376 -379 24419 -347
rect 24301 -422 24419 -379
rect 24461 -347 24579 -304
rect 24461 -379 24504 -347
rect 24504 -379 24536 -347
rect 24536 -379 24579 -347
rect 24461 -422 24579 -379
rect 24621 -347 24739 -304
rect 24806 -319 24924 -276
rect 24621 -379 24664 -347
rect 24664 -379 24696 -347
rect 24696 -379 24739 -347
rect 24621 -422 24739 -379
rect 3261 -5621 3379 -5578
rect 3261 -5653 3304 -5621
rect 3304 -5653 3336 -5621
rect 3336 -5653 3379 -5621
rect 3076 -5724 3194 -5681
rect 3261 -5696 3379 -5653
rect 3421 -5621 3539 -5578
rect 3421 -5653 3464 -5621
rect 3464 -5653 3496 -5621
rect 3496 -5653 3539 -5621
rect 3421 -5696 3539 -5653
rect 3581 -5621 3699 -5578
rect 3581 -5653 3624 -5621
rect 3624 -5653 3656 -5621
rect 3656 -5653 3699 -5621
rect 3581 -5696 3699 -5653
rect 3741 -5621 3859 -5578
rect 3741 -5653 3784 -5621
rect 3784 -5653 3816 -5621
rect 3816 -5653 3859 -5621
rect 3741 -5696 3859 -5653
rect 3901 -5621 4019 -5578
rect 3901 -5653 3944 -5621
rect 3944 -5653 3976 -5621
rect 3976 -5653 4019 -5621
rect 3901 -5696 4019 -5653
rect 4061 -5621 4179 -5578
rect 4061 -5653 4104 -5621
rect 4104 -5653 4136 -5621
rect 4136 -5653 4179 -5621
rect 4061 -5696 4179 -5653
rect 4221 -5621 4339 -5578
rect 4221 -5653 4264 -5621
rect 4264 -5653 4296 -5621
rect 4296 -5653 4339 -5621
rect 4221 -5696 4339 -5653
rect 4381 -5621 4499 -5578
rect 4381 -5653 4424 -5621
rect 4424 -5653 4456 -5621
rect 4456 -5653 4499 -5621
rect 4381 -5696 4499 -5653
rect 4541 -5621 4659 -5578
rect 4541 -5653 4584 -5621
rect 4584 -5653 4616 -5621
rect 4616 -5653 4659 -5621
rect 4541 -5696 4659 -5653
rect 4701 -5621 4819 -5578
rect 4701 -5653 4744 -5621
rect 4744 -5653 4776 -5621
rect 4776 -5653 4819 -5621
rect 4701 -5696 4819 -5653
rect 4861 -5621 4979 -5578
rect 4861 -5653 4904 -5621
rect 4904 -5653 4936 -5621
rect 4936 -5653 4979 -5621
rect 4861 -5696 4979 -5653
rect 5021 -5621 5139 -5578
rect 5021 -5653 5064 -5621
rect 5064 -5653 5096 -5621
rect 5096 -5653 5139 -5621
rect 5021 -5696 5139 -5653
rect 5181 -5621 5299 -5578
rect 5181 -5653 5224 -5621
rect 5224 -5653 5256 -5621
rect 5256 -5653 5299 -5621
rect 5181 -5696 5299 -5653
rect 5341 -5621 5459 -5578
rect 5341 -5653 5384 -5621
rect 5384 -5653 5416 -5621
rect 5416 -5653 5459 -5621
rect 5341 -5696 5459 -5653
rect 5501 -5621 5619 -5578
rect 5501 -5653 5544 -5621
rect 5544 -5653 5576 -5621
rect 5576 -5653 5619 -5621
rect 5501 -5696 5619 -5653
rect 5661 -5621 5779 -5578
rect 5661 -5653 5704 -5621
rect 5704 -5653 5736 -5621
rect 5736 -5653 5779 -5621
rect 5661 -5696 5779 -5653
rect 5821 -5621 5939 -5578
rect 5821 -5653 5864 -5621
rect 5864 -5653 5896 -5621
rect 5896 -5653 5939 -5621
rect 5821 -5696 5939 -5653
rect 5981 -5621 6099 -5578
rect 5981 -5653 6024 -5621
rect 6024 -5653 6056 -5621
rect 6056 -5653 6099 -5621
rect 5981 -5696 6099 -5653
rect 6141 -5621 6259 -5578
rect 6141 -5653 6184 -5621
rect 6184 -5653 6216 -5621
rect 6216 -5653 6259 -5621
rect 6141 -5696 6259 -5653
rect 6301 -5621 6419 -5578
rect 6301 -5653 6344 -5621
rect 6344 -5653 6376 -5621
rect 6376 -5653 6419 -5621
rect 6301 -5696 6419 -5653
rect 6461 -5621 6579 -5578
rect 6461 -5653 6504 -5621
rect 6504 -5653 6536 -5621
rect 6536 -5653 6579 -5621
rect 6461 -5696 6579 -5653
rect 6621 -5621 6739 -5578
rect 6621 -5653 6664 -5621
rect 6664 -5653 6696 -5621
rect 6696 -5653 6739 -5621
rect 6621 -5696 6739 -5653
rect 3076 -5756 3119 -5724
rect 3119 -5756 3151 -5724
rect 3151 -5756 3194 -5724
rect 3076 -5799 3194 -5756
rect 6809 -5724 6927 -5681
rect 6809 -5756 6852 -5724
rect 6852 -5756 6884 -5724
rect 6884 -5756 6927 -5724
rect 3076 -5884 3194 -5841
rect 3076 -5916 3119 -5884
rect 3119 -5916 3151 -5884
rect 3151 -5916 3194 -5884
rect 3076 -5959 3194 -5916
rect 3076 -6044 3194 -6001
rect 3076 -6076 3119 -6044
rect 3119 -6076 3151 -6044
rect 3151 -6076 3194 -6044
rect 3076 -6119 3194 -6076
rect 3076 -6204 3194 -6161
rect 3076 -6236 3119 -6204
rect 3119 -6236 3151 -6204
rect 3151 -6236 3194 -6204
rect 3076 -6279 3194 -6236
rect 3076 -6364 3194 -6321
rect 3076 -6396 3119 -6364
rect 3119 -6396 3151 -6364
rect 3151 -6396 3194 -6364
rect 3076 -6439 3194 -6396
rect 3076 -6524 3194 -6481
rect 3076 -6556 3119 -6524
rect 3119 -6556 3151 -6524
rect 3151 -6556 3194 -6524
rect 3076 -6599 3194 -6556
rect 3076 -6684 3194 -6641
rect 3076 -6716 3119 -6684
rect 3119 -6716 3151 -6684
rect 3151 -6716 3194 -6684
rect 3076 -6759 3194 -6716
rect 3076 -6844 3194 -6801
rect 3076 -6876 3119 -6844
rect 3119 -6876 3151 -6844
rect 3151 -6876 3194 -6844
rect 3076 -6919 3194 -6876
rect 3076 -7004 3194 -6961
rect 3076 -7036 3119 -7004
rect 3119 -7036 3151 -7004
rect 3151 -7036 3194 -7004
rect 3076 -7079 3194 -7036
rect 3076 -7164 3194 -7121
rect 3076 -7196 3119 -7164
rect 3119 -7196 3151 -7164
rect 3151 -7196 3194 -7164
rect 3076 -7239 3194 -7196
rect 3076 -7324 3194 -7281
rect 3076 -7356 3119 -7324
rect 3119 -7356 3151 -7324
rect 3151 -7356 3194 -7324
rect 3076 -7399 3194 -7356
rect 3076 -7484 3194 -7441
rect 3076 -7516 3119 -7484
rect 3119 -7516 3151 -7484
rect 3151 -7516 3194 -7484
rect 3076 -7559 3194 -7516
rect 3076 -7644 3194 -7601
rect 3076 -7676 3119 -7644
rect 3119 -7676 3151 -7644
rect 3151 -7676 3194 -7644
rect 3076 -7719 3194 -7676
rect 3076 -7804 3194 -7761
rect 3076 -7836 3119 -7804
rect 3119 -7836 3151 -7804
rect 3151 -7836 3194 -7804
rect 3076 -7879 3194 -7836
rect 3076 -7964 3194 -7921
rect 3076 -7996 3119 -7964
rect 3119 -7996 3151 -7964
rect 3151 -7996 3194 -7964
rect 3076 -8039 3194 -7996
rect 3076 -8124 3194 -8081
rect 3076 -8156 3119 -8124
rect 3119 -8156 3151 -8124
rect 3151 -8156 3194 -8124
rect 3076 -8199 3194 -8156
rect 3076 -8284 3194 -8241
rect 3076 -8316 3119 -8284
rect 3119 -8316 3151 -8284
rect 3151 -8316 3194 -8284
rect 3076 -8359 3194 -8316
rect 3076 -8444 3194 -8401
rect 3076 -8476 3119 -8444
rect 3119 -8476 3151 -8444
rect 3151 -8476 3194 -8444
rect 3076 -8519 3194 -8476
rect 3076 -8604 3194 -8561
rect 3076 -8636 3119 -8604
rect 3119 -8636 3151 -8604
rect 3151 -8636 3194 -8604
rect 3076 -8679 3194 -8636
rect 3076 -8764 3194 -8721
rect 3076 -8796 3119 -8764
rect 3119 -8796 3151 -8764
rect 3151 -8796 3194 -8764
rect 3076 -8839 3194 -8796
rect 3076 -8924 3194 -8881
rect 3076 -8956 3119 -8924
rect 3119 -8956 3151 -8924
rect 3151 -8956 3194 -8924
rect 3076 -8999 3194 -8956
rect 3076 -9084 3194 -9041
rect 3076 -9116 3119 -9084
rect 3119 -9116 3151 -9084
rect 3151 -9116 3194 -9084
rect 3076 -9159 3194 -9116
rect 3076 -9244 3194 -9201
rect 6809 -5799 6927 -5756
rect 6809 -5884 6927 -5841
rect 6809 -5916 6852 -5884
rect 6852 -5916 6884 -5884
rect 6884 -5916 6927 -5884
rect 6809 -5959 6927 -5916
rect 6809 -6044 6927 -6001
rect 6809 -6076 6852 -6044
rect 6852 -6076 6884 -6044
rect 6884 -6076 6927 -6044
rect 6809 -6119 6927 -6076
rect 6809 -6204 6927 -6161
rect 6809 -6236 6852 -6204
rect 6852 -6236 6884 -6204
rect 6884 -6236 6927 -6204
rect 6809 -6279 6927 -6236
rect 6809 -6364 6927 -6321
rect 6809 -6396 6852 -6364
rect 6852 -6396 6884 -6364
rect 6884 -6396 6927 -6364
rect 6809 -6439 6927 -6396
rect 6809 -6524 6927 -6481
rect 6809 -6556 6852 -6524
rect 6852 -6556 6884 -6524
rect 6884 -6556 6927 -6524
rect 6809 -6599 6927 -6556
rect 6809 -6684 6927 -6641
rect 6809 -6716 6852 -6684
rect 6852 -6716 6884 -6684
rect 6884 -6716 6927 -6684
rect 6809 -6759 6927 -6716
rect 6809 -6844 6927 -6801
rect 6809 -6876 6852 -6844
rect 6852 -6876 6884 -6844
rect 6884 -6876 6927 -6844
rect 6809 -6919 6927 -6876
rect 6809 -7004 6927 -6961
rect 6809 -7036 6852 -7004
rect 6852 -7036 6884 -7004
rect 6884 -7036 6927 -7004
rect 6809 -7079 6927 -7036
rect 6809 -7164 6927 -7121
rect 6809 -7196 6852 -7164
rect 6852 -7196 6884 -7164
rect 6884 -7196 6927 -7164
rect 6809 -7239 6927 -7196
rect 6809 -7324 6927 -7281
rect 6809 -7356 6852 -7324
rect 6852 -7356 6884 -7324
rect 6884 -7356 6927 -7324
rect 6809 -7399 6927 -7356
rect 6809 -7484 6927 -7441
rect 6809 -7516 6852 -7484
rect 6852 -7516 6884 -7484
rect 6884 -7516 6927 -7484
rect 6809 -7559 6927 -7516
rect 6809 -7644 6927 -7601
rect 6809 -7676 6852 -7644
rect 6852 -7676 6884 -7644
rect 6884 -7676 6927 -7644
rect 6809 -7719 6927 -7676
rect 6809 -7804 6927 -7761
rect 6809 -7836 6852 -7804
rect 6852 -7836 6884 -7804
rect 6884 -7836 6927 -7804
rect 6809 -7879 6927 -7836
rect 6809 -7964 6927 -7921
rect 6809 -7996 6852 -7964
rect 6852 -7996 6884 -7964
rect 6884 -7996 6927 -7964
rect 6809 -8039 6927 -7996
rect 6809 -8124 6927 -8081
rect 6809 -8156 6852 -8124
rect 6852 -8156 6884 -8124
rect 6884 -8156 6927 -8124
rect 6809 -8199 6927 -8156
rect 6809 -8284 6927 -8241
rect 6809 -8316 6852 -8284
rect 6852 -8316 6884 -8284
rect 6884 -8316 6927 -8284
rect 6809 -8359 6927 -8316
rect 6809 -8444 6927 -8401
rect 6809 -8476 6852 -8444
rect 6852 -8476 6884 -8444
rect 6884 -8476 6927 -8444
rect 6809 -8519 6927 -8476
rect 6809 -8604 6927 -8561
rect 6809 -8636 6852 -8604
rect 6852 -8636 6884 -8604
rect 6884 -8636 6927 -8604
rect 6809 -8679 6927 -8636
rect 6809 -8764 6927 -8721
rect 6809 -8796 6852 -8764
rect 6852 -8796 6884 -8764
rect 6884 -8796 6927 -8764
rect 6809 -8839 6927 -8796
rect 6809 -8924 6927 -8881
rect 6809 -8956 6852 -8924
rect 6852 -8956 6884 -8924
rect 6884 -8956 6927 -8924
rect 6809 -8999 6927 -8956
rect 6809 -9084 6927 -9041
rect 6809 -9116 6852 -9084
rect 6852 -9116 6884 -9084
rect 6884 -9116 6927 -9084
rect 6809 -9159 6927 -9116
rect 3076 -9276 3119 -9244
rect 3119 -9276 3151 -9244
rect 3151 -9276 3194 -9244
rect 3076 -9319 3194 -9276
rect 6809 -9244 6927 -9201
rect 6809 -9276 6852 -9244
rect 6852 -9276 6884 -9244
rect 6884 -9276 6927 -9244
rect 3261 -9349 3379 -9306
rect 3261 -9381 3304 -9349
rect 3304 -9381 3336 -9349
rect 3336 -9381 3379 -9349
rect 3261 -9424 3379 -9381
rect 3421 -9349 3539 -9306
rect 3421 -9381 3464 -9349
rect 3464 -9381 3496 -9349
rect 3496 -9381 3539 -9349
rect 3421 -9424 3539 -9381
rect 3581 -9349 3699 -9306
rect 3581 -9381 3624 -9349
rect 3624 -9381 3656 -9349
rect 3656 -9381 3699 -9349
rect 3581 -9424 3699 -9381
rect 3741 -9349 3859 -9306
rect 3741 -9381 3784 -9349
rect 3784 -9381 3816 -9349
rect 3816 -9381 3859 -9349
rect 3741 -9424 3859 -9381
rect 3901 -9349 4019 -9306
rect 3901 -9381 3944 -9349
rect 3944 -9381 3976 -9349
rect 3976 -9381 4019 -9349
rect 3901 -9424 4019 -9381
rect 4061 -9349 4179 -9306
rect 4061 -9381 4104 -9349
rect 4104 -9381 4136 -9349
rect 4136 -9381 4179 -9349
rect 4061 -9424 4179 -9381
rect 4221 -9349 4339 -9306
rect 4221 -9381 4264 -9349
rect 4264 -9381 4296 -9349
rect 4296 -9381 4339 -9349
rect 4221 -9424 4339 -9381
rect 4381 -9349 4499 -9306
rect 4381 -9381 4424 -9349
rect 4424 -9381 4456 -9349
rect 4456 -9381 4499 -9349
rect 4381 -9424 4499 -9381
rect 4541 -9349 4659 -9306
rect 4541 -9381 4584 -9349
rect 4584 -9381 4616 -9349
rect 4616 -9381 4659 -9349
rect 4541 -9424 4659 -9381
rect 4701 -9349 4819 -9306
rect 4701 -9381 4744 -9349
rect 4744 -9381 4776 -9349
rect 4776 -9381 4819 -9349
rect 4701 -9424 4819 -9381
rect 4861 -9349 4979 -9306
rect 4861 -9381 4904 -9349
rect 4904 -9381 4936 -9349
rect 4936 -9381 4979 -9349
rect 4861 -9424 4979 -9381
rect 5021 -9349 5139 -9306
rect 5021 -9381 5064 -9349
rect 5064 -9381 5096 -9349
rect 5096 -9381 5139 -9349
rect 5021 -9424 5139 -9381
rect 5181 -9349 5299 -9306
rect 5181 -9381 5224 -9349
rect 5224 -9381 5256 -9349
rect 5256 -9381 5299 -9349
rect 5181 -9424 5299 -9381
rect 5341 -9349 5459 -9306
rect 5341 -9381 5384 -9349
rect 5384 -9381 5416 -9349
rect 5416 -9381 5459 -9349
rect 5341 -9424 5459 -9381
rect 5501 -9349 5619 -9306
rect 5501 -9381 5544 -9349
rect 5544 -9381 5576 -9349
rect 5576 -9381 5619 -9349
rect 5501 -9424 5619 -9381
rect 5661 -9349 5779 -9306
rect 5661 -9381 5704 -9349
rect 5704 -9381 5736 -9349
rect 5736 -9381 5779 -9349
rect 5661 -9424 5779 -9381
rect 5821 -9349 5939 -9306
rect 5821 -9381 5864 -9349
rect 5864 -9381 5896 -9349
rect 5896 -9381 5939 -9349
rect 5821 -9424 5939 -9381
rect 5981 -9349 6099 -9306
rect 5981 -9381 6024 -9349
rect 6024 -9381 6056 -9349
rect 6056 -9381 6099 -9349
rect 5981 -9424 6099 -9381
rect 6141 -9349 6259 -9306
rect 6141 -9381 6184 -9349
rect 6184 -9381 6216 -9349
rect 6216 -9381 6259 -9349
rect 6141 -9424 6259 -9381
rect 6301 -9349 6419 -9306
rect 6301 -9381 6344 -9349
rect 6344 -9381 6376 -9349
rect 6376 -9381 6419 -9349
rect 6301 -9424 6419 -9381
rect 6461 -9349 6579 -9306
rect 6461 -9381 6504 -9349
rect 6504 -9381 6536 -9349
rect 6536 -9381 6579 -9349
rect 6461 -9424 6579 -9381
rect 6621 -9349 6739 -9306
rect 6809 -9319 6927 -9276
rect 6621 -9381 6664 -9349
rect 6664 -9381 6696 -9349
rect 6696 -9381 6739 -9349
rect 6621 -9424 6739 -9381
rect 9261 -5621 9379 -5578
rect 9261 -5653 9304 -5621
rect 9304 -5653 9336 -5621
rect 9336 -5653 9379 -5621
rect 9076 -5724 9194 -5681
rect 9261 -5696 9379 -5653
rect 9421 -5621 9539 -5578
rect 9421 -5653 9464 -5621
rect 9464 -5653 9496 -5621
rect 9496 -5653 9539 -5621
rect 9421 -5696 9539 -5653
rect 9581 -5621 9699 -5578
rect 9581 -5653 9624 -5621
rect 9624 -5653 9656 -5621
rect 9656 -5653 9699 -5621
rect 9581 -5696 9699 -5653
rect 9741 -5621 9859 -5578
rect 9741 -5653 9784 -5621
rect 9784 -5653 9816 -5621
rect 9816 -5653 9859 -5621
rect 9741 -5696 9859 -5653
rect 9901 -5621 10019 -5578
rect 9901 -5653 9944 -5621
rect 9944 -5653 9976 -5621
rect 9976 -5653 10019 -5621
rect 9901 -5696 10019 -5653
rect 10061 -5621 10179 -5578
rect 10061 -5653 10104 -5621
rect 10104 -5653 10136 -5621
rect 10136 -5653 10179 -5621
rect 10061 -5696 10179 -5653
rect 10221 -5621 10339 -5578
rect 10221 -5653 10264 -5621
rect 10264 -5653 10296 -5621
rect 10296 -5653 10339 -5621
rect 10221 -5696 10339 -5653
rect 10381 -5621 10499 -5578
rect 10381 -5653 10424 -5621
rect 10424 -5653 10456 -5621
rect 10456 -5653 10499 -5621
rect 10381 -5696 10499 -5653
rect 10541 -5621 10659 -5578
rect 10541 -5653 10584 -5621
rect 10584 -5653 10616 -5621
rect 10616 -5653 10659 -5621
rect 10541 -5696 10659 -5653
rect 10701 -5621 10819 -5578
rect 10701 -5653 10744 -5621
rect 10744 -5653 10776 -5621
rect 10776 -5653 10819 -5621
rect 10701 -5696 10819 -5653
rect 10861 -5621 10979 -5578
rect 10861 -5653 10904 -5621
rect 10904 -5653 10936 -5621
rect 10936 -5653 10979 -5621
rect 10861 -5696 10979 -5653
rect 11021 -5621 11139 -5578
rect 11021 -5653 11064 -5621
rect 11064 -5653 11096 -5621
rect 11096 -5653 11139 -5621
rect 11021 -5696 11139 -5653
rect 11181 -5621 11299 -5578
rect 11181 -5653 11224 -5621
rect 11224 -5653 11256 -5621
rect 11256 -5653 11299 -5621
rect 11181 -5696 11299 -5653
rect 11341 -5621 11459 -5578
rect 11341 -5653 11384 -5621
rect 11384 -5653 11416 -5621
rect 11416 -5653 11459 -5621
rect 11341 -5696 11459 -5653
rect 11501 -5621 11619 -5578
rect 11501 -5653 11544 -5621
rect 11544 -5653 11576 -5621
rect 11576 -5653 11619 -5621
rect 11501 -5696 11619 -5653
rect 11661 -5621 11779 -5578
rect 11661 -5653 11704 -5621
rect 11704 -5653 11736 -5621
rect 11736 -5653 11779 -5621
rect 11661 -5696 11779 -5653
rect 11821 -5621 11939 -5578
rect 11821 -5653 11864 -5621
rect 11864 -5653 11896 -5621
rect 11896 -5653 11939 -5621
rect 11821 -5696 11939 -5653
rect 11981 -5621 12099 -5578
rect 11981 -5653 12024 -5621
rect 12024 -5653 12056 -5621
rect 12056 -5653 12099 -5621
rect 11981 -5696 12099 -5653
rect 12141 -5621 12259 -5578
rect 12141 -5653 12184 -5621
rect 12184 -5653 12216 -5621
rect 12216 -5653 12259 -5621
rect 12141 -5696 12259 -5653
rect 12301 -5621 12419 -5578
rect 12301 -5653 12344 -5621
rect 12344 -5653 12376 -5621
rect 12376 -5653 12419 -5621
rect 12301 -5696 12419 -5653
rect 12461 -5621 12579 -5578
rect 12461 -5653 12504 -5621
rect 12504 -5653 12536 -5621
rect 12536 -5653 12579 -5621
rect 12461 -5696 12579 -5653
rect 12621 -5621 12739 -5578
rect 12621 -5653 12664 -5621
rect 12664 -5653 12696 -5621
rect 12696 -5653 12739 -5621
rect 12621 -5696 12739 -5653
rect 9076 -5756 9119 -5724
rect 9119 -5756 9151 -5724
rect 9151 -5756 9194 -5724
rect 9076 -5799 9194 -5756
rect 12809 -5724 12927 -5681
rect 12809 -5756 12852 -5724
rect 12852 -5756 12884 -5724
rect 12884 -5756 12927 -5724
rect 9076 -5884 9194 -5841
rect 9076 -5916 9119 -5884
rect 9119 -5916 9151 -5884
rect 9151 -5916 9194 -5884
rect 9076 -5959 9194 -5916
rect 9076 -6044 9194 -6001
rect 9076 -6076 9119 -6044
rect 9119 -6076 9151 -6044
rect 9151 -6076 9194 -6044
rect 9076 -6119 9194 -6076
rect 9076 -6204 9194 -6161
rect 9076 -6236 9119 -6204
rect 9119 -6236 9151 -6204
rect 9151 -6236 9194 -6204
rect 9076 -6279 9194 -6236
rect 9076 -6364 9194 -6321
rect 9076 -6396 9119 -6364
rect 9119 -6396 9151 -6364
rect 9151 -6396 9194 -6364
rect 9076 -6439 9194 -6396
rect 9076 -6524 9194 -6481
rect 9076 -6556 9119 -6524
rect 9119 -6556 9151 -6524
rect 9151 -6556 9194 -6524
rect 9076 -6599 9194 -6556
rect 9076 -6684 9194 -6641
rect 9076 -6716 9119 -6684
rect 9119 -6716 9151 -6684
rect 9151 -6716 9194 -6684
rect 9076 -6759 9194 -6716
rect 9076 -6844 9194 -6801
rect 9076 -6876 9119 -6844
rect 9119 -6876 9151 -6844
rect 9151 -6876 9194 -6844
rect 9076 -6919 9194 -6876
rect 9076 -7004 9194 -6961
rect 9076 -7036 9119 -7004
rect 9119 -7036 9151 -7004
rect 9151 -7036 9194 -7004
rect 9076 -7079 9194 -7036
rect 9076 -7164 9194 -7121
rect 9076 -7196 9119 -7164
rect 9119 -7196 9151 -7164
rect 9151 -7196 9194 -7164
rect 9076 -7239 9194 -7196
rect 9076 -7324 9194 -7281
rect 9076 -7356 9119 -7324
rect 9119 -7356 9151 -7324
rect 9151 -7356 9194 -7324
rect 9076 -7399 9194 -7356
rect 9076 -7484 9194 -7441
rect 9076 -7516 9119 -7484
rect 9119 -7516 9151 -7484
rect 9151 -7516 9194 -7484
rect 9076 -7559 9194 -7516
rect 9076 -7644 9194 -7601
rect 9076 -7676 9119 -7644
rect 9119 -7676 9151 -7644
rect 9151 -7676 9194 -7644
rect 9076 -7719 9194 -7676
rect 9076 -7804 9194 -7761
rect 9076 -7836 9119 -7804
rect 9119 -7836 9151 -7804
rect 9151 -7836 9194 -7804
rect 9076 -7879 9194 -7836
rect 9076 -7964 9194 -7921
rect 9076 -7996 9119 -7964
rect 9119 -7996 9151 -7964
rect 9151 -7996 9194 -7964
rect 9076 -8039 9194 -7996
rect 9076 -8124 9194 -8081
rect 9076 -8156 9119 -8124
rect 9119 -8156 9151 -8124
rect 9151 -8156 9194 -8124
rect 9076 -8199 9194 -8156
rect 9076 -8284 9194 -8241
rect 9076 -8316 9119 -8284
rect 9119 -8316 9151 -8284
rect 9151 -8316 9194 -8284
rect 9076 -8359 9194 -8316
rect 9076 -8444 9194 -8401
rect 9076 -8476 9119 -8444
rect 9119 -8476 9151 -8444
rect 9151 -8476 9194 -8444
rect 9076 -8519 9194 -8476
rect 9076 -8604 9194 -8561
rect 9076 -8636 9119 -8604
rect 9119 -8636 9151 -8604
rect 9151 -8636 9194 -8604
rect 9076 -8679 9194 -8636
rect 9076 -8764 9194 -8721
rect 9076 -8796 9119 -8764
rect 9119 -8796 9151 -8764
rect 9151 -8796 9194 -8764
rect 9076 -8839 9194 -8796
rect 9076 -8924 9194 -8881
rect 9076 -8956 9119 -8924
rect 9119 -8956 9151 -8924
rect 9151 -8956 9194 -8924
rect 9076 -8999 9194 -8956
rect 9076 -9084 9194 -9041
rect 9076 -9116 9119 -9084
rect 9119 -9116 9151 -9084
rect 9151 -9116 9194 -9084
rect 9076 -9159 9194 -9116
rect 9076 -9244 9194 -9201
rect 12809 -5799 12927 -5756
rect 12809 -5884 12927 -5841
rect 12809 -5916 12852 -5884
rect 12852 -5916 12884 -5884
rect 12884 -5916 12927 -5884
rect 12809 -5959 12927 -5916
rect 12809 -6044 12927 -6001
rect 12809 -6076 12852 -6044
rect 12852 -6076 12884 -6044
rect 12884 -6076 12927 -6044
rect 12809 -6119 12927 -6076
rect 12809 -6204 12927 -6161
rect 12809 -6236 12852 -6204
rect 12852 -6236 12884 -6204
rect 12884 -6236 12927 -6204
rect 12809 -6279 12927 -6236
rect 12809 -6364 12927 -6321
rect 12809 -6396 12852 -6364
rect 12852 -6396 12884 -6364
rect 12884 -6396 12927 -6364
rect 12809 -6439 12927 -6396
rect 12809 -6524 12927 -6481
rect 12809 -6556 12852 -6524
rect 12852 -6556 12884 -6524
rect 12884 -6556 12927 -6524
rect 12809 -6599 12927 -6556
rect 12809 -6684 12927 -6641
rect 12809 -6716 12852 -6684
rect 12852 -6716 12884 -6684
rect 12884 -6716 12927 -6684
rect 12809 -6759 12927 -6716
rect 12809 -6844 12927 -6801
rect 12809 -6876 12852 -6844
rect 12852 -6876 12884 -6844
rect 12884 -6876 12927 -6844
rect 12809 -6919 12927 -6876
rect 12809 -7004 12927 -6961
rect 12809 -7036 12852 -7004
rect 12852 -7036 12884 -7004
rect 12884 -7036 12927 -7004
rect 12809 -7079 12927 -7036
rect 12809 -7164 12927 -7121
rect 12809 -7196 12852 -7164
rect 12852 -7196 12884 -7164
rect 12884 -7196 12927 -7164
rect 12809 -7239 12927 -7196
rect 12809 -7324 12927 -7281
rect 12809 -7356 12852 -7324
rect 12852 -7356 12884 -7324
rect 12884 -7356 12927 -7324
rect 12809 -7399 12927 -7356
rect 12809 -7484 12927 -7441
rect 12809 -7516 12852 -7484
rect 12852 -7516 12884 -7484
rect 12884 -7516 12927 -7484
rect 12809 -7559 12927 -7516
rect 12809 -7644 12927 -7601
rect 12809 -7676 12852 -7644
rect 12852 -7676 12884 -7644
rect 12884 -7676 12927 -7644
rect 12809 -7719 12927 -7676
rect 12809 -7804 12927 -7761
rect 12809 -7836 12852 -7804
rect 12852 -7836 12884 -7804
rect 12884 -7836 12927 -7804
rect 12809 -7879 12927 -7836
rect 12809 -7964 12927 -7921
rect 12809 -7996 12852 -7964
rect 12852 -7996 12884 -7964
rect 12884 -7996 12927 -7964
rect 12809 -8039 12927 -7996
rect 12809 -8124 12927 -8081
rect 12809 -8156 12852 -8124
rect 12852 -8156 12884 -8124
rect 12884 -8156 12927 -8124
rect 12809 -8199 12927 -8156
rect 12809 -8284 12927 -8241
rect 12809 -8316 12852 -8284
rect 12852 -8316 12884 -8284
rect 12884 -8316 12927 -8284
rect 12809 -8359 12927 -8316
rect 12809 -8444 12927 -8401
rect 12809 -8476 12852 -8444
rect 12852 -8476 12884 -8444
rect 12884 -8476 12927 -8444
rect 12809 -8519 12927 -8476
rect 12809 -8604 12927 -8561
rect 12809 -8636 12852 -8604
rect 12852 -8636 12884 -8604
rect 12884 -8636 12927 -8604
rect 12809 -8679 12927 -8636
rect 12809 -8764 12927 -8721
rect 12809 -8796 12852 -8764
rect 12852 -8796 12884 -8764
rect 12884 -8796 12927 -8764
rect 12809 -8839 12927 -8796
rect 12809 -8924 12927 -8881
rect 12809 -8956 12852 -8924
rect 12852 -8956 12884 -8924
rect 12884 -8956 12927 -8924
rect 12809 -8999 12927 -8956
rect 12809 -9084 12927 -9041
rect 12809 -9116 12852 -9084
rect 12852 -9116 12884 -9084
rect 12884 -9116 12927 -9084
rect 12809 -9159 12927 -9116
rect 9076 -9276 9119 -9244
rect 9119 -9276 9151 -9244
rect 9151 -9276 9194 -9244
rect 9076 -9319 9194 -9276
rect 12809 -9244 12927 -9201
rect 12809 -9276 12852 -9244
rect 12852 -9276 12884 -9244
rect 12884 -9276 12927 -9244
rect 9261 -9349 9379 -9306
rect 9261 -9381 9304 -9349
rect 9304 -9381 9336 -9349
rect 9336 -9381 9379 -9349
rect 9261 -9424 9379 -9381
rect 9421 -9349 9539 -9306
rect 9421 -9381 9464 -9349
rect 9464 -9381 9496 -9349
rect 9496 -9381 9539 -9349
rect 9421 -9424 9539 -9381
rect 9581 -9349 9699 -9306
rect 9581 -9381 9624 -9349
rect 9624 -9381 9656 -9349
rect 9656 -9381 9699 -9349
rect 9581 -9424 9699 -9381
rect 9741 -9349 9859 -9306
rect 9741 -9381 9784 -9349
rect 9784 -9381 9816 -9349
rect 9816 -9381 9859 -9349
rect 9741 -9424 9859 -9381
rect 9901 -9349 10019 -9306
rect 9901 -9381 9944 -9349
rect 9944 -9381 9976 -9349
rect 9976 -9381 10019 -9349
rect 9901 -9424 10019 -9381
rect 10061 -9349 10179 -9306
rect 10061 -9381 10104 -9349
rect 10104 -9381 10136 -9349
rect 10136 -9381 10179 -9349
rect 10061 -9424 10179 -9381
rect 10221 -9349 10339 -9306
rect 10221 -9381 10264 -9349
rect 10264 -9381 10296 -9349
rect 10296 -9381 10339 -9349
rect 10221 -9424 10339 -9381
rect 10381 -9349 10499 -9306
rect 10381 -9381 10424 -9349
rect 10424 -9381 10456 -9349
rect 10456 -9381 10499 -9349
rect 10381 -9424 10499 -9381
rect 10541 -9349 10659 -9306
rect 10541 -9381 10584 -9349
rect 10584 -9381 10616 -9349
rect 10616 -9381 10659 -9349
rect 10541 -9424 10659 -9381
rect 10701 -9349 10819 -9306
rect 10701 -9381 10744 -9349
rect 10744 -9381 10776 -9349
rect 10776 -9381 10819 -9349
rect 10701 -9424 10819 -9381
rect 10861 -9349 10979 -9306
rect 10861 -9381 10904 -9349
rect 10904 -9381 10936 -9349
rect 10936 -9381 10979 -9349
rect 10861 -9424 10979 -9381
rect 11021 -9349 11139 -9306
rect 11021 -9381 11064 -9349
rect 11064 -9381 11096 -9349
rect 11096 -9381 11139 -9349
rect 11021 -9424 11139 -9381
rect 11181 -9349 11299 -9306
rect 11181 -9381 11224 -9349
rect 11224 -9381 11256 -9349
rect 11256 -9381 11299 -9349
rect 11181 -9424 11299 -9381
rect 11341 -9349 11459 -9306
rect 11341 -9381 11384 -9349
rect 11384 -9381 11416 -9349
rect 11416 -9381 11459 -9349
rect 11341 -9424 11459 -9381
rect 11501 -9349 11619 -9306
rect 11501 -9381 11544 -9349
rect 11544 -9381 11576 -9349
rect 11576 -9381 11619 -9349
rect 11501 -9424 11619 -9381
rect 11661 -9349 11779 -9306
rect 11661 -9381 11704 -9349
rect 11704 -9381 11736 -9349
rect 11736 -9381 11779 -9349
rect 11661 -9424 11779 -9381
rect 11821 -9349 11939 -9306
rect 11821 -9381 11864 -9349
rect 11864 -9381 11896 -9349
rect 11896 -9381 11939 -9349
rect 11821 -9424 11939 -9381
rect 11981 -9349 12099 -9306
rect 11981 -9381 12024 -9349
rect 12024 -9381 12056 -9349
rect 12056 -9381 12099 -9349
rect 11981 -9424 12099 -9381
rect 12141 -9349 12259 -9306
rect 12141 -9381 12184 -9349
rect 12184 -9381 12216 -9349
rect 12216 -9381 12259 -9349
rect 12141 -9424 12259 -9381
rect 12301 -9349 12419 -9306
rect 12301 -9381 12344 -9349
rect 12344 -9381 12376 -9349
rect 12376 -9381 12419 -9349
rect 12301 -9424 12419 -9381
rect 12461 -9349 12579 -9306
rect 12461 -9381 12504 -9349
rect 12504 -9381 12536 -9349
rect 12536 -9381 12579 -9349
rect 12461 -9424 12579 -9381
rect 12621 -9349 12739 -9306
rect 12809 -9319 12927 -9276
rect 12621 -9381 12664 -9349
rect 12664 -9381 12696 -9349
rect 12696 -9381 12739 -9349
rect 12621 -9424 12739 -9381
rect 15261 -5621 15379 -5578
rect 15261 -5653 15304 -5621
rect 15304 -5653 15336 -5621
rect 15336 -5653 15379 -5621
rect 15076 -5724 15194 -5681
rect 15261 -5696 15379 -5653
rect 15421 -5621 15539 -5578
rect 15421 -5653 15464 -5621
rect 15464 -5653 15496 -5621
rect 15496 -5653 15539 -5621
rect 15421 -5696 15539 -5653
rect 15581 -5621 15699 -5578
rect 15581 -5653 15624 -5621
rect 15624 -5653 15656 -5621
rect 15656 -5653 15699 -5621
rect 15581 -5696 15699 -5653
rect 15741 -5621 15859 -5578
rect 15741 -5653 15784 -5621
rect 15784 -5653 15816 -5621
rect 15816 -5653 15859 -5621
rect 15741 -5696 15859 -5653
rect 15901 -5621 16019 -5578
rect 15901 -5653 15944 -5621
rect 15944 -5653 15976 -5621
rect 15976 -5653 16019 -5621
rect 15901 -5696 16019 -5653
rect 16061 -5621 16179 -5578
rect 16061 -5653 16104 -5621
rect 16104 -5653 16136 -5621
rect 16136 -5653 16179 -5621
rect 16061 -5696 16179 -5653
rect 16221 -5621 16339 -5578
rect 16221 -5653 16264 -5621
rect 16264 -5653 16296 -5621
rect 16296 -5653 16339 -5621
rect 16221 -5696 16339 -5653
rect 16381 -5621 16499 -5578
rect 16381 -5653 16424 -5621
rect 16424 -5653 16456 -5621
rect 16456 -5653 16499 -5621
rect 16381 -5696 16499 -5653
rect 16541 -5621 16659 -5578
rect 16541 -5653 16584 -5621
rect 16584 -5653 16616 -5621
rect 16616 -5653 16659 -5621
rect 16541 -5696 16659 -5653
rect 16701 -5621 16819 -5578
rect 16701 -5653 16744 -5621
rect 16744 -5653 16776 -5621
rect 16776 -5653 16819 -5621
rect 16701 -5696 16819 -5653
rect 16861 -5621 16979 -5578
rect 16861 -5653 16904 -5621
rect 16904 -5653 16936 -5621
rect 16936 -5653 16979 -5621
rect 16861 -5696 16979 -5653
rect 17021 -5621 17139 -5578
rect 17021 -5653 17064 -5621
rect 17064 -5653 17096 -5621
rect 17096 -5653 17139 -5621
rect 17021 -5696 17139 -5653
rect 17181 -5621 17299 -5578
rect 17181 -5653 17224 -5621
rect 17224 -5653 17256 -5621
rect 17256 -5653 17299 -5621
rect 17181 -5696 17299 -5653
rect 17341 -5621 17459 -5578
rect 17341 -5653 17384 -5621
rect 17384 -5653 17416 -5621
rect 17416 -5653 17459 -5621
rect 17341 -5696 17459 -5653
rect 17501 -5621 17619 -5578
rect 17501 -5653 17544 -5621
rect 17544 -5653 17576 -5621
rect 17576 -5653 17619 -5621
rect 17501 -5696 17619 -5653
rect 17661 -5621 17779 -5578
rect 17661 -5653 17704 -5621
rect 17704 -5653 17736 -5621
rect 17736 -5653 17779 -5621
rect 17661 -5696 17779 -5653
rect 17821 -5621 17939 -5578
rect 17821 -5653 17864 -5621
rect 17864 -5653 17896 -5621
rect 17896 -5653 17939 -5621
rect 17821 -5696 17939 -5653
rect 17981 -5621 18099 -5578
rect 17981 -5653 18024 -5621
rect 18024 -5653 18056 -5621
rect 18056 -5653 18099 -5621
rect 17981 -5696 18099 -5653
rect 18141 -5621 18259 -5578
rect 18141 -5653 18184 -5621
rect 18184 -5653 18216 -5621
rect 18216 -5653 18259 -5621
rect 18141 -5696 18259 -5653
rect 18301 -5621 18419 -5578
rect 18301 -5653 18344 -5621
rect 18344 -5653 18376 -5621
rect 18376 -5653 18419 -5621
rect 18301 -5696 18419 -5653
rect 18461 -5621 18579 -5578
rect 18461 -5653 18504 -5621
rect 18504 -5653 18536 -5621
rect 18536 -5653 18579 -5621
rect 18461 -5696 18579 -5653
rect 18621 -5621 18739 -5578
rect 18621 -5653 18664 -5621
rect 18664 -5653 18696 -5621
rect 18696 -5653 18739 -5621
rect 18621 -5696 18739 -5653
rect 15076 -5756 15119 -5724
rect 15119 -5756 15151 -5724
rect 15151 -5756 15194 -5724
rect 15076 -5799 15194 -5756
rect 18809 -5724 18927 -5681
rect 18809 -5756 18852 -5724
rect 18852 -5756 18884 -5724
rect 18884 -5756 18927 -5724
rect 15076 -5884 15194 -5841
rect 15076 -5916 15119 -5884
rect 15119 -5916 15151 -5884
rect 15151 -5916 15194 -5884
rect 15076 -5959 15194 -5916
rect 15076 -6044 15194 -6001
rect 15076 -6076 15119 -6044
rect 15119 -6076 15151 -6044
rect 15151 -6076 15194 -6044
rect 15076 -6119 15194 -6076
rect 15076 -6204 15194 -6161
rect 15076 -6236 15119 -6204
rect 15119 -6236 15151 -6204
rect 15151 -6236 15194 -6204
rect 15076 -6279 15194 -6236
rect 15076 -6364 15194 -6321
rect 15076 -6396 15119 -6364
rect 15119 -6396 15151 -6364
rect 15151 -6396 15194 -6364
rect 15076 -6439 15194 -6396
rect 15076 -6524 15194 -6481
rect 15076 -6556 15119 -6524
rect 15119 -6556 15151 -6524
rect 15151 -6556 15194 -6524
rect 15076 -6599 15194 -6556
rect 15076 -6684 15194 -6641
rect 15076 -6716 15119 -6684
rect 15119 -6716 15151 -6684
rect 15151 -6716 15194 -6684
rect 15076 -6759 15194 -6716
rect 15076 -6844 15194 -6801
rect 15076 -6876 15119 -6844
rect 15119 -6876 15151 -6844
rect 15151 -6876 15194 -6844
rect 15076 -6919 15194 -6876
rect 15076 -7004 15194 -6961
rect 15076 -7036 15119 -7004
rect 15119 -7036 15151 -7004
rect 15151 -7036 15194 -7004
rect 15076 -7079 15194 -7036
rect 15076 -7164 15194 -7121
rect 15076 -7196 15119 -7164
rect 15119 -7196 15151 -7164
rect 15151 -7196 15194 -7164
rect 15076 -7239 15194 -7196
rect 15076 -7324 15194 -7281
rect 15076 -7356 15119 -7324
rect 15119 -7356 15151 -7324
rect 15151 -7356 15194 -7324
rect 15076 -7399 15194 -7356
rect 15076 -7484 15194 -7441
rect 15076 -7516 15119 -7484
rect 15119 -7516 15151 -7484
rect 15151 -7516 15194 -7484
rect 15076 -7559 15194 -7516
rect 15076 -7644 15194 -7601
rect 15076 -7676 15119 -7644
rect 15119 -7676 15151 -7644
rect 15151 -7676 15194 -7644
rect 15076 -7719 15194 -7676
rect 15076 -7804 15194 -7761
rect 15076 -7836 15119 -7804
rect 15119 -7836 15151 -7804
rect 15151 -7836 15194 -7804
rect 15076 -7879 15194 -7836
rect 15076 -7964 15194 -7921
rect 15076 -7996 15119 -7964
rect 15119 -7996 15151 -7964
rect 15151 -7996 15194 -7964
rect 15076 -8039 15194 -7996
rect 15076 -8124 15194 -8081
rect 15076 -8156 15119 -8124
rect 15119 -8156 15151 -8124
rect 15151 -8156 15194 -8124
rect 15076 -8199 15194 -8156
rect 15076 -8284 15194 -8241
rect 15076 -8316 15119 -8284
rect 15119 -8316 15151 -8284
rect 15151 -8316 15194 -8284
rect 15076 -8359 15194 -8316
rect 15076 -8444 15194 -8401
rect 15076 -8476 15119 -8444
rect 15119 -8476 15151 -8444
rect 15151 -8476 15194 -8444
rect 15076 -8519 15194 -8476
rect 15076 -8604 15194 -8561
rect 15076 -8636 15119 -8604
rect 15119 -8636 15151 -8604
rect 15151 -8636 15194 -8604
rect 15076 -8679 15194 -8636
rect 15076 -8764 15194 -8721
rect 15076 -8796 15119 -8764
rect 15119 -8796 15151 -8764
rect 15151 -8796 15194 -8764
rect 15076 -8839 15194 -8796
rect 15076 -8924 15194 -8881
rect 15076 -8956 15119 -8924
rect 15119 -8956 15151 -8924
rect 15151 -8956 15194 -8924
rect 15076 -8999 15194 -8956
rect 15076 -9084 15194 -9041
rect 15076 -9116 15119 -9084
rect 15119 -9116 15151 -9084
rect 15151 -9116 15194 -9084
rect 15076 -9159 15194 -9116
rect 15076 -9244 15194 -9201
rect 18809 -5799 18927 -5756
rect 21261 -5621 21379 -5578
rect 21261 -5653 21304 -5621
rect 21304 -5653 21336 -5621
rect 21336 -5653 21379 -5621
rect 21076 -5724 21194 -5681
rect 21261 -5696 21379 -5653
rect 21421 -5621 21539 -5578
rect 21421 -5653 21464 -5621
rect 21464 -5653 21496 -5621
rect 21496 -5653 21539 -5621
rect 21421 -5696 21539 -5653
rect 21581 -5621 21699 -5578
rect 21581 -5653 21624 -5621
rect 21624 -5653 21656 -5621
rect 21656 -5653 21699 -5621
rect 21581 -5696 21699 -5653
rect 21741 -5621 21859 -5578
rect 21741 -5653 21784 -5621
rect 21784 -5653 21816 -5621
rect 21816 -5653 21859 -5621
rect 21741 -5696 21859 -5653
rect 21901 -5621 22019 -5578
rect 21901 -5653 21944 -5621
rect 21944 -5653 21976 -5621
rect 21976 -5653 22019 -5621
rect 21901 -5696 22019 -5653
rect 22061 -5621 22179 -5578
rect 22061 -5653 22104 -5621
rect 22104 -5653 22136 -5621
rect 22136 -5653 22179 -5621
rect 22061 -5696 22179 -5653
rect 22221 -5621 22339 -5578
rect 22221 -5653 22264 -5621
rect 22264 -5653 22296 -5621
rect 22296 -5653 22339 -5621
rect 22221 -5696 22339 -5653
rect 22381 -5621 22499 -5578
rect 22381 -5653 22424 -5621
rect 22424 -5653 22456 -5621
rect 22456 -5653 22499 -5621
rect 22381 -5696 22499 -5653
rect 22541 -5621 22659 -5578
rect 22541 -5653 22584 -5621
rect 22584 -5653 22616 -5621
rect 22616 -5653 22659 -5621
rect 22541 -5696 22659 -5653
rect 22701 -5621 22819 -5578
rect 22701 -5653 22744 -5621
rect 22744 -5653 22776 -5621
rect 22776 -5653 22819 -5621
rect 22701 -5696 22819 -5653
rect 22861 -5621 22979 -5578
rect 22861 -5653 22904 -5621
rect 22904 -5653 22936 -5621
rect 22936 -5653 22979 -5621
rect 22861 -5696 22979 -5653
rect 23021 -5621 23139 -5578
rect 23021 -5653 23064 -5621
rect 23064 -5653 23096 -5621
rect 23096 -5653 23139 -5621
rect 23021 -5696 23139 -5653
rect 23181 -5621 23299 -5578
rect 23181 -5653 23224 -5621
rect 23224 -5653 23256 -5621
rect 23256 -5653 23299 -5621
rect 23181 -5696 23299 -5653
rect 23341 -5621 23459 -5578
rect 23341 -5653 23384 -5621
rect 23384 -5653 23416 -5621
rect 23416 -5653 23459 -5621
rect 23341 -5696 23459 -5653
rect 23501 -5621 23619 -5578
rect 23501 -5653 23544 -5621
rect 23544 -5653 23576 -5621
rect 23576 -5653 23619 -5621
rect 23501 -5696 23619 -5653
rect 23661 -5621 23779 -5578
rect 23661 -5653 23704 -5621
rect 23704 -5653 23736 -5621
rect 23736 -5653 23779 -5621
rect 23661 -5696 23779 -5653
rect 23821 -5621 23939 -5578
rect 23821 -5653 23864 -5621
rect 23864 -5653 23896 -5621
rect 23896 -5653 23939 -5621
rect 23821 -5696 23939 -5653
rect 23981 -5621 24099 -5578
rect 23981 -5653 24024 -5621
rect 24024 -5653 24056 -5621
rect 24056 -5653 24099 -5621
rect 23981 -5696 24099 -5653
rect 24141 -5621 24259 -5578
rect 24141 -5653 24184 -5621
rect 24184 -5653 24216 -5621
rect 24216 -5653 24259 -5621
rect 24141 -5696 24259 -5653
rect 24301 -5621 24419 -5578
rect 24301 -5653 24344 -5621
rect 24344 -5653 24376 -5621
rect 24376 -5653 24419 -5621
rect 24301 -5696 24419 -5653
rect 24461 -5621 24579 -5578
rect 24461 -5653 24504 -5621
rect 24504 -5653 24536 -5621
rect 24536 -5653 24579 -5621
rect 24461 -5696 24579 -5653
rect 24621 -5621 24739 -5578
rect 24621 -5653 24664 -5621
rect 24664 -5653 24696 -5621
rect 24696 -5653 24739 -5621
rect 24621 -5696 24739 -5653
rect 18809 -5884 18927 -5841
rect 18809 -5916 18852 -5884
rect 18852 -5916 18884 -5884
rect 18884 -5916 18927 -5884
rect 18809 -5959 18927 -5916
rect 18809 -6044 18927 -6001
rect 18809 -6076 18852 -6044
rect 18852 -6076 18884 -6044
rect 18884 -6076 18927 -6044
rect 18809 -6119 18927 -6076
rect 18809 -6204 18927 -6161
rect 18809 -6236 18852 -6204
rect 18852 -6236 18884 -6204
rect 18884 -6236 18927 -6204
rect 18809 -6279 18927 -6236
rect 18809 -6364 18927 -6321
rect 18809 -6396 18852 -6364
rect 18852 -6396 18884 -6364
rect 18884 -6396 18927 -6364
rect 18809 -6439 18927 -6396
rect 18809 -6524 18927 -6481
rect 18809 -6556 18852 -6524
rect 18852 -6556 18884 -6524
rect 18884 -6556 18927 -6524
rect 18809 -6599 18927 -6556
rect 18809 -6684 18927 -6641
rect 18809 -6716 18852 -6684
rect 18852 -6716 18884 -6684
rect 18884 -6716 18927 -6684
rect 18809 -6759 18927 -6716
rect 18809 -6844 18927 -6801
rect 18809 -6876 18852 -6844
rect 18852 -6876 18884 -6844
rect 18884 -6876 18927 -6844
rect 18809 -6919 18927 -6876
rect 18809 -7004 18927 -6961
rect 18809 -7036 18852 -7004
rect 18852 -7036 18884 -7004
rect 18884 -7036 18927 -7004
rect 18809 -7079 18927 -7036
rect 18809 -7164 18927 -7121
rect 18809 -7196 18852 -7164
rect 18852 -7196 18884 -7164
rect 18884 -7196 18927 -7164
rect 18809 -7239 18927 -7196
rect 18809 -7324 18927 -7281
rect 18809 -7356 18852 -7324
rect 18852 -7356 18884 -7324
rect 18884 -7356 18927 -7324
rect 18809 -7399 18927 -7356
rect 18809 -7484 18927 -7441
rect 18809 -7516 18852 -7484
rect 18852 -7516 18884 -7484
rect 18884 -7516 18927 -7484
rect 18809 -7559 18927 -7516
rect 18809 -7644 18927 -7601
rect 18809 -7676 18852 -7644
rect 18852 -7676 18884 -7644
rect 18884 -7676 18927 -7644
rect 18809 -7719 18927 -7676
rect 18809 -7804 18927 -7761
rect 18809 -7836 18852 -7804
rect 18852 -7836 18884 -7804
rect 18884 -7836 18927 -7804
rect 18809 -7879 18927 -7836
rect 18809 -7964 18927 -7921
rect 18809 -7996 18852 -7964
rect 18852 -7996 18884 -7964
rect 18884 -7996 18927 -7964
rect 18809 -8039 18927 -7996
rect 18809 -8124 18927 -8081
rect 18809 -8156 18852 -8124
rect 18852 -8156 18884 -8124
rect 18884 -8156 18927 -8124
rect 18809 -8199 18927 -8156
rect 18809 -8284 18927 -8241
rect 18809 -8316 18852 -8284
rect 18852 -8316 18884 -8284
rect 18884 -8316 18927 -8284
rect 18809 -8359 18927 -8316
rect 18809 -8444 18927 -8401
rect 18809 -8476 18852 -8444
rect 18852 -8476 18884 -8444
rect 18884 -8476 18927 -8444
rect 18809 -8519 18927 -8476
rect 18809 -8604 18927 -8561
rect 18809 -8636 18852 -8604
rect 18852 -8636 18884 -8604
rect 18884 -8636 18927 -8604
rect 18809 -8679 18927 -8636
rect 18809 -8764 18927 -8721
rect 18809 -8796 18852 -8764
rect 18852 -8796 18884 -8764
rect 18884 -8796 18927 -8764
rect 18809 -8839 18927 -8796
rect 18809 -8924 18927 -8881
rect 18809 -8956 18852 -8924
rect 18852 -8956 18884 -8924
rect 18884 -8956 18927 -8924
rect 18809 -8999 18927 -8956
rect 18809 -9084 18927 -9041
rect 18809 -9116 18852 -9084
rect 18852 -9116 18884 -9084
rect 18884 -9116 18927 -9084
rect 18809 -9159 18927 -9116
rect 15076 -9276 15119 -9244
rect 15119 -9276 15151 -9244
rect 15151 -9276 15194 -9244
rect 15076 -9319 15194 -9276
rect 18809 -9244 18927 -9201
rect 18809 -9276 18852 -9244
rect 18852 -9276 18884 -9244
rect 18884 -9276 18927 -9244
rect 15261 -9349 15379 -9306
rect 15261 -9381 15304 -9349
rect 15304 -9381 15336 -9349
rect 15336 -9381 15379 -9349
rect 15261 -9424 15379 -9381
rect 15421 -9349 15539 -9306
rect 15421 -9381 15464 -9349
rect 15464 -9381 15496 -9349
rect 15496 -9381 15539 -9349
rect 15421 -9424 15539 -9381
rect 15581 -9349 15699 -9306
rect 15581 -9381 15624 -9349
rect 15624 -9381 15656 -9349
rect 15656 -9381 15699 -9349
rect 15581 -9424 15699 -9381
rect 15741 -9349 15859 -9306
rect 15741 -9381 15784 -9349
rect 15784 -9381 15816 -9349
rect 15816 -9381 15859 -9349
rect 15741 -9424 15859 -9381
rect 15901 -9349 16019 -9306
rect 15901 -9381 15944 -9349
rect 15944 -9381 15976 -9349
rect 15976 -9381 16019 -9349
rect 15901 -9424 16019 -9381
rect 16061 -9349 16179 -9306
rect 16061 -9381 16104 -9349
rect 16104 -9381 16136 -9349
rect 16136 -9381 16179 -9349
rect 16061 -9424 16179 -9381
rect 16221 -9349 16339 -9306
rect 16221 -9381 16264 -9349
rect 16264 -9381 16296 -9349
rect 16296 -9381 16339 -9349
rect 16221 -9424 16339 -9381
rect 16381 -9349 16499 -9306
rect 16381 -9381 16424 -9349
rect 16424 -9381 16456 -9349
rect 16456 -9381 16499 -9349
rect 16381 -9424 16499 -9381
rect 16541 -9349 16659 -9306
rect 16541 -9381 16584 -9349
rect 16584 -9381 16616 -9349
rect 16616 -9381 16659 -9349
rect 16541 -9424 16659 -9381
rect 16701 -9349 16819 -9306
rect 16701 -9381 16744 -9349
rect 16744 -9381 16776 -9349
rect 16776 -9381 16819 -9349
rect 16701 -9424 16819 -9381
rect 16861 -9349 16979 -9306
rect 16861 -9381 16904 -9349
rect 16904 -9381 16936 -9349
rect 16936 -9381 16979 -9349
rect 16861 -9424 16979 -9381
rect 17021 -9349 17139 -9306
rect 17021 -9381 17064 -9349
rect 17064 -9381 17096 -9349
rect 17096 -9381 17139 -9349
rect 17021 -9424 17139 -9381
rect 17181 -9349 17299 -9306
rect 17181 -9381 17224 -9349
rect 17224 -9381 17256 -9349
rect 17256 -9381 17299 -9349
rect 17181 -9424 17299 -9381
rect 17341 -9349 17459 -9306
rect 17341 -9381 17384 -9349
rect 17384 -9381 17416 -9349
rect 17416 -9381 17459 -9349
rect 17341 -9424 17459 -9381
rect 17501 -9349 17619 -9306
rect 17501 -9381 17544 -9349
rect 17544 -9381 17576 -9349
rect 17576 -9381 17619 -9349
rect 17501 -9424 17619 -9381
rect 17661 -9349 17779 -9306
rect 17661 -9381 17704 -9349
rect 17704 -9381 17736 -9349
rect 17736 -9381 17779 -9349
rect 17661 -9424 17779 -9381
rect 17821 -9349 17939 -9306
rect 17821 -9381 17864 -9349
rect 17864 -9381 17896 -9349
rect 17896 -9381 17939 -9349
rect 17821 -9424 17939 -9381
rect 17981 -9349 18099 -9306
rect 17981 -9381 18024 -9349
rect 18024 -9381 18056 -9349
rect 18056 -9381 18099 -9349
rect 17981 -9424 18099 -9381
rect 18141 -9349 18259 -9306
rect 18141 -9381 18184 -9349
rect 18184 -9381 18216 -9349
rect 18216 -9381 18259 -9349
rect 18141 -9424 18259 -9381
rect 18301 -9349 18419 -9306
rect 18301 -9381 18344 -9349
rect 18344 -9381 18376 -9349
rect 18376 -9381 18419 -9349
rect 18301 -9424 18419 -9381
rect 18461 -9349 18579 -9306
rect 18461 -9381 18504 -9349
rect 18504 -9381 18536 -9349
rect 18536 -9381 18579 -9349
rect 18461 -9424 18579 -9381
rect 18621 -9349 18739 -9306
rect 18809 -9319 18927 -9276
rect 18621 -9381 18664 -9349
rect 18664 -9381 18696 -9349
rect 18696 -9381 18739 -9349
rect 18621 -9424 18739 -9381
rect 21076 -5756 21119 -5724
rect 21119 -5756 21151 -5724
rect 21151 -5756 21194 -5724
rect 21076 -5799 21194 -5756
rect 24809 -5724 24927 -5681
rect 24809 -5756 24852 -5724
rect 24852 -5756 24884 -5724
rect 24884 -5756 24927 -5724
rect 21076 -5884 21194 -5841
rect 21076 -5916 21119 -5884
rect 21119 -5916 21151 -5884
rect 21151 -5916 21194 -5884
rect 21076 -5959 21194 -5916
rect 21076 -6044 21194 -6001
rect 21076 -6076 21119 -6044
rect 21119 -6076 21151 -6044
rect 21151 -6076 21194 -6044
rect 21076 -6119 21194 -6076
rect 21076 -6204 21194 -6161
rect 21076 -6236 21119 -6204
rect 21119 -6236 21151 -6204
rect 21151 -6236 21194 -6204
rect 21076 -6279 21194 -6236
rect 21076 -6364 21194 -6321
rect 21076 -6396 21119 -6364
rect 21119 -6396 21151 -6364
rect 21151 -6396 21194 -6364
rect 21076 -6439 21194 -6396
rect 21076 -6524 21194 -6481
rect 21076 -6556 21119 -6524
rect 21119 -6556 21151 -6524
rect 21151 -6556 21194 -6524
rect 21076 -6599 21194 -6556
rect 21076 -6684 21194 -6641
rect 21076 -6716 21119 -6684
rect 21119 -6716 21151 -6684
rect 21151 -6716 21194 -6684
rect 21076 -6759 21194 -6716
rect 21076 -6844 21194 -6801
rect 21076 -6876 21119 -6844
rect 21119 -6876 21151 -6844
rect 21151 -6876 21194 -6844
rect 21076 -6919 21194 -6876
rect 21076 -7004 21194 -6961
rect 21076 -7036 21119 -7004
rect 21119 -7036 21151 -7004
rect 21151 -7036 21194 -7004
rect 21076 -7079 21194 -7036
rect 21076 -7164 21194 -7121
rect 21076 -7196 21119 -7164
rect 21119 -7196 21151 -7164
rect 21151 -7196 21194 -7164
rect 21076 -7239 21194 -7196
rect 21076 -7324 21194 -7281
rect 21076 -7356 21119 -7324
rect 21119 -7356 21151 -7324
rect 21151 -7356 21194 -7324
rect 21076 -7399 21194 -7356
rect 21076 -7484 21194 -7441
rect 21076 -7516 21119 -7484
rect 21119 -7516 21151 -7484
rect 21151 -7516 21194 -7484
rect 21076 -7559 21194 -7516
rect 21076 -7644 21194 -7601
rect 21076 -7676 21119 -7644
rect 21119 -7676 21151 -7644
rect 21151 -7676 21194 -7644
rect 21076 -7719 21194 -7676
rect 21076 -7804 21194 -7761
rect 21076 -7836 21119 -7804
rect 21119 -7836 21151 -7804
rect 21151 -7836 21194 -7804
rect 21076 -7879 21194 -7836
rect 21076 -7964 21194 -7921
rect 21076 -7996 21119 -7964
rect 21119 -7996 21151 -7964
rect 21151 -7996 21194 -7964
rect 21076 -8039 21194 -7996
rect 21076 -8124 21194 -8081
rect 21076 -8156 21119 -8124
rect 21119 -8156 21151 -8124
rect 21151 -8156 21194 -8124
rect 21076 -8199 21194 -8156
rect 21076 -8284 21194 -8241
rect 21076 -8316 21119 -8284
rect 21119 -8316 21151 -8284
rect 21151 -8316 21194 -8284
rect 21076 -8359 21194 -8316
rect 21076 -8444 21194 -8401
rect 21076 -8476 21119 -8444
rect 21119 -8476 21151 -8444
rect 21151 -8476 21194 -8444
rect 21076 -8519 21194 -8476
rect 21076 -8604 21194 -8561
rect 21076 -8636 21119 -8604
rect 21119 -8636 21151 -8604
rect 21151 -8636 21194 -8604
rect 21076 -8679 21194 -8636
rect 21076 -8764 21194 -8721
rect 21076 -8796 21119 -8764
rect 21119 -8796 21151 -8764
rect 21151 -8796 21194 -8764
rect 21076 -8839 21194 -8796
rect 21076 -8924 21194 -8881
rect 21076 -8956 21119 -8924
rect 21119 -8956 21151 -8924
rect 21151 -8956 21194 -8924
rect 21076 -8999 21194 -8956
rect 21076 -9084 21194 -9041
rect 21076 -9116 21119 -9084
rect 21119 -9116 21151 -9084
rect 21151 -9116 21194 -9084
rect 21076 -9159 21194 -9116
rect 21076 -9244 21194 -9201
rect 24809 -5799 24927 -5756
rect 24809 -5884 24927 -5841
rect 24809 -5916 24852 -5884
rect 24852 -5916 24884 -5884
rect 24884 -5916 24927 -5884
rect 24809 -5959 24927 -5916
rect 24809 -6044 24927 -6001
rect 24809 -6076 24852 -6044
rect 24852 -6076 24884 -6044
rect 24884 -6076 24927 -6044
rect 24809 -6119 24927 -6076
rect 24809 -6204 24927 -6161
rect 24809 -6236 24852 -6204
rect 24852 -6236 24884 -6204
rect 24884 -6236 24927 -6204
rect 24809 -6279 24927 -6236
rect 24809 -6364 24927 -6321
rect 24809 -6396 24852 -6364
rect 24852 -6396 24884 -6364
rect 24884 -6396 24927 -6364
rect 24809 -6439 24927 -6396
rect 24809 -6524 24927 -6481
rect 24809 -6556 24852 -6524
rect 24852 -6556 24884 -6524
rect 24884 -6556 24927 -6524
rect 24809 -6599 24927 -6556
rect 24809 -6684 24927 -6641
rect 24809 -6716 24852 -6684
rect 24852 -6716 24884 -6684
rect 24884 -6716 24927 -6684
rect 24809 -6759 24927 -6716
rect 24809 -6844 24927 -6801
rect 24809 -6876 24852 -6844
rect 24852 -6876 24884 -6844
rect 24884 -6876 24927 -6844
rect 24809 -6919 24927 -6876
rect 24809 -7004 24927 -6961
rect 24809 -7036 24852 -7004
rect 24852 -7036 24884 -7004
rect 24884 -7036 24927 -7004
rect 24809 -7079 24927 -7036
rect 24809 -7164 24927 -7121
rect 24809 -7196 24852 -7164
rect 24852 -7196 24884 -7164
rect 24884 -7196 24927 -7164
rect 24809 -7239 24927 -7196
rect 24809 -7324 24927 -7281
rect 24809 -7356 24852 -7324
rect 24852 -7356 24884 -7324
rect 24884 -7356 24927 -7324
rect 24809 -7399 24927 -7356
rect 24809 -7484 24927 -7441
rect 24809 -7516 24852 -7484
rect 24852 -7516 24884 -7484
rect 24884 -7516 24927 -7484
rect 24809 -7559 24927 -7516
rect 24809 -7644 24927 -7601
rect 24809 -7676 24852 -7644
rect 24852 -7676 24884 -7644
rect 24884 -7676 24927 -7644
rect 24809 -7719 24927 -7676
rect 24809 -7804 24927 -7761
rect 24809 -7836 24852 -7804
rect 24852 -7836 24884 -7804
rect 24884 -7836 24927 -7804
rect 24809 -7879 24927 -7836
rect 24809 -7964 24927 -7921
rect 24809 -7996 24852 -7964
rect 24852 -7996 24884 -7964
rect 24884 -7996 24927 -7964
rect 24809 -8039 24927 -7996
rect 24809 -8124 24927 -8081
rect 24809 -8156 24852 -8124
rect 24852 -8156 24884 -8124
rect 24884 -8156 24927 -8124
rect 24809 -8199 24927 -8156
rect 24809 -8284 24927 -8241
rect 24809 -8316 24852 -8284
rect 24852 -8316 24884 -8284
rect 24884 -8316 24927 -8284
rect 24809 -8359 24927 -8316
rect 24809 -8444 24927 -8401
rect 24809 -8476 24852 -8444
rect 24852 -8476 24884 -8444
rect 24884 -8476 24927 -8444
rect 24809 -8519 24927 -8476
rect 24809 -8604 24927 -8561
rect 24809 -8636 24852 -8604
rect 24852 -8636 24884 -8604
rect 24884 -8636 24927 -8604
rect 24809 -8679 24927 -8636
rect 24809 -8764 24927 -8721
rect 24809 -8796 24852 -8764
rect 24852 -8796 24884 -8764
rect 24884 -8796 24927 -8764
rect 24809 -8839 24927 -8796
rect 24809 -8924 24927 -8881
rect 24809 -8956 24852 -8924
rect 24852 -8956 24884 -8924
rect 24884 -8956 24927 -8924
rect 24809 -8999 24927 -8956
rect 24809 -9084 24927 -9041
rect 24809 -9116 24852 -9084
rect 24852 -9116 24884 -9084
rect 24884 -9116 24927 -9084
rect 24809 -9159 24927 -9116
rect 21076 -9276 21119 -9244
rect 21119 -9276 21151 -9244
rect 21151 -9276 21194 -9244
rect 21076 -9319 21194 -9276
rect 24809 -9244 24927 -9201
rect 24809 -9276 24852 -9244
rect 24852 -9276 24884 -9244
rect 24884 -9276 24927 -9244
rect 21261 -9349 21379 -9306
rect 21261 -9381 21304 -9349
rect 21304 -9381 21336 -9349
rect 21336 -9381 21379 -9349
rect 21261 -9424 21379 -9381
rect 21421 -9349 21539 -9306
rect 21421 -9381 21464 -9349
rect 21464 -9381 21496 -9349
rect 21496 -9381 21539 -9349
rect 21421 -9424 21539 -9381
rect 21581 -9349 21699 -9306
rect 21581 -9381 21624 -9349
rect 21624 -9381 21656 -9349
rect 21656 -9381 21699 -9349
rect 21581 -9424 21699 -9381
rect 21741 -9349 21859 -9306
rect 21741 -9381 21784 -9349
rect 21784 -9381 21816 -9349
rect 21816 -9381 21859 -9349
rect 21741 -9424 21859 -9381
rect 21901 -9349 22019 -9306
rect 21901 -9381 21944 -9349
rect 21944 -9381 21976 -9349
rect 21976 -9381 22019 -9349
rect 21901 -9424 22019 -9381
rect 22061 -9349 22179 -9306
rect 22061 -9381 22104 -9349
rect 22104 -9381 22136 -9349
rect 22136 -9381 22179 -9349
rect 22061 -9424 22179 -9381
rect 22221 -9349 22339 -9306
rect 22221 -9381 22264 -9349
rect 22264 -9381 22296 -9349
rect 22296 -9381 22339 -9349
rect 22221 -9424 22339 -9381
rect 22381 -9349 22499 -9306
rect 22381 -9381 22424 -9349
rect 22424 -9381 22456 -9349
rect 22456 -9381 22499 -9349
rect 22381 -9424 22499 -9381
rect 22541 -9349 22659 -9306
rect 22541 -9381 22584 -9349
rect 22584 -9381 22616 -9349
rect 22616 -9381 22659 -9349
rect 22541 -9424 22659 -9381
rect 22701 -9349 22819 -9306
rect 22701 -9381 22744 -9349
rect 22744 -9381 22776 -9349
rect 22776 -9381 22819 -9349
rect 22701 -9424 22819 -9381
rect 22861 -9349 22979 -9306
rect 22861 -9381 22904 -9349
rect 22904 -9381 22936 -9349
rect 22936 -9381 22979 -9349
rect 22861 -9424 22979 -9381
rect 23021 -9349 23139 -9306
rect 23021 -9381 23064 -9349
rect 23064 -9381 23096 -9349
rect 23096 -9381 23139 -9349
rect 23021 -9424 23139 -9381
rect 23181 -9349 23299 -9306
rect 23181 -9381 23224 -9349
rect 23224 -9381 23256 -9349
rect 23256 -9381 23299 -9349
rect 23181 -9424 23299 -9381
rect 23341 -9349 23459 -9306
rect 23341 -9381 23384 -9349
rect 23384 -9381 23416 -9349
rect 23416 -9381 23459 -9349
rect 23341 -9424 23459 -9381
rect 23501 -9349 23619 -9306
rect 23501 -9381 23544 -9349
rect 23544 -9381 23576 -9349
rect 23576 -9381 23619 -9349
rect 23501 -9424 23619 -9381
rect 23661 -9349 23779 -9306
rect 23661 -9381 23704 -9349
rect 23704 -9381 23736 -9349
rect 23736 -9381 23779 -9349
rect 23661 -9424 23779 -9381
rect 23821 -9349 23939 -9306
rect 23821 -9381 23864 -9349
rect 23864 -9381 23896 -9349
rect 23896 -9381 23939 -9349
rect 23821 -9424 23939 -9381
rect 23981 -9349 24099 -9306
rect 23981 -9381 24024 -9349
rect 24024 -9381 24056 -9349
rect 24056 -9381 24099 -9349
rect 23981 -9424 24099 -9381
rect 24141 -9349 24259 -9306
rect 24141 -9381 24184 -9349
rect 24184 -9381 24216 -9349
rect 24216 -9381 24259 -9349
rect 24141 -9424 24259 -9381
rect 24301 -9349 24419 -9306
rect 24301 -9381 24344 -9349
rect 24344 -9381 24376 -9349
rect 24376 -9381 24419 -9349
rect 24301 -9424 24419 -9381
rect 24461 -9349 24579 -9306
rect 24461 -9381 24504 -9349
rect 24504 -9381 24536 -9349
rect 24536 -9381 24579 -9349
rect 24461 -9424 24579 -9381
rect 24621 -9349 24739 -9306
rect 24809 -9319 24927 -9276
rect 24621 -9381 24664 -9349
rect 24664 -9381 24696 -9349
rect 24696 -9381 24739 -9349
rect 24621 -9424 24739 -9381
rect 3261 -11621 3379 -11578
rect 3261 -11653 3304 -11621
rect 3304 -11653 3336 -11621
rect 3336 -11653 3379 -11621
rect 3076 -11724 3194 -11681
rect 3261 -11696 3379 -11653
rect 3421 -11621 3539 -11578
rect 3421 -11653 3464 -11621
rect 3464 -11653 3496 -11621
rect 3496 -11653 3539 -11621
rect 3421 -11696 3539 -11653
rect 3581 -11621 3699 -11578
rect 3581 -11653 3624 -11621
rect 3624 -11653 3656 -11621
rect 3656 -11653 3699 -11621
rect 3581 -11696 3699 -11653
rect 3741 -11621 3859 -11578
rect 3741 -11653 3784 -11621
rect 3784 -11653 3816 -11621
rect 3816 -11653 3859 -11621
rect 3741 -11696 3859 -11653
rect 3901 -11621 4019 -11578
rect 3901 -11653 3944 -11621
rect 3944 -11653 3976 -11621
rect 3976 -11653 4019 -11621
rect 3901 -11696 4019 -11653
rect 4061 -11621 4179 -11578
rect 4061 -11653 4104 -11621
rect 4104 -11653 4136 -11621
rect 4136 -11653 4179 -11621
rect 4061 -11696 4179 -11653
rect 4221 -11621 4339 -11578
rect 4221 -11653 4264 -11621
rect 4264 -11653 4296 -11621
rect 4296 -11653 4339 -11621
rect 4221 -11696 4339 -11653
rect 4381 -11621 4499 -11578
rect 4381 -11653 4424 -11621
rect 4424 -11653 4456 -11621
rect 4456 -11653 4499 -11621
rect 4381 -11696 4499 -11653
rect 4541 -11621 4659 -11578
rect 4541 -11653 4584 -11621
rect 4584 -11653 4616 -11621
rect 4616 -11653 4659 -11621
rect 4541 -11696 4659 -11653
rect 4701 -11621 4819 -11578
rect 4701 -11653 4744 -11621
rect 4744 -11653 4776 -11621
rect 4776 -11653 4819 -11621
rect 4701 -11696 4819 -11653
rect 4861 -11621 4979 -11578
rect 4861 -11653 4904 -11621
rect 4904 -11653 4936 -11621
rect 4936 -11653 4979 -11621
rect 4861 -11696 4979 -11653
rect 5021 -11621 5139 -11578
rect 5021 -11653 5064 -11621
rect 5064 -11653 5096 -11621
rect 5096 -11653 5139 -11621
rect 5021 -11696 5139 -11653
rect 5181 -11621 5299 -11578
rect 5181 -11653 5224 -11621
rect 5224 -11653 5256 -11621
rect 5256 -11653 5299 -11621
rect 5181 -11696 5299 -11653
rect 5341 -11621 5459 -11578
rect 5341 -11653 5384 -11621
rect 5384 -11653 5416 -11621
rect 5416 -11653 5459 -11621
rect 5341 -11696 5459 -11653
rect 5501 -11621 5619 -11578
rect 5501 -11653 5544 -11621
rect 5544 -11653 5576 -11621
rect 5576 -11653 5619 -11621
rect 5501 -11696 5619 -11653
rect 5661 -11621 5779 -11578
rect 5661 -11653 5704 -11621
rect 5704 -11653 5736 -11621
rect 5736 -11653 5779 -11621
rect 5661 -11696 5779 -11653
rect 5821 -11621 5939 -11578
rect 5821 -11653 5864 -11621
rect 5864 -11653 5896 -11621
rect 5896 -11653 5939 -11621
rect 5821 -11696 5939 -11653
rect 5981 -11621 6099 -11578
rect 5981 -11653 6024 -11621
rect 6024 -11653 6056 -11621
rect 6056 -11653 6099 -11621
rect 5981 -11696 6099 -11653
rect 6141 -11621 6259 -11578
rect 6141 -11653 6184 -11621
rect 6184 -11653 6216 -11621
rect 6216 -11653 6259 -11621
rect 6141 -11696 6259 -11653
rect 6301 -11621 6419 -11578
rect 6301 -11653 6344 -11621
rect 6344 -11653 6376 -11621
rect 6376 -11653 6419 -11621
rect 6301 -11696 6419 -11653
rect 6461 -11621 6579 -11578
rect 6461 -11653 6504 -11621
rect 6504 -11653 6536 -11621
rect 6536 -11653 6579 -11621
rect 6461 -11696 6579 -11653
rect 6621 -11621 6739 -11578
rect 6621 -11653 6664 -11621
rect 6664 -11653 6696 -11621
rect 6696 -11653 6739 -11621
rect 6621 -11696 6739 -11653
rect 3076 -11756 3119 -11724
rect 3119 -11756 3151 -11724
rect 3151 -11756 3194 -11724
rect 3076 -11799 3194 -11756
rect 6809 -11724 6927 -11681
rect 6809 -11756 6852 -11724
rect 6852 -11756 6884 -11724
rect 6884 -11756 6927 -11724
rect 3076 -11884 3194 -11841
rect 3076 -11916 3119 -11884
rect 3119 -11916 3151 -11884
rect 3151 -11916 3194 -11884
rect 3076 -11959 3194 -11916
rect 3076 -12044 3194 -12001
rect 3076 -12076 3119 -12044
rect 3119 -12076 3151 -12044
rect 3151 -12076 3194 -12044
rect 3076 -12119 3194 -12076
rect 3076 -12204 3194 -12161
rect 3076 -12236 3119 -12204
rect 3119 -12236 3151 -12204
rect 3151 -12236 3194 -12204
rect 3076 -12279 3194 -12236
rect 3076 -12364 3194 -12321
rect 3076 -12396 3119 -12364
rect 3119 -12396 3151 -12364
rect 3151 -12396 3194 -12364
rect 3076 -12439 3194 -12396
rect 3076 -12524 3194 -12481
rect 3076 -12556 3119 -12524
rect 3119 -12556 3151 -12524
rect 3151 -12556 3194 -12524
rect 3076 -12599 3194 -12556
rect 3076 -12684 3194 -12641
rect 3076 -12716 3119 -12684
rect 3119 -12716 3151 -12684
rect 3151 -12716 3194 -12684
rect 3076 -12759 3194 -12716
rect 3076 -12844 3194 -12801
rect 3076 -12876 3119 -12844
rect 3119 -12876 3151 -12844
rect 3151 -12876 3194 -12844
rect 3076 -12919 3194 -12876
rect 3076 -13004 3194 -12961
rect 3076 -13036 3119 -13004
rect 3119 -13036 3151 -13004
rect 3151 -13036 3194 -13004
rect 3076 -13079 3194 -13036
rect 3076 -13164 3194 -13121
rect 3076 -13196 3119 -13164
rect 3119 -13196 3151 -13164
rect 3151 -13196 3194 -13164
rect 3076 -13239 3194 -13196
rect 3076 -13324 3194 -13281
rect 3076 -13356 3119 -13324
rect 3119 -13356 3151 -13324
rect 3151 -13356 3194 -13324
rect 3076 -13399 3194 -13356
rect 3076 -13484 3194 -13441
rect 3076 -13516 3119 -13484
rect 3119 -13516 3151 -13484
rect 3151 -13516 3194 -13484
rect 3076 -13559 3194 -13516
rect 3076 -13644 3194 -13601
rect 3076 -13676 3119 -13644
rect 3119 -13676 3151 -13644
rect 3151 -13676 3194 -13644
rect 3076 -13719 3194 -13676
rect 3076 -13804 3194 -13761
rect 3076 -13836 3119 -13804
rect 3119 -13836 3151 -13804
rect 3151 -13836 3194 -13804
rect 3076 -13879 3194 -13836
rect 3076 -13964 3194 -13921
rect 3076 -13996 3119 -13964
rect 3119 -13996 3151 -13964
rect 3151 -13996 3194 -13964
rect 3076 -14039 3194 -13996
rect 3076 -14124 3194 -14081
rect 3076 -14156 3119 -14124
rect 3119 -14156 3151 -14124
rect 3151 -14156 3194 -14124
rect 3076 -14199 3194 -14156
rect 3076 -14284 3194 -14241
rect 3076 -14316 3119 -14284
rect 3119 -14316 3151 -14284
rect 3151 -14316 3194 -14284
rect 3076 -14359 3194 -14316
rect 3076 -14444 3194 -14401
rect 3076 -14476 3119 -14444
rect 3119 -14476 3151 -14444
rect 3151 -14476 3194 -14444
rect 3076 -14519 3194 -14476
rect 3076 -14604 3194 -14561
rect 3076 -14636 3119 -14604
rect 3119 -14636 3151 -14604
rect 3151 -14636 3194 -14604
rect 3076 -14679 3194 -14636
rect 3076 -14764 3194 -14721
rect 3076 -14796 3119 -14764
rect 3119 -14796 3151 -14764
rect 3151 -14796 3194 -14764
rect 3076 -14839 3194 -14796
rect 3076 -14924 3194 -14881
rect 3076 -14956 3119 -14924
rect 3119 -14956 3151 -14924
rect 3151 -14956 3194 -14924
rect 3076 -14999 3194 -14956
rect 3076 -15084 3194 -15041
rect 3076 -15116 3119 -15084
rect 3119 -15116 3151 -15084
rect 3151 -15116 3194 -15084
rect 3076 -15159 3194 -15116
rect 3076 -15244 3194 -15201
rect 6809 -11799 6927 -11756
rect 6809 -11884 6927 -11841
rect 6809 -11916 6852 -11884
rect 6852 -11916 6884 -11884
rect 6884 -11916 6927 -11884
rect 6809 -11959 6927 -11916
rect 6809 -12044 6927 -12001
rect 6809 -12076 6852 -12044
rect 6852 -12076 6884 -12044
rect 6884 -12076 6927 -12044
rect 6809 -12119 6927 -12076
rect 6809 -12204 6927 -12161
rect 6809 -12236 6852 -12204
rect 6852 -12236 6884 -12204
rect 6884 -12236 6927 -12204
rect 6809 -12279 6927 -12236
rect 6809 -12364 6927 -12321
rect 6809 -12396 6852 -12364
rect 6852 -12396 6884 -12364
rect 6884 -12396 6927 -12364
rect 6809 -12439 6927 -12396
rect 6809 -12524 6927 -12481
rect 6809 -12556 6852 -12524
rect 6852 -12556 6884 -12524
rect 6884 -12556 6927 -12524
rect 6809 -12599 6927 -12556
rect 6809 -12684 6927 -12641
rect 6809 -12716 6852 -12684
rect 6852 -12716 6884 -12684
rect 6884 -12716 6927 -12684
rect 6809 -12759 6927 -12716
rect 6809 -12844 6927 -12801
rect 6809 -12876 6852 -12844
rect 6852 -12876 6884 -12844
rect 6884 -12876 6927 -12844
rect 6809 -12919 6927 -12876
rect 6809 -13004 6927 -12961
rect 6809 -13036 6852 -13004
rect 6852 -13036 6884 -13004
rect 6884 -13036 6927 -13004
rect 6809 -13079 6927 -13036
rect 6809 -13164 6927 -13121
rect 6809 -13196 6852 -13164
rect 6852 -13196 6884 -13164
rect 6884 -13196 6927 -13164
rect 6809 -13239 6927 -13196
rect 6809 -13324 6927 -13281
rect 6809 -13356 6852 -13324
rect 6852 -13356 6884 -13324
rect 6884 -13356 6927 -13324
rect 6809 -13399 6927 -13356
rect 6809 -13484 6927 -13441
rect 6809 -13516 6852 -13484
rect 6852 -13516 6884 -13484
rect 6884 -13516 6927 -13484
rect 6809 -13559 6927 -13516
rect 6809 -13644 6927 -13601
rect 6809 -13676 6852 -13644
rect 6852 -13676 6884 -13644
rect 6884 -13676 6927 -13644
rect 6809 -13719 6927 -13676
rect 6809 -13804 6927 -13761
rect 6809 -13836 6852 -13804
rect 6852 -13836 6884 -13804
rect 6884 -13836 6927 -13804
rect 6809 -13879 6927 -13836
rect 6809 -13964 6927 -13921
rect 6809 -13996 6852 -13964
rect 6852 -13996 6884 -13964
rect 6884 -13996 6927 -13964
rect 6809 -14039 6927 -13996
rect 6809 -14124 6927 -14081
rect 6809 -14156 6852 -14124
rect 6852 -14156 6884 -14124
rect 6884 -14156 6927 -14124
rect 6809 -14199 6927 -14156
rect 6809 -14284 6927 -14241
rect 6809 -14316 6852 -14284
rect 6852 -14316 6884 -14284
rect 6884 -14316 6927 -14284
rect 6809 -14359 6927 -14316
rect 6809 -14444 6927 -14401
rect 6809 -14476 6852 -14444
rect 6852 -14476 6884 -14444
rect 6884 -14476 6927 -14444
rect 6809 -14519 6927 -14476
rect 6809 -14604 6927 -14561
rect 6809 -14636 6852 -14604
rect 6852 -14636 6884 -14604
rect 6884 -14636 6927 -14604
rect 6809 -14679 6927 -14636
rect 6809 -14764 6927 -14721
rect 6809 -14796 6852 -14764
rect 6852 -14796 6884 -14764
rect 6884 -14796 6927 -14764
rect 6809 -14839 6927 -14796
rect 6809 -14924 6927 -14881
rect 6809 -14956 6852 -14924
rect 6852 -14956 6884 -14924
rect 6884 -14956 6927 -14924
rect 6809 -14999 6927 -14956
rect 6809 -15084 6927 -15041
rect 6809 -15116 6852 -15084
rect 6852 -15116 6884 -15084
rect 6884 -15116 6927 -15084
rect 6809 -15159 6927 -15116
rect 3076 -15276 3119 -15244
rect 3119 -15276 3151 -15244
rect 3151 -15276 3194 -15244
rect 3076 -15319 3194 -15276
rect 6809 -15244 6927 -15201
rect 6809 -15276 6852 -15244
rect 6852 -15276 6884 -15244
rect 6884 -15276 6927 -15244
rect 3261 -15349 3379 -15306
rect 3261 -15381 3304 -15349
rect 3304 -15381 3336 -15349
rect 3336 -15381 3379 -15349
rect 3261 -15424 3379 -15381
rect 3421 -15349 3539 -15306
rect 3421 -15381 3464 -15349
rect 3464 -15381 3496 -15349
rect 3496 -15381 3539 -15349
rect 3421 -15424 3539 -15381
rect 3581 -15349 3699 -15306
rect 3581 -15381 3624 -15349
rect 3624 -15381 3656 -15349
rect 3656 -15381 3699 -15349
rect 3581 -15424 3699 -15381
rect 3741 -15349 3859 -15306
rect 3741 -15381 3784 -15349
rect 3784 -15381 3816 -15349
rect 3816 -15381 3859 -15349
rect 3741 -15424 3859 -15381
rect 3901 -15349 4019 -15306
rect 3901 -15381 3944 -15349
rect 3944 -15381 3976 -15349
rect 3976 -15381 4019 -15349
rect 3901 -15424 4019 -15381
rect 4061 -15349 4179 -15306
rect 4061 -15381 4104 -15349
rect 4104 -15381 4136 -15349
rect 4136 -15381 4179 -15349
rect 4061 -15424 4179 -15381
rect 4221 -15349 4339 -15306
rect 4221 -15381 4264 -15349
rect 4264 -15381 4296 -15349
rect 4296 -15381 4339 -15349
rect 4221 -15424 4339 -15381
rect 4381 -15349 4499 -15306
rect 4381 -15381 4424 -15349
rect 4424 -15381 4456 -15349
rect 4456 -15381 4499 -15349
rect 4381 -15424 4499 -15381
rect 4541 -15349 4659 -15306
rect 4541 -15381 4584 -15349
rect 4584 -15381 4616 -15349
rect 4616 -15381 4659 -15349
rect 4541 -15424 4659 -15381
rect 4701 -15349 4819 -15306
rect 4701 -15381 4744 -15349
rect 4744 -15381 4776 -15349
rect 4776 -15381 4819 -15349
rect 4701 -15424 4819 -15381
rect 4861 -15349 4979 -15306
rect 4861 -15381 4904 -15349
rect 4904 -15381 4936 -15349
rect 4936 -15381 4979 -15349
rect 4861 -15424 4979 -15381
rect 5021 -15349 5139 -15306
rect 5021 -15381 5064 -15349
rect 5064 -15381 5096 -15349
rect 5096 -15381 5139 -15349
rect 5021 -15424 5139 -15381
rect 5181 -15349 5299 -15306
rect 5181 -15381 5224 -15349
rect 5224 -15381 5256 -15349
rect 5256 -15381 5299 -15349
rect 5181 -15424 5299 -15381
rect 5341 -15349 5459 -15306
rect 5341 -15381 5384 -15349
rect 5384 -15381 5416 -15349
rect 5416 -15381 5459 -15349
rect 5341 -15424 5459 -15381
rect 5501 -15349 5619 -15306
rect 5501 -15381 5544 -15349
rect 5544 -15381 5576 -15349
rect 5576 -15381 5619 -15349
rect 5501 -15424 5619 -15381
rect 5661 -15349 5779 -15306
rect 5661 -15381 5704 -15349
rect 5704 -15381 5736 -15349
rect 5736 -15381 5779 -15349
rect 5661 -15424 5779 -15381
rect 5821 -15349 5939 -15306
rect 5821 -15381 5864 -15349
rect 5864 -15381 5896 -15349
rect 5896 -15381 5939 -15349
rect 5821 -15424 5939 -15381
rect 5981 -15349 6099 -15306
rect 5981 -15381 6024 -15349
rect 6024 -15381 6056 -15349
rect 6056 -15381 6099 -15349
rect 5981 -15424 6099 -15381
rect 6141 -15349 6259 -15306
rect 6141 -15381 6184 -15349
rect 6184 -15381 6216 -15349
rect 6216 -15381 6259 -15349
rect 6141 -15424 6259 -15381
rect 6301 -15349 6419 -15306
rect 6301 -15381 6344 -15349
rect 6344 -15381 6376 -15349
rect 6376 -15381 6419 -15349
rect 6301 -15424 6419 -15381
rect 6461 -15349 6579 -15306
rect 6461 -15381 6504 -15349
rect 6504 -15381 6536 -15349
rect 6536 -15381 6579 -15349
rect 6461 -15424 6579 -15381
rect 6621 -15349 6739 -15306
rect 6809 -15319 6927 -15276
rect 6621 -15381 6664 -15349
rect 6664 -15381 6696 -15349
rect 6696 -15381 6739 -15349
rect 6621 -15424 6739 -15381
rect 9261 -11621 9379 -11578
rect 9261 -11653 9304 -11621
rect 9304 -11653 9336 -11621
rect 9336 -11653 9379 -11621
rect 9076 -11724 9194 -11681
rect 9261 -11696 9379 -11653
rect 9421 -11621 9539 -11578
rect 9421 -11653 9464 -11621
rect 9464 -11653 9496 -11621
rect 9496 -11653 9539 -11621
rect 9421 -11696 9539 -11653
rect 9581 -11621 9699 -11578
rect 9581 -11653 9624 -11621
rect 9624 -11653 9656 -11621
rect 9656 -11653 9699 -11621
rect 9581 -11696 9699 -11653
rect 9741 -11621 9859 -11578
rect 9741 -11653 9784 -11621
rect 9784 -11653 9816 -11621
rect 9816 -11653 9859 -11621
rect 9741 -11696 9859 -11653
rect 9901 -11621 10019 -11578
rect 9901 -11653 9944 -11621
rect 9944 -11653 9976 -11621
rect 9976 -11653 10019 -11621
rect 9901 -11696 10019 -11653
rect 10061 -11621 10179 -11578
rect 10061 -11653 10104 -11621
rect 10104 -11653 10136 -11621
rect 10136 -11653 10179 -11621
rect 10061 -11696 10179 -11653
rect 10221 -11621 10339 -11578
rect 10221 -11653 10264 -11621
rect 10264 -11653 10296 -11621
rect 10296 -11653 10339 -11621
rect 10221 -11696 10339 -11653
rect 10381 -11621 10499 -11578
rect 10381 -11653 10424 -11621
rect 10424 -11653 10456 -11621
rect 10456 -11653 10499 -11621
rect 10381 -11696 10499 -11653
rect 10541 -11621 10659 -11578
rect 10541 -11653 10584 -11621
rect 10584 -11653 10616 -11621
rect 10616 -11653 10659 -11621
rect 10541 -11696 10659 -11653
rect 10701 -11621 10819 -11578
rect 10701 -11653 10744 -11621
rect 10744 -11653 10776 -11621
rect 10776 -11653 10819 -11621
rect 10701 -11696 10819 -11653
rect 10861 -11621 10979 -11578
rect 10861 -11653 10904 -11621
rect 10904 -11653 10936 -11621
rect 10936 -11653 10979 -11621
rect 10861 -11696 10979 -11653
rect 11021 -11621 11139 -11578
rect 11021 -11653 11064 -11621
rect 11064 -11653 11096 -11621
rect 11096 -11653 11139 -11621
rect 11021 -11696 11139 -11653
rect 11181 -11621 11299 -11578
rect 11181 -11653 11224 -11621
rect 11224 -11653 11256 -11621
rect 11256 -11653 11299 -11621
rect 11181 -11696 11299 -11653
rect 11341 -11621 11459 -11578
rect 11341 -11653 11384 -11621
rect 11384 -11653 11416 -11621
rect 11416 -11653 11459 -11621
rect 11341 -11696 11459 -11653
rect 11501 -11621 11619 -11578
rect 11501 -11653 11544 -11621
rect 11544 -11653 11576 -11621
rect 11576 -11653 11619 -11621
rect 11501 -11696 11619 -11653
rect 11661 -11621 11779 -11578
rect 11661 -11653 11704 -11621
rect 11704 -11653 11736 -11621
rect 11736 -11653 11779 -11621
rect 11661 -11696 11779 -11653
rect 11821 -11621 11939 -11578
rect 11821 -11653 11864 -11621
rect 11864 -11653 11896 -11621
rect 11896 -11653 11939 -11621
rect 11821 -11696 11939 -11653
rect 11981 -11621 12099 -11578
rect 11981 -11653 12024 -11621
rect 12024 -11653 12056 -11621
rect 12056 -11653 12099 -11621
rect 11981 -11696 12099 -11653
rect 12141 -11621 12259 -11578
rect 12141 -11653 12184 -11621
rect 12184 -11653 12216 -11621
rect 12216 -11653 12259 -11621
rect 12141 -11696 12259 -11653
rect 12301 -11621 12419 -11578
rect 12301 -11653 12344 -11621
rect 12344 -11653 12376 -11621
rect 12376 -11653 12419 -11621
rect 12301 -11696 12419 -11653
rect 12461 -11621 12579 -11578
rect 12461 -11653 12504 -11621
rect 12504 -11653 12536 -11621
rect 12536 -11653 12579 -11621
rect 12461 -11696 12579 -11653
rect 12621 -11621 12739 -11578
rect 12621 -11653 12664 -11621
rect 12664 -11653 12696 -11621
rect 12696 -11653 12739 -11621
rect 12621 -11696 12739 -11653
rect 9076 -11756 9119 -11724
rect 9119 -11756 9151 -11724
rect 9151 -11756 9194 -11724
rect 9076 -11799 9194 -11756
rect 12809 -11724 12927 -11681
rect 12809 -11756 12852 -11724
rect 12852 -11756 12884 -11724
rect 12884 -11756 12927 -11724
rect 9076 -11884 9194 -11841
rect 9076 -11916 9119 -11884
rect 9119 -11916 9151 -11884
rect 9151 -11916 9194 -11884
rect 9076 -11959 9194 -11916
rect 9076 -12044 9194 -12001
rect 9076 -12076 9119 -12044
rect 9119 -12076 9151 -12044
rect 9151 -12076 9194 -12044
rect 9076 -12119 9194 -12076
rect 9076 -12204 9194 -12161
rect 9076 -12236 9119 -12204
rect 9119 -12236 9151 -12204
rect 9151 -12236 9194 -12204
rect 9076 -12279 9194 -12236
rect 9076 -12364 9194 -12321
rect 9076 -12396 9119 -12364
rect 9119 -12396 9151 -12364
rect 9151 -12396 9194 -12364
rect 9076 -12439 9194 -12396
rect 9076 -12524 9194 -12481
rect 9076 -12556 9119 -12524
rect 9119 -12556 9151 -12524
rect 9151 -12556 9194 -12524
rect 9076 -12599 9194 -12556
rect 9076 -12684 9194 -12641
rect 9076 -12716 9119 -12684
rect 9119 -12716 9151 -12684
rect 9151 -12716 9194 -12684
rect 9076 -12759 9194 -12716
rect 9076 -12844 9194 -12801
rect 9076 -12876 9119 -12844
rect 9119 -12876 9151 -12844
rect 9151 -12876 9194 -12844
rect 9076 -12919 9194 -12876
rect 9076 -13004 9194 -12961
rect 9076 -13036 9119 -13004
rect 9119 -13036 9151 -13004
rect 9151 -13036 9194 -13004
rect 9076 -13079 9194 -13036
rect 9076 -13164 9194 -13121
rect 9076 -13196 9119 -13164
rect 9119 -13196 9151 -13164
rect 9151 -13196 9194 -13164
rect 9076 -13239 9194 -13196
rect 9076 -13324 9194 -13281
rect 9076 -13356 9119 -13324
rect 9119 -13356 9151 -13324
rect 9151 -13356 9194 -13324
rect 9076 -13399 9194 -13356
rect 9076 -13484 9194 -13441
rect 9076 -13516 9119 -13484
rect 9119 -13516 9151 -13484
rect 9151 -13516 9194 -13484
rect 9076 -13559 9194 -13516
rect 9076 -13644 9194 -13601
rect 9076 -13676 9119 -13644
rect 9119 -13676 9151 -13644
rect 9151 -13676 9194 -13644
rect 9076 -13719 9194 -13676
rect 9076 -13804 9194 -13761
rect 9076 -13836 9119 -13804
rect 9119 -13836 9151 -13804
rect 9151 -13836 9194 -13804
rect 9076 -13879 9194 -13836
rect 9076 -13964 9194 -13921
rect 9076 -13996 9119 -13964
rect 9119 -13996 9151 -13964
rect 9151 -13996 9194 -13964
rect 9076 -14039 9194 -13996
rect 9076 -14124 9194 -14081
rect 9076 -14156 9119 -14124
rect 9119 -14156 9151 -14124
rect 9151 -14156 9194 -14124
rect 9076 -14199 9194 -14156
rect 9076 -14284 9194 -14241
rect 9076 -14316 9119 -14284
rect 9119 -14316 9151 -14284
rect 9151 -14316 9194 -14284
rect 9076 -14359 9194 -14316
rect 9076 -14444 9194 -14401
rect 9076 -14476 9119 -14444
rect 9119 -14476 9151 -14444
rect 9151 -14476 9194 -14444
rect 9076 -14519 9194 -14476
rect 9076 -14604 9194 -14561
rect 9076 -14636 9119 -14604
rect 9119 -14636 9151 -14604
rect 9151 -14636 9194 -14604
rect 9076 -14679 9194 -14636
rect 9076 -14764 9194 -14721
rect 9076 -14796 9119 -14764
rect 9119 -14796 9151 -14764
rect 9151 -14796 9194 -14764
rect 9076 -14839 9194 -14796
rect 9076 -14924 9194 -14881
rect 9076 -14956 9119 -14924
rect 9119 -14956 9151 -14924
rect 9151 -14956 9194 -14924
rect 9076 -14999 9194 -14956
rect 9076 -15084 9194 -15041
rect 9076 -15116 9119 -15084
rect 9119 -15116 9151 -15084
rect 9151 -15116 9194 -15084
rect 9076 -15159 9194 -15116
rect 9076 -15244 9194 -15201
rect 12809 -11799 12927 -11756
rect 12809 -11884 12927 -11841
rect 12809 -11916 12852 -11884
rect 12852 -11916 12884 -11884
rect 12884 -11916 12927 -11884
rect 12809 -11959 12927 -11916
rect 12809 -12044 12927 -12001
rect 12809 -12076 12852 -12044
rect 12852 -12076 12884 -12044
rect 12884 -12076 12927 -12044
rect 12809 -12119 12927 -12076
rect 12809 -12204 12927 -12161
rect 12809 -12236 12852 -12204
rect 12852 -12236 12884 -12204
rect 12884 -12236 12927 -12204
rect 12809 -12279 12927 -12236
rect 12809 -12364 12927 -12321
rect 12809 -12396 12852 -12364
rect 12852 -12396 12884 -12364
rect 12884 -12396 12927 -12364
rect 12809 -12439 12927 -12396
rect 12809 -12524 12927 -12481
rect 12809 -12556 12852 -12524
rect 12852 -12556 12884 -12524
rect 12884 -12556 12927 -12524
rect 12809 -12599 12927 -12556
rect 12809 -12684 12927 -12641
rect 12809 -12716 12852 -12684
rect 12852 -12716 12884 -12684
rect 12884 -12716 12927 -12684
rect 12809 -12759 12927 -12716
rect 12809 -12844 12927 -12801
rect 12809 -12876 12852 -12844
rect 12852 -12876 12884 -12844
rect 12884 -12876 12927 -12844
rect 12809 -12919 12927 -12876
rect 12809 -13004 12927 -12961
rect 12809 -13036 12852 -13004
rect 12852 -13036 12884 -13004
rect 12884 -13036 12927 -13004
rect 12809 -13079 12927 -13036
rect 12809 -13164 12927 -13121
rect 12809 -13196 12852 -13164
rect 12852 -13196 12884 -13164
rect 12884 -13196 12927 -13164
rect 12809 -13239 12927 -13196
rect 12809 -13324 12927 -13281
rect 12809 -13356 12852 -13324
rect 12852 -13356 12884 -13324
rect 12884 -13356 12927 -13324
rect 12809 -13399 12927 -13356
rect 12809 -13484 12927 -13441
rect 12809 -13516 12852 -13484
rect 12852 -13516 12884 -13484
rect 12884 -13516 12927 -13484
rect 12809 -13559 12927 -13516
rect 12809 -13644 12927 -13601
rect 12809 -13676 12852 -13644
rect 12852 -13676 12884 -13644
rect 12884 -13676 12927 -13644
rect 12809 -13719 12927 -13676
rect 12809 -13804 12927 -13761
rect 12809 -13836 12852 -13804
rect 12852 -13836 12884 -13804
rect 12884 -13836 12927 -13804
rect 12809 -13879 12927 -13836
rect 12809 -13964 12927 -13921
rect 12809 -13996 12852 -13964
rect 12852 -13996 12884 -13964
rect 12884 -13996 12927 -13964
rect 12809 -14039 12927 -13996
rect 12809 -14124 12927 -14081
rect 12809 -14156 12852 -14124
rect 12852 -14156 12884 -14124
rect 12884 -14156 12927 -14124
rect 12809 -14199 12927 -14156
rect 12809 -14284 12927 -14241
rect 12809 -14316 12852 -14284
rect 12852 -14316 12884 -14284
rect 12884 -14316 12927 -14284
rect 12809 -14359 12927 -14316
rect 12809 -14444 12927 -14401
rect 12809 -14476 12852 -14444
rect 12852 -14476 12884 -14444
rect 12884 -14476 12927 -14444
rect 12809 -14519 12927 -14476
rect 12809 -14604 12927 -14561
rect 12809 -14636 12852 -14604
rect 12852 -14636 12884 -14604
rect 12884 -14636 12927 -14604
rect 12809 -14679 12927 -14636
rect 12809 -14764 12927 -14721
rect 12809 -14796 12852 -14764
rect 12852 -14796 12884 -14764
rect 12884 -14796 12927 -14764
rect 12809 -14839 12927 -14796
rect 12809 -14924 12927 -14881
rect 12809 -14956 12852 -14924
rect 12852 -14956 12884 -14924
rect 12884 -14956 12927 -14924
rect 12809 -14999 12927 -14956
rect 12809 -15084 12927 -15041
rect 12809 -15116 12852 -15084
rect 12852 -15116 12884 -15084
rect 12884 -15116 12927 -15084
rect 12809 -15159 12927 -15116
rect 9076 -15276 9119 -15244
rect 9119 -15276 9151 -15244
rect 9151 -15276 9194 -15244
rect 9076 -15319 9194 -15276
rect 12809 -15244 12927 -15201
rect 12809 -15276 12852 -15244
rect 12852 -15276 12884 -15244
rect 12884 -15276 12927 -15244
rect 9261 -15349 9379 -15306
rect 9261 -15381 9304 -15349
rect 9304 -15381 9336 -15349
rect 9336 -15381 9379 -15349
rect 9261 -15424 9379 -15381
rect 9421 -15349 9539 -15306
rect 9421 -15381 9464 -15349
rect 9464 -15381 9496 -15349
rect 9496 -15381 9539 -15349
rect 9421 -15424 9539 -15381
rect 9581 -15349 9699 -15306
rect 9581 -15381 9624 -15349
rect 9624 -15381 9656 -15349
rect 9656 -15381 9699 -15349
rect 9581 -15424 9699 -15381
rect 9741 -15349 9859 -15306
rect 9741 -15381 9784 -15349
rect 9784 -15381 9816 -15349
rect 9816 -15381 9859 -15349
rect 9741 -15424 9859 -15381
rect 9901 -15349 10019 -15306
rect 9901 -15381 9944 -15349
rect 9944 -15381 9976 -15349
rect 9976 -15381 10019 -15349
rect 9901 -15424 10019 -15381
rect 10061 -15349 10179 -15306
rect 10061 -15381 10104 -15349
rect 10104 -15381 10136 -15349
rect 10136 -15381 10179 -15349
rect 10061 -15424 10179 -15381
rect 10221 -15349 10339 -15306
rect 10221 -15381 10264 -15349
rect 10264 -15381 10296 -15349
rect 10296 -15381 10339 -15349
rect 10221 -15424 10339 -15381
rect 10381 -15349 10499 -15306
rect 10381 -15381 10424 -15349
rect 10424 -15381 10456 -15349
rect 10456 -15381 10499 -15349
rect 10381 -15424 10499 -15381
rect 10541 -15349 10659 -15306
rect 10541 -15381 10584 -15349
rect 10584 -15381 10616 -15349
rect 10616 -15381 10659 -15349
rect 10541 -15424 10659 -15381
rect 10701 -15349 10819 -15306
rect 10701 -15381 10744 -15349
rect 10744 -15381 10776 -15349
rect 10776 -15381 10819 -15349
rect 10701 -15424 10819 -15381
rect 10861 -15349 10979 -15306
rect 10861 -15381 10904 -15349
rect 10904 -15381 10936 -15349
rect 10936 -15381 10979 -15349
rect 10861 -15424 10979 -15381
rect 11021 -15349 11139 -15306
rect 11021 -15381 11064 -15349
rect 11064 -15381 11096 -15349
rect 11096 -15381 11139 -15349
rect 11021 -15424 11139 -15381
rect 11181 -15349 11299 -15306
rect 11181 -15381 11224 -15349
rect 11224 -15381 11256 -15349
rect 11256 -15381 11299 -15349
rect 11181 -15424 11299 -15381
rect 11341 -15349 11459 -15306
rect 11341 -15381 11384 -15349
rect 11384 -15381 11416 -15349
rect 11416 -15381 11459 -15349
rect 11341 -15424 11459 -15381
rect 11501 -15349 11619 -15306
rect 11501 -15381 11544 -15349
rect 11544 -15381 11576 -15349
rect 11576 -15381 11619 -15349
rect 11501 -15424 11619 -15381
rect 11661 -15349 11779 -15306
rect 11661 -15381 11704 -15349
rect 11704 -15381 11736 -15349
rect 11736 -15381 11779 -15349
rect 11661 -15424 11779 -15381
rect 11821 -15349 11939 -15306
rect 11821 -15381 11864 -15349
rect 11864 -15381 11896 -15349
rect 11896 -15381 11939 -15349
rect 11821 -15424 11939 -15381
rect 11981 -15349 12099 -15306
rect 11981 -15381 12024 -15349
rect 12024 -15381 12056 -15349
rect 12056 -15381 12099 -15349
rect 11981 -15424 12099 -15381
rect 12141 -15349 12259 -15306
rect 12141 -15381 12184 -15349
rect 12184 -15381 12216 -15349
rect 12216 -15381 12259 -15349
rect 12141 -15424 12259 -15381
rect 12301 -15349 12419 -15306
rect 12301 -15381 12344 -15349
rect 12344 -15381 12376 -15349
rect 12376 -15381 12419 -15349
rect 12301 -15424 12419 -15381
rect 12461 -15349 12579 -15306
rect 12461 -15381 12504 -15349
rect 12504 -15381 12536 -15349
rect 12536 -15381 12579 -15349
rect 12461 -15424 12579 -15381
rect 12621 -15349 12739 -15306
rect 12809 -15319 12927 -15276
rect 12621 -15381 12664 -15349
rect 12664 -15381 12696 -15349
rect 12696 -15381 12739 -15349
rect 12621 -15424 12739 -15381
rect 15261 -11621 15379 -11578
rect 15261 -11653 15304 -11621
rect 15304 -11653 15336 -11621
rect 15336 -11653 15379 -11621
rect 15076 -11724 15194 -11681
rect 15261 -11696 15379 -11653
rect 15421 -11621 15539 -11578
rect 15421 -11653 15464 -11621
rect 15464 -11653 15496 -11621
rect 15496 -11653 15539 -11621
rect 15421 -11696 15539 -11653
rect 15581 -11621 15699 -11578
rect 15581 -11653 15624 -11621
rect 15624 -11653 15656 -11621
rect 15656 -11653 15699 -11621
rect 15581 -11696 15699 -11653
rect 15741 -11621 15859 -11578
rect 15741 -11653 15784 -11621
rect 15784 -11653 15816 -11621
rect 15816 -11653 15859 -11621
rect 15741 -11696 15859 -11653
rect 15901 -11621 16019 -11578
rect 15901 -11653 15944 -11621
rect 15944 -11653 15976 -11621
rect 15976 -11653 16019 -11621
rect 15901 -11696 16019 -11653
rect 16061 -11621 16179 -11578
rect 16061 -11653 16104 -11621
rect 16104 -11653 16136 -11621
rect 16136 -11653 16179 -11621
rect 16061 -11696 16179 -11653
rect 16221 -11621 16339 -11578
rect 16221 -11653 16264 -11621
rect 16264 -11653 16296 -11621
rect 16296 -11653 16339 -11621
rect 16221 -11696 16339 -11653
rect 16381 -11621 16499 -11578
rect 16381 -11653 16424 -11621
rect 16424 -11653 16456 -11621
rect 16456 -11653 16499 -11621
rect 16381 -11696 16499 -11653
rect 16541 -11621 16659 -11578
rect 16541 -11653 16584 -11621
rect 16584 -11653 16616 -11621
rect 16616 -11653 16659 -11621
rect 16541 -11696 16659 -11653
rect 16701 -11621 16819 -11578
rect 16701 -11653 16744 -11621
rect 16744 -11653 16776 -11621
rect 16776 -11653 16819 -11621
rect 16701 -11696 16819 -11653
rect 16861 -11621 16979 -11578
rect 16861 -11653 16904 -11621
rect 16904 -11653 16936 -11621
rect 16936 -11653 16979 -11621
rect 16861 -11696 16979 -11653
rect 17021 -11621 17139 -11578
rect 17021 -11653 17064 -11621
rect 17064 -11653 17096 -11621
rect 17096 -11653 17139 -11621
rect 17021 -11696 17139 -11653
rect 17181 -11621 17299 -11578
rect 17181 -11653 17224 -11621
rect 17224 -11653 17256 -11621
rect 17256 -11653 17299 -11621
rect 17181 -11696 17299 -11653
rect 17341 -11621 17459 -11578
rect 17341 -11653 17384 -11621
rect 17384 -11653 17416 -11621
rect 17416 -11653 17459 -11621
rect 17341 -11696 17459 -11653
rect 17501 -11621 17619 -11578
rect 17501 -11653 17544 -11621
rect 17544 -11653 17576 -11621
rect 17576 -11653 17619 -11621
rect 17501 -11696 17619 -11653
rect 17661 -11621 17779 -11578
rect 17661 -11653 17704 -11621
rect 17704 -11653 17736 -11621
rect 17736 -11653 17779 -11621
rect 17661 -11696 17779 -11653
rect 17821 -11621 17939 -11578
rect 17821 -11653 17864 -11621
rect 17864 -11653 17896 -11621
rect 17896 -11653 17939 -11621
rect 17821 -11696 17939 -11653
rect 17981 -11621 18099 -11578
rect 17981 -11653 18024 -11621
rect 18024 -11653 18056 -11621
rect 18056 -11653 18099 -11621
rect 17981 -11696 18099 -11653
rect 18141 -11621 18259 -11578
rect 18141 -11653 18184 -11621
rect 18184 -11653 18216 -11621
rect 18216 -11653 18259 -11621
rect 18141 -11696 18259 -11653
rect 18301 -11621 18419 -11578
rect 18301 -11653 18344 -11621
rect 18344 -11653 18376 -11621
rect 18376 -11653 18419 -11621
rect 18301 -11696 18419 -11653
rect 18461 -11621 18579 -11578
rect 18461 -11653 18504 -11621
rect 18504 -11653 18536 -11621
rect 18536 -11653 18579 -11621
rect 18461 -11696 18579 -11653
rect 18621 -11621 18739 -11578
rect 18621 -11653 18664 -11621
rect 18664 -11653 18696 -11621
rect 18696 -11653 18739 -11621
rect 18621 -11696 18739 -11653
rect 15076 -11756 15119 -11724
rect 15119 -11756 15151 -11724
rect 15151 -11756 15194 -11724
rect 15076 -11799 15194 -11756
rect 18809 -11724 18927 -11681
rect 18809 -11756 18852 -11724
rect 18852 -11756 18884 -11724
rect 18884 -11756 18927 -11724
rect 15076 -11884 15194 -11841
rect 15076 -11916 15119 -11884
rect 15119 -11916 15151 -11884
rect 15151 -11916 15194 -11884
rect 15076 -11959 15194 -11916
rect 15076 -12044 15194 -12001
rect 15076 -12076 15119 -12044
rect 15119 -12076 15151 -12044
rect 15151 -12076 15194 -12044
rect 15076 -12119 15194 -12076
rect 15076 -12204 15194 -12161
rect 15076 -12236 15119 -12204
rect 15119 -12236 15151 -12204
rect 15151 -12236 15194 -12204
rect 15076 -12279 15194 -12236
rect 15076 -12364 15194 -12321
rect 15076 -12396 15119 -12364
rect 15119 -12396 15151 -12364
rect 15151 -12396 15194 -12364
rect 15076 -12439 15194 -12396
rect 15076 -12524 15194 -12481
rect 15076 -12556 15119 -12524
rect 15119 -12556 15151 -12524
rect 15151 -12556 15194 -12524
rect 15076 -12599 15194 -12556
rect 15076 -12684 15194 -12641
rect 15076 -12716 15119 -12684
rect 15119 -12716 15151 -12684
rect 15151 -12716 15194 -12684
rect 15076 -12759 15194 -12716
rect 15076 -12844 15194 -12801
rect 15076 -12876 15119 -12844
rect 15119 -12876 15151 -12844
rect 15151 -12876 15194 -12844
rect 15076 -12919 15194 -12876
rect 15076 -13004 15194 -12961
rect 15076 -13036 15119 -13004
rect 15119 -13036 15151 -13004
rect 15151 -13036 15194 -13004
rect 15076 -13079 15194 -13036
rect 15076 -13164 15194 -13121
rect 15076 -13196 15119 -13164
rect 15119 -13196 15151 -13164
rect 15151 -13196 15194 -13164
rect 15076 -13239 15194 -13196
rect 15076 -13324 15194 -13281
rect 15076 -13356 15119 -13324
rect 15119 -13356 15151 -13324
rect 15151 -13356 15194 -13324
rect 15076 -13399 15194 -13356
rect 15076 -13484 15194 -13441
rect 15076 -13516 15119 -13484
rect 15119 -13516 15151 -13484
rect 15151 -13516 15194 -13484
rect 15076 -13559 15194 -13516
rect 15076 -13644 15194 -13601
rect 15076 -13676 15119 -13644
rect 15119 -13676 15151 -13644
rect 15151 -13676 15194 -13644
rect 15076 -13719 15194 -13676
rect 15076 -13804 15194 -13761
rect 15076 -13836 15119 -13804
rect 15119 -13836 15151 -13804
rect 15151 -13836 15194 -13804
rect 15076 -13879 15194 -13836
rect 15076 -13964 15194 -13921
rect 15076 -13996 15119 -13964
rect 15119 -13996 15151 -13964
rect 15151 -13996 15194 -13964
rect 15076 -14039 15194 -13996
rect 15076 -14124 15194 -14081
rect 15076 -14156 15119 -14124
rect 15119 -14156 15151 -14124
rect 15151 -14156 15194 -14124
rect 15076 -14199 15194 -14156
rect 15076 -14284 15194 -14241
rect 15076 -14316 15119 -14284
rect 15119 -14316 15151 -14284
rect 15151 -14316 15194 -14284
rect 15076 -14359 15194 -14316
rect 15076 -14444 15194 -14401
rect 15076 -14476 15119 -14444
rect 15119 -14476 15151 -14444
rect 15151 -14476 15194 -14444
rect 15076 -14519 15194 -14476
rect 15076 -14604 15194 -14561
rect 15076 -14636 15119 -14604
rect 15119 -14636 15151 -14604
rect 15151 -14636 15194 -14604
rect 15076 -14679 15194 -14636
rect 15076 -14764 15194 -14721
rect 15076 -14796 15119 -14764
rect 15119 -14796 15151 -14764
rect 15151 -14796 15194 -14764
rect 15076 -14839 15194 -14796
rect 15076 -14924 15194 -14881
rect 15076 -14956 15119 -14924
rect 15119 -14956 15151 -14924
rect 15151 -14956 15194 -14924
rect 15076 -14999 15194 -14956
rect 15076 -15084 15194 -15041
rect 15076 -15116 15119 -15084
rect 15119 -15116 15151 -15084
rect 15151 -15116 15194 -15084
rect 15076 -15159 15194 -15116
rect 15076 -15244 15194 -15201
rect 18809 -11799 18927 -11756
rect 18809 -11884 18927 -11841
rect 18809 -11916 18852 -11884
rect 18852 -11916 18884 -11884
rect 18884 -11916 18927 -11884
rect 18809 -11959 18927 -11916
rect 18809 -12044 18927 -12001
rect 18809 -12076 18852 -12044
rect 18852 -12076 18884 -12044
rect 18884 -12076 18927 -12044
rect 18809 -12119 18927 -12076
rect 18809 -12204 18927 -12161
rect 18809 -12236 18852 -12204
rect 18852 -12236 18884 -12204
rect 18884 -12236 18927 -12204
rect 18809 -12279 18927 -12236
rect 18809 -12364 18927 -12321
rect 18809 -12396 18852 -12364
rect 18852 -12396 18884 -12364
rect 18884 -12396 18927 -12364
rect 18809 -12439 18927 -12396
rect 18809 -12524 18927 -12481
rect 18809 -12556 18852 -12524
rect 18852 -12556 18884 -12524
rect 18884 -12556 18927 -12524
rect 18809 -12599 18927 -12556
rect 18809 -12684 18927 -12641
rect 18809 -12716 18852 -12684
rect 18852 -12716 18884 -12684
rect 18884 -12716 18927 -12684
rect 18809 -12759 18927 -12716
rect 18809 -12844 18927 -12801
rect 18809 -12876 18852 -12844
rect 18852 -12876 18884 -12844
rect 18884 -12876 18927 -12844
rect 18809 -12919 18927 -12876
rect 18809 -13004 18927 -12961
rect 18809 -13036 18852 -13004
rect 18852 -13036 18884 -13004
rect 18884 -13036 18927 -13004
rect 18809 -13079 18927 -13036
rect 18809 -13164 18927 -13121
rect 18809 -13196 18852 -13164
rect 18852 -13196 18884 -13164
rect 18884 -13196 18927 -13164
rect 18809 -13239 18927 -13196
rect 18809 -13324 18927 -13281
rect 18809 -13356 18852 -13324
rect 18852 -13356 18884 -13324
rect 18884 -13356 18927 -13324
rect 18809 -13399 18927 -13356
rect 18809 -13484 18927 -13441
rect 18809 -13516 18852 -13484
rect 18852 -13516 18884 -13484
rect 18884 -13516 18927 -13484
rect 18809 -13559 18927 -13516
rect 18809 -13644 18927 -13601
rect 18809 -13676 18852 -13644
rect 18852 -13676 18884 -13644
rect 18884 -13676 18927 -13644
rect 18809 -13719 18927 -13676
rect 18809 -13804 18927 -13761
rect 18809 -13836 18852 -13804
rect 18852 -13836 18884 -13804
rect 18884 -13836 18927 -13804
rect 18809 -13879 18927 -13836
rect 18809 -13964 18927 -13921
rect 18809 -13996 18852 -13964
rect 18852 -13996 18884 -13964
rect 18884 -13996 18927 -13964
rect 18809 -14039 18927 -13996
rect 18809 -14124 18927 -14081
rect 18809 -14156 18852 -14124
rect 18852 -14156 18884 -14124
rect 18884 -14156 18927 -14124
rect 18809 -14199 18927 -14156
rect 18809 -14284 18927 -14241
rect 18809 -14316 18852 -14284
rect 18852 -14316 18884 -14284
rect 18884 -14316 18927 -14284
rect 18809 -14359 18927 -14316
rect 18809 -14444 18927 -14401
rect 18809 -14476 18852 -14444
rect 18852 -14476 18884 -14444
rect 18884 -14476 18927 -14444
rect 18809 -14519 18927 -14476
rect 18809 -14604 18927 -14561
rect 18809 -14636 18852 -14604
rect 18852 -14636 18884 -14604
rect 18884 -14636 18927 -14604
rect 18809 -14679 18927 -14636
rect 18809 -14764 18927 -14721
rect 18809 -14796 18852 -14764
rect 18852 -14796 18884 -14764
rect 18884 -14796 18927 -14764
rect 18809 -14839 18927 -14796
rect 18809 -14924 18927 -14881
rect 18809 -14956 18852 -14924
rect 18852 -14956 18884 -14924
rect 18884 -14956 18927 -14924
rect 18809 -14999 18927 -14956
rect 18809 -15084 18927 -15041
rect 18809 -15116 18852 -15084
rect 18852 -15116 18884 -15084
rect 18884 -15116 18927 -15084
rect 18809 -15159 18927 -15116
rect 15076 -15276 15119 -15244
rect 15119 -15276 15151 -15244
rect 15151 -15276 15194 -15244
rect 15076 -15319 15194 -15276
rect 18809 -15244 18927 -15201
rect 18809 -15276 18852 -15244
rect 18852 -15276 18884 -15244
rect 18884 -15276 18927 -15244
rect 15261 -15349 15379 -15306
rect 15261 -15381 15304 -15349
rect 15304 -15381 15336 -15349
rect 15336 -15381 15379 -15349
rect 15261 -15424 15379 -15381
rect 15421 -15349 15539 -15306
rect 15421 -15381 15464 -15349
rect 15464 -15381 15496 -15349
rect 15496 -15381 15539 -15349
rect 15421 -15424 15539 -15381
rect 15581 -15349 15699 -15306
rect 15581 -15381 15624 -15349
rect 15624 -15381 15656 -15349
rect 15656 -15381 15699 -15349
rect 15581 -15424 15699 -15381
rect 15741 -15349 15859 -15306
rect 15741 -15381 15784 -15349
rect 15784 -15381 15816 -15349
rect 15816 -15381 15859 -15349
rect 15741 -15424 15859 -15381
rect 15901 -15349 16019 -15306
rect 15901 -15381 15944 -15349
rect 15944 -15381 15976 -15349
rect 15976 -15381 16019 -15349
rect 15901 -15424 16019 -15381
rect 16061 -15349 16179 -15306
rect 16061 -15381 16104 -15349
rect 16104 -15381 16136 -15349
rect 16136 -15381 16179 -15349
rect 16061 -15424 16179 -15381
rect 16221 -15349 16339 -15306
rect 16221 -15381 16264 -15349
rect 16264 -15381 16296 -15349
rect 16296 -15381 16339 -15349
rect 16221 -15424 16339 -15381
rect 16381 -15349 16499 -15306
rect 16381 -15381 16424 -15349
rect 16424 -15381 16456 -15349
rect 16456 -15381 16499 -15349
rect 16381 -15424 16499 -15381
rect 16541 -15349 16659 -15306
rect 16541 -15381 16584 -15349
rect 16584 -15381 16616 -15349
rect 16616 -15381 16659 -15349
rect 16541 -15424 16659 -15381
rect 16701 -15349 16819 -15306
rect 16701 -15381 16744 -15349
rect 16744 -15381 16776 -15349
rect 16776 -15381 16819 -15349
rect 16701 -15424 16819 -15381
rect 16861 -15349 16979 -15306
rect 16861 -15381 16904 -15349
rect 16904 -15381 16936 -15349
rect 16936 -15381 16979 -15349
rect 16861 -15424 16979 -15381
rect 17021 -15349 17139 -15306
rect 17021 -15381 17064 -15349
rect 17064 -15381 17096 -15349
rect 17096 -15381 17139 -15349
rect 17021 -15424 17139 -15381
rect 17181 -15349 17299 -15306
rect 17181 -15381 17224 -15349
rect 17224 -15381 17256 -15349
rect 17256 -15381 17299 -15349
rect 17181 -15424 17299 -15381
rect 17341 -15349 17459 -15306
rect 17341 -15381 17384 -15349
rect 17384 -15381 17416 -15349
rect 17416 -15381 17459 -15349
rect 17341 -15424 17459 -15381
rect 17501 -15349 17619 -15306
rect 17501 -15381 17544 -15349
rect 17544 -15381 17576 -15349
rect 17576 -15381 17619 -15349
rect 17501 -15424 17619 -15381
rect 17661 -15349 17779 -15306
rect 17661 -15381 17704 -15349
rect 17704 -15381 17736 -15349
rect 17736 -15381 17779 -15349
rect 17661 -15424 17779 -15381
rect 17821 -15349 17939 -15306
rect 17821 -15381 17864 -15349
rect 17864 -15381 17896 -15349
rect 17896 -15381 17939 -15349
rect 17821 -15424 17939 -15381
rect 17981 -15349 18099 -15306
rect 17981 -15381 18024 -15349
rect 18024 -15381 18056 -15349
rect 18056 -15381 18099 -15349
rect 17981 -15424 18099 -15381
rect 18141 -15349 18259 -15306
rect 18141 -15381 18184 -15349
rect 18184 -15381 18216 -15349
rect 18216 -15381 18259 -15349
rect 18141 -15424 18259 -15381
rect 18301 -15349 18419 -15306
rect 18301 -15381 18344 -15349
rect 18344 -15381 18376 -15349
rect 18376 -15381 18419 -15349
rect 18301 -15424 18419 -15381
rect 18461 -15349 18579 -15306
rect 18461 -15381 18504 -15349
rect 18504 -15381 18536 -15349
rect 18536 -15381 18579 -15349
rect 18461 -15424 18579 -15381
rect 18621 -15349 18739 -15306
rect 18809 -15319 18927 -15276
rect 18621 -15381 18664 -15349
rect 18664 -15381 18696 -15349
rect 18696 -15381 18739 -15349
rect 18621 -15424 18739 -15381
rect 21261 -11621 21379 -11578
rect 21261 -11653 21304 -11621
rect 21304 -11653 21336 -11621
rect 21336 -11653 21379 -11621
rect 21076 -11724 21194 -11681
rect 21261 -11696 21379 -11653
rect 21421 -11621 21539 -11578
rect 21421 -11653 21464 -11621
rect 21464 -11653 21496 -11621
rect 21496 -11653 21539 -11621
rect 21421 -11696 21539 -11653
rect 21581 -11621 21699 -11578
rect 21581 -11653 21624 -11621
rect 21624 -11653 21656 -11621
rect 21656 -11653 21699 -11621
rect 21581 -11696 21699 -11653
rect 21741 -11621 21859 -11578
rect 21741 -11653 21784 -11621
rect 21784 -11653 21816 -11621
rect 21816 -11653 21859 -11621
rect 21741 -11696 21859 -11653
rect 21901 -11621 22019 -11578
rect 21901 -11653 21944 -11621
rect 21944 -11653 21976 -11621
rect 21976 -11653 22019 -11621
rect 21901 -11696 22019 -11653
rect 22061 -11621 22179 -11578
rect 22061 -11653 22104 -11621
rect 22104 -11653 22136 -11621
rect 22136 -11653 22179 -11621
rect 22061 -11696 22179 -11653
rect 22221 -11621 22339 -11578
rect 22221 -11653 22264 -11621
rect 22264 -11653 22296 -11621
rect 22296 -11653 22339 -11621
rect 22221 -11696 22339 -11653
rect 22381 -11621 22499 -11578
rect 22381 -11653 22424 -11621
rect 22424 -11653 22456 -11621
rect 22456 -11653 22499 -11621
rect 22381 -11696 22499 -11653
rect 22541 -11621 22659 -11578
rect 22541 -11653 22584 -11621
rect 22584 -11653 22616 -11621
rect 22616 -11653 22659 -11621
rect 22541 -11696 22659 -11653
rect 22701 -11621 22819 -11578
rect 22701 -11653 22744 -11621
rect 22744 -11653 22776 -11621
rect 22776 -11653 22819 -11621
rect 22701 -11696 22819 -11653
rect 22861 -11621 22979 -11578
rect 22861 -11653 22904 -11621
rect 22904 -11653 22936 -11621
rect 22936 -11653 22979 -11621
rect 22861 -11696 22979 -11653
rect 23021 -11621 23139 -11578
rect 23021 -11653 23064 -11621
rect 23064 -11653 23096 -11621
rect 23096 -11653 23139 -11621
rect 23021 -11696 23139 -11653
rect 23181 -11621 23299 -11578
rect 23181 -11653 23224 -11621
rect 23224 -11653 23256 -11621
rect 23256 -11653 23299 -11621
rect 23181 -11696 23299 -11653
rect 23341 -11621 23459 -11578
rect 23341 -11653 23384 -11621
rect 23384 -11653 23416 -11621
rect 23416 -11653 23459 -11621
rect 23341 -11696 23459 -11653
rect 23501 -11621 23619 -11578
rect 23501 -11653 23544 -11621
rect 23544 -11653 23576 -11621
rect 23576 -11653 23619 -11621
rect 23501 -11696 23619 -11653
rect 23661 -11621 23779 -11578
rect 23661 -11653 23704 -11621
rect 23704 -11653 23736 -11621
rect 23736 -11653 23779 -11621
rect 23661 -11696 23779 -11653
rect 23821 -11621 23939 -11578
rect 23821 -11653 23864 -11621
rect 23864 -11653 23896 -11621
rect 23896 -11653 23939 -11621
rect 23821 -11696 23939 -11653
rect 23981 -11621 24099 -11578
rect 23981 -11653 24024 -11621
rect 24024 -11653 24056 -11621
rect 24056 -11653 24099 -11621
rect 23981 -11696 24099 -11653
rect 24141 -11621 24259 -11578
rect 24141 -11653 24184 -11621
rect 24184 -11653 24216 -11621
rect 24216 -11653 24259 -11621
rect 24141 -11696 24259 -11653
rect 24301 -11621 24419 -11578
rect 24301 -11653 24344 -11621
rect 24344 -11653 24376 -11621
rect 24376 -11653 24419 -11621
rect 24301 -11696 24419 -11653
rect 24461 -11621 24579 -11578
rect 24461 -11653 24504 -11621
rect 24504 -11653 24536 -11621
rect 24536 -11653 24579 -11621
rect 24461 -11696 24579 -11653
rect 24621 -11621 24739 -11578
rect 24621 -11653 24664 -11621
rect 24664 -11653 24696 -11621
rect 24696 -11653 24739 -11621
rect 24621 -11696 24739 -11653
rect 21076 -11756 21119 -11724
rect 21119 -11756 21151 -11724
rect 21151 -11756 21194 -11724
rect 21076 -11799 21194 -11756
rect 24809 -11724 24927 -11681
rect 24809 -11756 24852 -11724
rect 24852 -11756 24884 -11724
rect 24884 -11756 24927 -11724
rect 21076 -11884 21194 -11841
rect 21076 -11916 21119 -11884
rect 21119 -11916 21151 -11884
rect 21151 -11916 21194 -11884
rect 21076 -11959 21194 -11916
rect 21076 -12044 21194 -12001
rect 21076 -12076 21119 -12044
rect 21119 -12076 21151 -12044
rect 21151 -12076 21194 -12044
rect 21076 -12119 21194 -12076
rect 21076 -12204 21194 -12161
rect 21076 -12236 21119 -12204
rect 21119 -12236 21151 -12204
rect 21151 -12236 21194 -12204
rect 21076 -12279 21194 -12236
rect 21076 -12364 21194 -12321
rect 21076 -12396 21119 -12364
rect 21119 -12396 21151 -12364
rect 21151 -12396 21194 -12364
rect 21076 -12439 21194 -12396
rect 21076 -12524 21194 -12481
rect 21076 -12556 21119 -12524
rect 21119 -12556 21151 -12524
rect 21151 -12556 21194 -12524
rect 21076 -12599 21194 -12556
rect 21076 -12684 21194 -12641
rect 21076 -12716 21119 -12684
rect 21119 -12716 21151 -12684
rect 21151 -12716 21194 -12684
rect 21076 -12759 21194 -12716
rect 21076 -12844 21194 -12801
rect 21076 -12876 21119 -12844
rect 21119 -12876 21151 -12844
rect 21151 -12876 21194 -12844
rect 21076 -12919 21194 -12876
rect 21076 -13004 21194 -12961
rect 21076 -13036 21119 -13004
rect 21119 -13036 21151 -13004
rect 21151 -13036 21194 -13004
rect 21076 -13079 21194 -13036
rect 21076 -13164 21194 -13121
rect 21076 -13196 21119 -13164
rect 21119 -13196 21151 -13164
rect 21151 -13196 21194 -13164
rect 21076 -13239 21194 -13196
rect 21076 -13324 21194 -13281
rect 21076 -13356 21119 -13324
rect 21119 -13356 21151 -13324
rect 21151 -13356 21194 -13324
rect 21076 -13399 21194 -13356
rect 21076 -13484 21194 -13441
rect 21076 -13516 21119 -13484
rect 21119 -13516 21151 -13484
rect 21151 -13516 21194 -13484
rect 21076 -13559 21194 -13516
rect 21076 -13644 21194 -13601
rect 21076 -13676 21119 -13644
rect 21119 -13676 21151 -13644
rect 21151 -13676 21194 -13644
rect 21076 -13719 21194 -13676
rect 21076 -13804 21194 -13761
rect 21076 -13836 21119 -13804
rect 21119 -13836 21151 -13804
rect 21151 -13836 21194 -13804
rect 21076 -13879 21194 -13836
rect 21076 -13964 21194 -13921
rect 21076 -13996 21119 -13964
rect 21119 -13996 21151 -13964
rect 21151 -13996 21194 -13964
rect 21076 -14039 21194 -13996
rect 21076 -14124 21194 -14081
rect 21076 -14156 21119 -14124
rect 21119 -14156 21151 -14124
rect 21151 -14156 21194 -14124
rect 21076 -14199 21194 -14156
rect 21076 -14284 21194 -14241
rect 21076 -14316 21119 -14284
rect 21119 -14316 21151 -14284
rect 21151 -14316 21194 -14284
rect 21076 -14359 21194 -14316
rect 21076 -14444 21194 -14401
rect 21076 -14476 21119 -14444
rect 21119 -14476 21151 -14444
rect 21151 -14476 21194 -14444
rect 21076 -14519 21194 -14476
rect 21076 -14604 21194 -14561
rect 21076 -14636 21119 -14604
rect 21119 -14636 21151 -14604
rect 21151 -14636 21194 -14604
rect 21076 -14679 21194 -14636
rect 21076 -14764 21194 -14721
rect 21076 -14796 21119 -14764
rect 21119 -14796 21151 -14764
rect 21151 -14796 21194 -14764
rect 21076 -14839 21194 -14796
rect 21076 -14924 21194 -14881
rect 21076 -14956 21119 -14924
rect 21119 -14956 21151 -14924
rect 21151 -14956 21194 -14924
rect 21076 -14999 21194 -14956
rect 21076 -15084 21194 -15041
rect 21076 -15116 21119 -15084
rect 21119 -15116 21151 -15084
rect 21151 -15116 21194 -15084
rect 21076 -15159 21194 -15116
rect 21076 -15244 21194 -15201
rect 24809 -11799 24927 -11756
rect 24809 -11884 24927 -11841
rect 24809 -11916 24852 -11884
rect 24852 -11916 24884 -11884
rect 24884 -11916 24927 -11884
rect 24809 -11959 24927 -11916
rect 24809 -12044 24927 -12001
rect 24809 -12076 24852 -12044
rect 24852 -12076 24884 -12044
rect 24884 -12076 24927 -12044
rect 24809 -12119 24927 -12076
rect 24809 -12204 24927 -12161
rect 24809 -12236 24852 -12204
rect 24852 -12236 24884 -12204
rect 24884 -12236 24927 -12204
rect 24809 -12279 24927 -12236
rect 24809 -12364 24927 -12321
rect 24809 -12396 24852 -12364
rect 24852 -12396 24884 -12364
rect 24884 -12396 24927 -12364
rect 24809 -12439 24927 -12396
rect 24809 -12524 24927 -12481
rect 24809 -12556 24852 -12524
rect 24852 -12556 24884 -12524
rect 24884 -12556 24927 -12524
rect 24809 -12599 24927 -12556
rect 24809 -12684 24927 -12641
rect 24809 -12716 24852 -12684
rect 24852 -12716 24884 -12684
rect 24884 -12716 24927 -12684
rect 24809 -12759 24927 -12716
rect 24809 -12844 24927 -12801
rect 24809 -12876 24852 -12844
rect 24852 -12876 24884 -12844
rect 24884 -12876 24927 -12844
rect 24809 -12919 24927 -12876
rect 24809 -13004 24927 -12961
rect 24809 -13036 24852 -13004
rect 24852 -13036 24884 -13004
rect 24884 -13036 24927 -13004
rect 24809 -13079 24927 -13036
rect 24809 -13164 24927 -13121
rect 24809 -13196 24852 -13164
rect 24852 -13196 24884 -13164
rect 24884 -13196 24927 -13164
rect 24809 -13239 24927 -13196
rect 24809 -13324 24927 -13281
rect 24809 -13356 24852 -13324
rect 24852 -13356 24884 -13324
rect 24884 -13356 24927 -13324
rect 24809 -13399 24927 -13356
rect 24809 -13484 24927 -13441
rect 24809 -13516 24852 -13484
rect 24852 -13516 24884 -13484
rect 24884 -13516 24927 -13484
rect 24809 -13559 24927 -13516
rect 24809 -13644 24927 -13601
rect 24809 -13676 24852 -13644
rect 24852 -13676 24884 -13644
rect 24884 -13676 24927 -13644
rect 24809 -13719 24927 -13676
rect 24809 -13804 24927 -13761
rect 24809 -13836 24852 -13804
rect 24852 -13836 24884 -13804
rect 24884 -13836 24927 -13804
rect 24809 -13879 24927 -13836
rect 24809 -13964 24927 -13921
rect 24809 -13996 24852 -13964
rect 24852 -13996 24884 -13964
rect 24884 -13996 24927 -13964
rect 24809 -14039 24927 -13996
rect 24809 -14124 24927 -14081
rect 24809 -14156 24852 -14124
rect 24852 -14156 24884 -14124
rect 24884 -14156 24927 -14124
rect 24809 -14199 24927 -14156
rect 24809 -14284 24927 -14241
rect 24809 -14316 24852 -14284
rect 24852 -14316 24884 -14284
rect 24884 -14316 24927 -14284
rect 24809 -14359 24927 -14316
rect 24809 -14444 24927 -14401
rect 24809 -14476 24852 -14444
rect 24852 -14476 24884 -14444
rect 24884 -14476 24927 -14444
rect 24809 -14519 24927 -14476
rect 24809 -14604 24927 -14561
rect 24809 -14636 24852 -14604
rect 24852 -14636 24884 -14604
rect 24884 -14636 24927 -14604
rect 24809 -14679 24927 -14636
rect 24809 -14764 24927 -14721
rect 24809 -14796 24852 -14764
rect 24852 -14796 24884 -14764
rect 24884 -14796 24927 -14764
rect 24809 -14839 24927 -14796
rect 24809 -14924 24927 -14881
rect 24809 -14956 24852 -14924
rect 24852 -14956 24884 -14924
rect 24884 -14956 24927 -14924
rect 24809 -14999 24927 -14956
rect 24809 -15084 24927 -15041
rect 24809 -15116 24852 -15084
rect 24852 -15116 24884 -15084
rect 24884 -15116 24927 -15084
rect 24809 -15159 24927 -15116
rect 21076 -15276 21119 -15244
rect 21119 -15276 21151 -15244
rect 21151 -15276 21194 -15244
rect 21076 -15319 21194 -15276
rect 24809 -15244 24927 -15201
rect 24809 -15276 24852 -15244
rect 24852 -15276 24884 -15244
rect 24884 -15276 24927 -15244
rect 21261 -15349 21379 -15306
rect 21261 -15381 21304 -15349
rect 21304 -15381 21336 -15349
rect 21336 -15381 21379 -15349
rect 21261 -15424 21379 -15381
rect 21421 -15349 21539 -15306
rect 21421 -15381 21464 -15349
rect 21464 -15381 21496 -15349
rect 21496 -15381 21539 -15349
rect 21421 -15424 21539 -15381
rect 21581 -15349 21699 -15306
rect 21581 -15381 21624 -15349
rect 21624 -15381 21656 -15349
rect 21656 -15381 21699 -15349
rect 21581 -15424 21699 -15381
rect 21741 -15349 21859 -15306
rect 21741 -15381 21784 -15349
rect 21784 -15381 21816 -15349
rect 21816 -15381 21859 -15349
rect 21741 -15424 21859 -15381
rect 21901 -15349 22019 -15306
rect 21901 -15381 21944 -15349
rect 21944 -15381 21976 -15349
rect 21976 -15381 22019 -15349
rect 21901 -15424 22019 -15381
rect 22061 -15349 22179 -15306
rect 22061 -15381 22104 -15349
rect 22104 -15381 22136 -15349
rect 22136 -15381 22179 -15349
rect 22061 -15424 22179 -15381
rect 22221 -15349 22339 -15306
rect 22221 -15381 22264 -15349
rect 22264 -15381 22296 -15349
rect 22296 -15381 22339 -15349
rect 22221 -15424 22339 -15381
rect 22381 -15349 22499 -15306
rect 22381 -15381 22424 -15349
rect 22424 -15381 22456 -15349
rect 22456 -15381 22499 -15349
rect 22381 -15424 22499 -15381
rect 22541 -15349 22659 -15306
rect 22541 -15381 22584 -15349
rect 22584 -15381 22616 -15349
rect 22616 -15381 22659 -15349
rect 22541 -15424 22659 -15381
rect 22701 -15349 22819 -15306
rect 22701 -15381 22744 -15349
rect 22744 -15381 22776 -15349
rect 22776 -15381 22819 -15349
rect 22701 -15424 22819 -15381
rect 22861 -15349 22979 -15306
rect 22861 -15381 22904 -15349
rect 22904 -15381 22936 -15349
rect 22936 -15381 22979 -15349
rect 22861 -15424 22979 -15381
rect 23021 -15349 23139 -15306
rect 23021 -15381 23064 -15349
rect 23064 -15381 23096 -15349
rect 23096 -15381 23139 -15349
rect 23021 -15424 23139 -15381
rect 23181 -15349 23299 -15306
rect 23181 -15381 23224 -15349
rect 23224 -15381 23256 -15349
rect 23256 -15381 23299 -15349
rect 23181 -15424 23299 -15381
rect 23341 -15349 23459 -15306
rect 23341 -15381 23384 -15349
rect 23384 -15381 23416 -15349
rect 23416 -15381 23459 -15349
rect 23341 -15424 23459 -15381
rect 23501 -15349 23619 -15306
rect 23501 -15381 23544 -15349
rect 23544 -15381 23576 -15349
rect 23576 -15381 23619 -15349
rect 23501 -15424 23619 -15381
rect 23661 -15349 23779 -15306
rect 23661 -15381 23704 -15349
rect 23704 -15381 23736 -15349
rect 23736 -15381 23779 -15349
rect 23661 -15424 23779 -15381
rect 23821 -15349 23939 -15306
rect 23821 -15381 23864 -15349
rect 23864 -15381 23896 -15349
rect 23896 -15381 23939 -15349
rect 23821 -15424 23939 -15381
rect 23981 -15349 24099 -15306
rect 23981 -15381 24024 -15349
rect 24024 -15381 24056 -15349
rect 24056 -15381 24099 -15349
rect 23981 -15424 24099 -15381
rect 24141 -15349 24259 -15306
rect 24141 -15381 24184 -15349
rect 24184 -15381 24216 -15349
rect 24216 -15381 24259 -15349
rect 24141 -15424 24259 -15381
rect 24301 -15349 24419 -15306
rect 24301 -15381 24344 -15349
rect 24344 -15381 24376 -15349
rect 24376 -15381 24419 -15349
rect 24301 -15424 24419 -15381
rect 24461 -15349 24579 -15306
rect 24461 -15381 24504 -15349
rect 24504 -15381 24536 -15349
rect 24536 -15381 24579 -15349
rect 24461 -15424 24579 -15381
rect 24621 -15349 24739 -15306
rect 24809 -15319 24927 -15276
rect 24621 -15381 24664 -15349
rect 24664 -15381 24696 -15349
rect 24696 -15381 24739 -15349
rect 24621 -15424 24739 -15381
<< metal5 >>
rect 3000 9424 7000 9500
rect 3000 9319 3261 9424
rect 3000 9201 3073 9319
rect 3191 9306 3261 9319
rect 3379 9306 3421 9424
rect 3539 9306 3581 9424
rect 3699 9306 3741 9424
rect 3859 9306 3901 9424
rect 4019 9306 4061 9424
rect 4179 9306 4221 9424
rect 4339 9306 4381 9424
rect 4499 9306 4541 9424
rect 4659 9306 4701 9424
rect 4819 9306 4861 9424
rect 4979 9306 5021 9424
rect 5139 9306 5181 9424
rect 5299 9306 5341 9424
rect 5459 9306 5501 9424
rect 5619 9306 5661 9424
rect 5779 9306 5821 9424
rect 5939 9306 5981 9424
rect 6099 9306 6141 9424
rect 6259 9306 6301 9424
rect 6419 9306 6461 9424
rect 6579 9306 6621 9424
rect 6739 9319 7000 9424
rect 6739 9306 6806 9319
rect 3191 9201 6806 9306
rect 6924 9201 7000 9319
rect 3000 9159 7000 9201
rect 3000 9041 3073 9159
rect 3191 9041 6806 9159
rect 6924 9041 7000 9159
rect 3000 8999 7000 9041
rect 3000 8881 3073 8999
rect 3191 8881 6806 8999
rect 6924 8881 7000 8999
rect 3000 8839 7000 8881
rect 3000 8721 3073 8839
rect 3191 8721 6806 8839
rect 6924 8721 7000 8839
rect 3000 8679 7000 8721
rect 3000 8561 3073 8679
rect 3191 8561 6806 8679
rect 6924 8561 7000 8679
rect 3000 8519 7000 8561
rect 3000 8401 3073 8519
rect 3191 8401 6806 8519
rect 6924 8401 7000 8519
rect 3000 8359 7000 8401
rect 3000 8241 3073 8359
rect 3191 8241 6806 8359
rect 6924 8241 7000 8359
rect 3000 8199 7000 8241
rect 3000 8081 3073 8199
rect 3191 8081 6806 8199
rect 6924 8081 7000 8199
rect 3000 8039 7000 8081
rect 3000 7921 3073 8039
rect 3191 7921 6806 8039
rect 6924 7921 7000 8039
rect 3000 7879 7000 7921
rect 3000 7761 3073 7879
rect 3191 7761 6806 7879
rect 6924 7761 7000 7879
rect 3000 7719 7000 7761
rect 3000 7601 3073 7719
rect 3191 7601 6806 7719
rect 6924 7601 7000 7719
rect 3000 7559 7000 7601
rect 3000 7441 3073 7559
rect 3191 7441 6806 7559
rect 6924 7441 7000 7559
rect 3000 7399 7000 7441
rect 3000 7281 3073 7399
rect 3191 7281 6806 7399
rect 6924 7281 7000 7399
rect 3000 7239 7000 7281
rect 3000 7121 3073 7239
rect 3191 7121 6806 7239
rect 6924 7121 7000 7239
rect 3000 7079 7000 7121
rect 3000 6961 3073 7079
rect 3191 6961 6806 7079
rect 6924 6961 7000 7079
rect 3000 6919 7000 6961
rect 3000 6801 3073 6919
rect 3191 6801 6806 6919
rect 6924 6801 7000 6919
rect 3000 6759 7000 6801
rect 3000 6641 3073 6759
rect 3191 6641 6806 6759
rect 6924 6641 7000 6759
rect 3000 6599 7000 6641
rect 3000 6481 3073 6599
rect 3191 6481 6806 6599
rect 6924 6481 7000 6599
rect 3000 6439 7000 6481
rect 3000 6321 3073 6439
rect 3191 6321 6806 6439
rect 6924 6321 7000 6439
rect 3000 6279 7000 6321
rect 3000 6161 3073 6279
rect 3191 6161 6806 6279
rect 6924 6161 7000 6279
rect 3000 6119 7000 6161
rect 3000 6001 3073 6119
rect 3191 6001 6806 6119
rect 6924 6001 7000 6119
rect 3000 5959 7000 6001
rect 3000 5841 3073 5959
rect 3191 5841 6806 5959
rect 6924 5841 7000 5959
rect 3000 5799 7000 5841
rect 3000 5681 3073 5799
rect 3191 5696 6806 5799
rect 3191 5681 3261 5696
rect 3000 5578 3261 5681
rect 3379 5578 3421 5696
rect 3539 5578 3581 5696
rect 3699 5578 3741 5696
rect 3859 5578 3901 5696
rect 4019 5578 4061 5696
rect 4179 5578 4221 5696
rect 4339 5578 4381 5696
rect 4499 5578 4541 5696
rect 4659 5578 4701 5696
rect 4819 5578 4861 5696
rect 4979 5578 5021 5696
rect 5139 5578 5181 5696
rect 5299 5578 5341 5696
rect 5459 5578 5501 5696
rect 5619 5578 5661 5696
rect 5779 5578 5821 5696
rect 5939 5578 5981 5696
rect 6099 5578 6141 5696
rect 6259 5578 6301 5696
rect 6419 5578 6461 5696
rect 6579 5578 6621 5696
rect 6739 5681 6806 5696
rect 6924 5681 7000 5799
rect 6739 5578 7000 5681
rect 3000 5500 7000 5578
rect 9000 9424 13000 9500
rect 9000 9319 9261 9424
rect 9000 9201 9073 9319
rect 9191 9306 9261 9319
rect 9379 9306 9421 9424
rect 9539 9306 9581 9424
rect 9699 9306 9741 9424
rect 9859 9306 9901 9424
rect 10019 9306 10061 9424
rect 10179 9306 10221 9424
rect 10339 9306 10381 9424
rect 10499 9306 10541 9424
rect 10659 9306 10701 9424
rect 10819 9306 10861 9424
rect 10979 9306 11021 9424
rect 11139 9306 11181 9424
rect 11299 9306 11341 9424
rect 11459 9306 11501 9424
rect 11619 9306 11661 9424
rect 11779 9306 11821 9424
rect 11939 9306 11981 9424
rect 12099 9306 12141 9424
rect 12259 9306 12301 9424
rect 12419 9306 12461 9424
rect 12579 9306 12621 9424
rect 12739 9319 13000 9424
rect 12739 9306 12806 9319
rect 9191 9201 12806 9306
rect 12924 9201 13000 9319
rect 9000 9159 13000 9201
rect 9000 9041 9073 9159
rect 9191 9041 12806 9159
rect 12924 9041 13000 9159
rect 9000 8999 13000 9041
rect 9000 8881 9073 8999
rect 9191 8881 12806 8999
rect 12924 8881 13000 8999
rect 9000 8839 13000 8881
rect 9000 8721 9073 8839
rect 9191 8721 12806 8839
rect 12924 8721 13000 8839
rect 9000 8679 13000 8721
rect 9000 8561 9073 8679
rect 9191 8561 12806 8679
rect 12924 8561 13000 8679
rect 9000 8519 13000 8561
rect 9000 8401 9073 8519
rect 9191 8401 12806 8519
rect 12924 8401 13000 8519
rect 9000 8359 13000 8401
rect 9000 8241 9073 8359
rect 9191 8241 12806 8359
rect 12924 8241 13000 8359
rect 9000 8199 13000 8241
rect 9000 8081 9073 8199
rect 9191 8081 12806 8199
rect 12924 8081 13000 8199
rect 9000 8039 13000 8081
rect 9000 7921 9073 8039
rect 9191 7921 12806 8039
rect 12924 7921 13000 8039
rect 9000 7879 13000 7921
rect 9000 7761 9073 7879
rect 9191 7761 12806 7879
rect 12924 7761 13000 7879
rect 9000 7719 13000 7761
rect 9000 7601 9073 7719
rect 9191 7601 12806 7719
rect 12924 7601 13000 7719
rect 9000 7559 13000 7601
rect 9000 7441 9073 7559
rect 9191 7441 12806 7559
rect 12924 7441 13000 7559
rect 9000 7399 13000 7441
rect 9000 7281 9073 7399
rect 9191 7281 12806 7399
rect 12924 7281 13000 7399
rect 9000 7239 13000 7281
rect 9000 7121 9073 7239
rect 9191 7121 12806 7239
rect 12924 7121 13000 7239
rect 9000 7079 13000 7121
rect 9000 6961 9073 7079
rect 9191 6961 12806 7079
rect 12924 6961 13000 7079
rect 9000 6919 13000 6961
rect 9000 6801 9073 6919
rect 9191 6801 12806 6919
rect 12924 6801 13000 6919
rect 9000 6759 13000 6801
rect 9000 6641 9073 6759
rect 9191 6641 12806 6759
rect 12924 6641 13000 6759
rect 9000 6599 13000 6641
rect 9000 6481 9073 6599
rect 9191 6481 12806 6599
rect 12924 6481 13000 6599
rect 9000 6439 13000 6481
rect 9000 6321 9073 6439
rect 9191 6321 12806 6439
rect 12924 6321 13000 6439
rect 9000 6279 13000 6321
rect 9000 6161 9073 6279
rect 9191 6161 12806 6279
rect 12924 6161 13000 6279
rect 9000 6119 13000 6161
rect 9000 6001 9073 6119
rect 9191 6001 12806 6119
rect 12924 6001 13000 6119
rect 9000 5959 13000 6001
rect 9000 5841 9073 5959
rect 9191 5841 12806 5959
rect 12924 5841 13000 5959
rect 9000 5799 13000 5841
rect 9000 5681 9073 5799
rect 9191 5696 12806 5799
rect 9191 5681 9261 5696
rect 9000 5578 9261 5681
rect 9379 5578 9421 5696
rect 9539 5578 9581 5696
rect 9699 5578 9741 5696
rect 9859 5578 9901 5696
rect 10019 5578 10061 5696
rect 10179 5578 10221 5696
rect 10339 5578 10381 5696
rect 10499 5578 10541 5696
rect 10659 5578 10701 5696
rect 10819 5578 10861 5696
rect 10979 5578 11021 5696
rect 11139 5578 11181 5696
rect 11299 5578 11341 5696
rect 11459 5578 11501 5696
rect 11619 5578 11661 5696
rect 11779 5578 11821 5696
rect 11939 5578 11981 5696
rect 12099 5578 12141 5696
rect 12259 5578 12301 5696
rect 12419 5578 12461 5696
rect 12579 5578 12621 5696
rect 12739 5681 12806 5696
rect 12924 5681 13000 5799
rect 12739 5578 13000 5681
rect 9000 5500 13000 5578
rect 15000 9424 19000 9500
rect 15000 9319 15261 9424
rect 15000 9201 15073 9319
rect 15191 9306 15261 9319
rect 15379 9306 15421 9424
rect 15539 9306 15581 9424
rect 15699 9306 15741 9424
rect 15859 9306 15901 9424
rect 16019 9306 16061 9424
rect 16179 9306 16221 9424
rect 16339 9306 16381 9424
rect 16499 9306 16541 9424
rect 16659 9306 16701 9424
rect 16819 9306 16861 9424
rect 16979 9306 17021 9424
rect 17139 9306 17181 9424
rect 17299 9306 17341 9424
rect 17459 9306 17501 9424
rect 17619 9306 17661 9424
rect 17779 9306 17821 9424
rect 17939 9306 17981 9424
rect 18099 9306 18141 9424
rect 18259 9306 18301 9424
rect 18419 9306 18461 9424
rect 18579 9306 18621 9424
rect 18739 9319 19000 9424
rect 18739 9306 18806 9319
rect 15191 9201 18806 9306
rect 18924 9201 19000 9319
rect 15000 9159 19000 9201
rect 15000 9041 15073 9159
rect 15191 9041 18806 9159
rect 18924 9041 19000 9159
rect 15000 8999 19000 9041
rect 15000 8881 15073 8999
rect 15191 8881 18806 8999
rect 18924 8881 19000 8999
rect 15000 8839 19000 8881
rect 15000 8721 15073 8839
rect 15191 8721 18806 8839
rect 18924 8721 19000 8839
rect 15000 8679 19000 8721
rect 15000 8561 15073 8679
rect 15191 8561 18806 8679
rect 18924 8561 19000 8679
rect 15000 8519 19000 8561
rect 15000 8401 15073 8519
rect 15191 8401 18806 8519
rect 18924 8401 19000 8519
rect 15000 8359 19000 8401
rect 15000 8241 15073 8359
rect 15191 8241 18806 8359
rect 18924 8241 19000 8359
rect 15000 8199 19000 8241
rect 15000 8081 15073 8199
rect 15191 8081 18806 8199
rect 18924 8081 19000 8199
rect 15000 8039 19000 8081
rect 15000 7921 15073 8039
rect 15191 7921 18806 8039
rect 18924 7921 19000 8039
rect 15000 7879 19000 7921
rect 15000 7761 15073 7879
rect 15191 7761 18806 7879
rect 18924 7761 19000 7879
rect 15000 7719 19000 7761
rect 15000 7601 15073 7719
rect 15191 7601 18806 7719
rect 18924 7601 19000 7719
rect 15000 7559 19000 7601
rect 15000 7441 15073 7559
rect 15191 7441 18806 7559
rect 18924 7441 19000 7559
rect 15000 7399 19000 7441
rect 15000 7281 15073 7399
rect 15191 7281 18806 7399
rect 18924 7281 19000 7399
rect 15000 7239 19000 7281
rect 15000 7121 15073 7239
rect 15191 7121 18806 7239
rect 18924 7121 19000 7239
rect 15000 7079 19000 7121
rect 15000 6961 15073 7079
rect 15191 6961 18806 7079
rect 18924 6961 19000 7079
rect 15000 6919 19000 6961
rect 15000 6801 15073 6919
rect 15191 6801 18806 6919
rect 18924 6801 19000 6919
rect 15000 6759 19000 6801
rect 15000 6641 15073 6759
rect 15191 6641 18806 6759
rect 18924 6641 19000 6759
rect 15000 6599 19000 6641
rect 15000 6481 15073 6599
rect 15191 6481 18806 6599
rect 18924 6481 19000 6599
rect 15000 6439 19000 6481
rect 15000 6321 15073 6439
rect 15191 6321 18806 6439
rect 18924 6321 19000 6439
rect 15000 6279 19000 6321
rect 15000 6161 15073 6279
rect 15191 6161 18806 6279
rect 18924 6161 19000 6279
rect 15000 6119 19000 6161
rect 15000 6001 15073 6119
rect 15191 6001 18806 6119
rect 18924 6001 19000 6119
rect 15000 5959 19000 6001
rect 15000 5841 15073 5959
rect 15191 5841 18806 5959
rect 18924 5841 19000 5959
rect 15000 5799 19000 5841
rect 15000 5681 15073 5799
rect 15191 5696 18806 5799
rect 15191 5681 15261 5696
rect 15000 5578 15261 5681
rect 15379 5578 15421 5696
rect 15539 5578 15581 5696
rect 15699 5578 15741 5696
rect 15859 5578 15901 5696
rect 16019 5578 16061 5696
rect 16179 5578 16221 5696
rect 16339 5578 16381 5696
rect 16499 5578 16541 5696
rect 16659 5578 16701 5696
rect 16819 5578 16861 5696
rect 16979 5578 17021 5696
rect 17139 5578 17181 5696
rect 17299 5578 17341 5696
rect 17459 5578 17501 5696
rect 17619 5578 17661 5696
rect 17779 5578 17821 5696
rect 17939 5578 17981 5696
rect 18099 5578 18141 5696
rect 18259 5578 18301 5696
rect 18419 5578 18461 5696
rect 18579 5578 18621 5696
rect 18739 5681 18806 5696
rect 18924 5681 19000 5799
rect 18739 5578 19000 5681
rect 15000 5500 19000 5578
rect 21000 9424 25000 9500
rect 21000 9319 21261 9424
rect 21000 9201 21073 9319
rect 21191 9306 21261 9319
rect 21379 9306 21421 9424
rect 21539 9306 21581 9424
rect 21699 9306 21741 9424
rect 21859 9306 21901 9424
rect 22019 9306 22061 9424
rect 22179 9306 22221 9424
rect 22339 9306 22381 9424
rect 22499 9306 22541 9424
rect 22659 9306 22701 9424
rect 22819 9306 22861 9424
rect 22979 9306 23021 9424
rect 23139 9306 23181 9424
rect 23299 9306 23341 9424
rect 23459 9306 23501 9424
rect 23619 9306 23661 9424
rect 23779 9306 23821 9424
rect 23939 9306 23981 9424
rect 24099 9306 24141 9424
rect 24259 9306 24301 9424
rect 24419 9306 24461 9424
rect 24579 9306 24621 9424
rect 24739 9319 25000 9424
rect 24739 9306 24806 9319
rect 21191 9201 24806 9306
rect 24924 9201 25000 9319
rect 21000 9159 25000 9201
rect 21000 9041 21073 9159
rect 21191 9041 24806 9159
rect 24924 9041 25000 9159
rect 21000 8999 25000 9041
rect 21000 8881 21073 8999
rect 21191 8881 24806 8999
rect 24924 8881 25000 8999
rect 21000 8839 25000 8881
rect 21000 8721 21073 8839
rect 21191 8721 24806 8839
rect 24924 8721 25000 8839
rect 21000 8679 25000 8721
rect 21000 8561 21073 8679
rect 21191 8561 24806 8679
rect 24924 8561 25000 8679
rect 21000 8519 25000 8561
rect 21000 8401 21073 8519
rect 21191 8401 24806 8519
rect 24924 8401 25000 8519
rect 21000 8359 25000 8401
rect 21000 8241 21073 8359
rect 21191 8241 24806 8359
rect 24924 8241 25000 8359
rect 21000 8199 25000 8241
rect 21000 8081 21073 8199
rect 21191 8081 24806 8199
rect 24924 8081 25000 8199
rect 21000 8039 25000 8081
rect 21000 7921 21073 8039
rect 21191 7921 24806 8039
rect 24924 7921 25000 8039
rect 21000 7879 25000 7921
rect 21000 7761 21073 7879
rect 21191 7761 24806 7879
rect 24924 7761 25000 7879
rect 21000 7719 25000 7761
rect 21000 7601 21073 7719
rect 21191 7601 24806 7719
rect 24924 7601 25000 7719
rect 21000 7559 25000 7601
rect 21000 7441 21073 7559
rect 21191 7441 24806 7559
rect 24924 7441 25000 7559
rect 21000 7399 25000 7441
rect 21000 7281 21073 7399
rect 21191 7281 24806 7399
rect 24924 7281 25000 7399
rect 21000 7239 25000 7281
rect 21000 7121 21073 7239
rect 21191 7121 24806 7239
rect 24924 7121 25000 7239
rect 21000 7079 25000 7121
rect 21000 6961 21073 7079
rect 21191 6961 24806 7079
rect 24924 6961 25000 7079
rect 21000 6919 25000 6961
rect 21000 6801 21073 6919
rect 21191 6801 24806 6919
rect 24924 6801 25000 6919
rect 21000 6759 25000 6801
rect 21000 6641 21073 6759
rect 21191 6641 24806 6759
rect 24924 6641 25000 6759
rect 21000 6599 25000 6641
rect 21000 6481 21073 6599
rect 21191 6481 24806 6599
rect 24924 6481 25000 6599
rect 21000 6439 25000 6481
rect 21000 6321 21073 6439
rect 21191 6321 24806 6439
rect 24924 6321 25000 6439
rect 21000 6279 25000 6321
rect 21000 6161 21073 6279
rect 21191 6161 24806 6279
rect 24924 6161 25000 6279
rect 21000 6119 25000 6161
rect 21000 6001 21073 6119
rect 21191 6001 24806 6119
rect 24924 6001 25000 6119
rect 21000 5959 25000 6001
rect 21000 5841 21073 5959
rect 21191 5841 24806 5959
rect 24924 5841 25000 5959
rect 21000 5799 25000 5841
rect 21000 5681 21073 5799
rect 21191 5696 24806 5799
rect 21191 5681 21261 5696
rect 21000 5578 21261 5681
rect 21379 5578 21421 5696
rect 21539 5578 21581 5696
rect 21699 5578 21741 5696
rect 21859 5578 21901 5696
rect 22019 5578 22061 5696
rect 22179 5578 22221 5696
rect 22339 5578 22381 5696
rect 22499 5578 22541 5696
rect 22659 5578 22701 5696
rect 22819 5578 22861 5696
rect 22979 5578 23021 5696
rect 23139 5578 23181 5696
rect 23299 5578 23341 5696
rect 23459 5578 23501 5696
rect 23619 5578 23661 5696
rect 23779 5578 23821 5696
rect 23939 5578 23981 5696
rect 24099 5578 24141 5696
rect 24259 5578 24301 5696
rect 24419 5578 24461 5696
rect 24579 5578 24621 5696
rect 24739 5681 24806 5696
rect 24924 5681 25000 5799
rect 24739 5578 25000 5681
rect 21000 5500 25000 5578
rect 3000 3424 7000 3500
rect 3000 3319 3261 3424
rect 3000 3201 3073 3319
rect 3191 3306 3261 3319
rect 3379 3306 3421 3424
rect 3539 3306 3581 3424
rect 3699 3306 3741 3424
rect 3859 3306 3901 3424
rect 4019 3306 4061 3424
rect 4179 3306 4221 3424
rect 4339 3306 4381 3424
rect 4499 3306 4541 3424
rect 4659 3306 4701 3424
rect 4819 3306 4861 3424
rect 4979 3306 5021 3424
rect 5139 3306 5181 3424
rect 5299 3306 5341 3424
rect 5459 3306 5501 3424
rect 5619 3306 5661 3424
rect 5779 3306 5821 3424
rect 5939 3306 5981 3424
rect 6099 3306 6141 3424
rect 6259 3306 6301 3424
rect 6419 3306 6461 3424
rect 6579 3306 6621 3424
rect 6739 3319 7000 3424
rect 6739 3306 6806 3319
rect 3191 3201 6806 3306
rect 6924 3201 7000 3319
rect 3000 3159 7000 3201
rect 3000 3041 3073 3159
rect 3191 3041 6806 3159
rect 6924 3041 7000 3159
rect 3000 2999 7000 3041
rect 3000 2881 3073 2999
rect 3191 2881 6806 2999
rect 6924 2881 7000 2999
rect 3000 2839 7000 2881
rect 3000 2721 3073 2839
rect 3191 2721 6806 2839
rect 6924 2721 7000 2839
rect 3000 2679 7000 2721
rect 3000 2561 3073 2679
rect 3191 2561 6806 2679
rect 6924 2561 7000 2679
rect 3000 2519 7000 2561
rect 3000 2401 3073 2519
rect 3191 2401 6806 2519
rect 6924 2401 7000 2519
rect 3000 2359 7000 2401
rect 3000 2241 3073 2359
rect 3191 2241 6806 2359
rect 6924 2241 7000 2359
rect 3000 2199 7000 2241
rect 3000 2081 3073 2199
rect 3191 2081 6806 2199
rect 6924 2081 7000 2199
rect 3000 2039 7000 2081
rect 3000 1921 3073 2039
rect 3191 1921 6806 2039
rect 6924 1921 7000 2039
rect 3000 1879 7000 1921
rect 3000 1761 3073 1879
rect 3191 1761 6806 1879
rect 6924 1761 7000 1879
rect 3000 1719 7000 1761
rect 3000 1601 3073 1719
rect 3191 1601 6806 1719
rect 6924 1601 7000 1719
rect 3000 1559 7000 1601
rect 3000 1441 3073 1559
rect 3191 1441 6806 1559
rect 6924 1441 7000 1559
rect 3000 1399 7000 1441
rect 3000 1281 3073 1399
rect 3191 1281 6806 1399
rect 6924 1281 7000 1399
rect 3000 1239 7000 1281
rect 3000 1121 3073 1239
rect 3191 1121 6806 1239
rect 6924 1121 7000 1239
rect 3000 1079 7000 1121
rect 3000 961 3073 1079
rect 3191 961 6806 1079
rect 6924 961 7000 1079
rect 3000 919 7000 961
rect 3000 801 3073 919
rect 3191 801 6806 919
rect 6924 801 7000 919
rect 3000 759 7000 801
rect 3000 641 3073 759
rect 3191 641 6806 759
rect 6924 641 7000 759
rect 3000 599 7000 641
rect 3000 481 3073 599
rect 3191 481 6806 599
rect 6924 481 7000 599
rect 3000 439 7000 481
rect 3000 321 3073 439
rect 3191 321 6806 439
rect 6924 321 7000 439
rect 3000 279 7000 321
rect 3000 161 3073 279
rect 3191 161 6806 279
rect 6924 161 7000 279
rect 3000 119 7000 161
rect 3000 1 3073 119
rect 3191 1 6806 119
rect 6924 1 7000 119
rect 3000 -41 7000 1
rect 3000 -159 3073 -41
rect 3191 -159 6806 -41
rect 6924 -159 7000 -41
rect 3000 -201 7000 -159
rect 3000 -319 3073 -201
rect 3191 -304 6806 -201
rect 3191 -319 3261 -304
rect 3000 -422 3261 -319
rect 3379 -422 3421 -304
rect 3539 -422 3581 -304
rect 3699 -422 3741 -304
rect 3859 -422 3901 -304
rect 4019 -422 4061 -304
rect 4179 -422 4221 -304
rect 4339 -422 4381 -304
rect 4499 -422 4541 -304
rect 4659 -422 4701 -304
rect 4819 -422 4861 -304
rect 4979 -422 5021 -304
rect 5139 -422 5181 -304
rect 5299 -422 5341 -304
rect 5459 -422 5501 -304
rect 5619 -422 5661 -304
rect 5779 -422 5821 -304
rect 5939 -422 5981 -304
rect 6099 -422 6141 -304
rect 6259 -422 6301 -304
rect 6419 -422 6461 -304
rect 6579 -422 6621 -304
rect 6739 -319 6806 -304
rect 6924 -319 7000 -201
rect 6739 -422 7000 -319
rect 3000 -500 7000 -422
rect 9000 3424 13000 3500
rect 9000 3319 9261 3424
rect 9000 3201 9073 3319
rect 9191 3306 9261 3319
rect 9379 3306 9421 3424
rect 9539 3306 9581 3424
rect 9699 3306 9741 3424
rect 9859 3306 9901 3424
rect 10019 3306 10061 3424
rect 10179 3306 10221 3424
rect 10339 3306 10381 3424
rect 10499 3306 10541 3424
rect 10659 3306 10701 3424
rect 10819 3306 10861 3424
rect 10979 3306 11021 3424
rect 11139 3306 11181 3424
rect 11299 3306 11341 3424
rect 11459 3306 11501 3424
rect 11619 3306 11661 3424
rect 11779 3306 11821 3424
rect 11939 3306 11981 3424
rect 12099 3306 12141 3424
rect 12259 3306 12301 3424
rect 12419 3306 12461 3424
rect 12579 3306 12621 3424
rect 12739 3319 13000 3424
rect 12739 3306 12806 3319
rect 9191 3201 12806 3306
rect 12924 3201 13000 3319
rect 9000 3159 13000 3201
rect 9000 3041 9073 3159
rect 9191 3041 12806 3159
rect 12924 3041 13000 3159
rect 9000 2999 13000 3041
rect 9000 2881 9073 2999
rect 9191 2881 12806 2999
rect 12924 2881 13000 2999
rect 9000 2839 13000 2881
rect 9000 2721 9073 2839
rect 9191 2721 12806 2839
rect 12924 2721 13000 2839
rect 9000 2679 13000 2721
rect 9000 2561 9073 2679
rect 9191 2561 12806 2679
rect 12924 2561 13000 2679
rect 9000 2519 13000 2561
rect 9000 2401 9073 2519
rect 9191 2401 12806 2519
rect 12924 2401 13000 2519
rect 9000 2359 13000 2401
rect 9000 2241 9073 2359
rect 9191 2241 12806 2359
rect 12924 2241 13000 2359
rect 9000 2199 13000 2241
rect 9000 2081 9073 2199
rect 9191 2081 12806 2199
rect 12924 2081 13000 2199
rect 9000 2039 13000 2081
rect 9000 1921 9073 2039
rect 9191 1921 12806 2039
rect 12924 1921 13000 2039
rect 9000 1879 13000 1921
rect 9000 1761 9073 1879
rect 9191 1761 12806 1879
rect 12924 1761 13000 1879
rect 9000 1719 13000 1761
rect 9000 1601 9073 1719
rect 9191 1601 12806 1719
rect 12924 1601 13000 1719
rect 9000 1559 13000 1601
rect 9000 1441 9073 1559
rect 9191 1441 12806 1559
rect 12924 1441 13000 1559
rect 9000 1399 13000 1441
rect 9000 1281 9073 1399
rect 9191 1281 12806 1399
rect 12924 1281 13000 1399
rect 9000 1239 13000 1281
rect 9000 1121 9073 1239
rect 9191 1121 12806 1239
rect 12924 1121 13000 1239
rect 9000 1079 13000 1121
rect 9000 961 9073 1079
rect 9191 961 12806 1079
rect 12924 961 13000 1079
rect 9000 919 13000 961
rect 9000 801 9073 919
rect 9191 801 12806 919
rect 12924 801 13000 919
rect 9000 759 13000 801
rect 9000 641 9073 759
rect 9191 641 12806 759
rect 12924 641 13000 759
rect 9000 599 13000 641
rect 9000 481 9073 599
rect 9191 481 12806 599
rect 12924 481 13000 599
rect 9000 439 13000 481
rect 9000 321 9073 439
rect 9191 321 12806 439
rect 12924 321 13000 439
rect 9000 279 13000 321
rect 9000 161 9073 279
rect 9191 161 12806 279
rect 12924 161 13000 279
rect 9000 119 13000 161
rect 9000 1 9073 119
rect 9191 1 12806 119
rect 12924 1 13000 119
rect 9000 -41 13000 1
rect 9000 -159 9073 -41
rect 9191 -159 12806 -41
rect 12924 -159 13000 -41
rect 9000 -201 13000 -159
rect 9000 -319 9073 -201
rect 9191 -304 12806 -201
rect 9191 -319 9261 -304
rect 9000 -422 9261 -319
rect 9379 -422 9421 -304
rect 9539 -422 9581 -304
rect 9699 -422 9741 -304
rect 9859 -422 9901 -304
rect 10019 -422 10061 -304
rect 10179 -422 10221 -304
rect 10339 -422 10381 -304
rect 10499 -422 10541 -304
rect 10659 -422 10701 -304
rect 10819 -422 10861 -304
rect 10979 -422 11021 -304
rect 11139 -422 11181 -304
rect 11299 -422 11341 -304
rect 11459 -422 11501 -304
rect 11619 -422 11661 -304
rect 11779 -422 11821 -304
rect 11939 -422 11981 -304
rect 12099 -422 12141 -304
rect 12259 -422 12301 -304
rect 12419 -422 12461 -304
rect 12579 -422 12621 -304
rect 12739 -319 12806 -304
rect 12924 -319 13000 -201
rect 12739 -422 13000 -319
rect 9000 -500 13000 -422
rect 15000 3424 19000 3500
rect 15000 3319 15261 3424
rect 15000 3201 15073 3319
rect 15191 3306 15261 3319
rect 15379 3306 15421 3424
rect 15539 3306 15581 3424
rect 15699 3306 15741 3424
rect 15859 3306 15901 3424
rect 16019 3306 16061 3424
rect 16179 3306 16221 3424
rect 16339 3306 16381 3424
rect 16499 3306 16541 3424
rect 16659 3306 16701 3424
rect 16819 3306 16861 3424
rect 16979 3306 17021 3424
rect 17139 3306 17181 3424
rect 17299 3306 17341 3424
rect 17459 3306 17501 3424
rect 17619 3306 17661 3424
rect 17779 3306 17821 3424
rect 17939 3306 17981 3424
rect 18099 3306 18141 3424
rect 18259 3306 18301 3424
rect 18419 3306 18461 3424
rect 18579 3306 18621 3424
rect 18739 3319 19000 3424
rect 18739 3306 18806 3319
rect 15191 3201 18806 3306
rect 18924 3201 19000 3319
rect 15000 3159 19000 3201
rect 15000 3041 15073 3159
rect 15191 3041 18806 3159
rect 18924 3041 19000 3159
rect 15000 2999 19000 3041
rect 15000 2881 15073 2999
rect 15191 2881 18806 2999
rect 18924 2881 19000 2999
rect 15000 2839 19000 2881
rect 15000 2721 15073 2839
rect 15191 2721 18806 2839
rect 18924 2721 19000 2839
rect 15000 2679 19000 2721
rect 15000 2561 15073 2679
rect 15191 2561 18806 2679
rect 18924 2561 19000 2679
rect 15000 2519 19000 2561
rect 15000 2401 15073 2519
rect 15191 2401 18806 2519
rect 18924 2401 19000 2519
rect 15000 2359 19000 2401
rect 15000 2241 15073 2359
rect 15191 2241 18806 2359
rect 18924 2241 19000 2359
rect 15000 2199 19000 2241
rect 15000 2081 15073 2199
rect 15191 2081 18806 2199
rect 18924 2081 19000 2199
rect 15000 2039 19000 2081
rect 15000 1921 15073 2039
rect 15191 1921 18806 2039
rect 18924 1921 19000 2039
rect 15000 1879 19000 1921
rect 15000 1761 15073 1879
rect 15191 1761 18806 1879
rect 18924 1761 19000 1879
rect 15000 1719 19000 1761
rect 15000 1601 15073 1719
rect 15191 1601 18806 1719
rect 18924 1601 19000 1719
rect 15000 1559 19000 1601
rect 15000 1441 15073 1559
rect 15191 1441 18806 1559
rect 18924 1441 19000 1559
rect 15000 1399 19000 1441
rect 15000 1281 15073 1399
rect 15191 1281 18806 1399
rect 18924 1281 19000 1399
rect 15000 1239 19000 1281
rect 15000 1121 15073 1239
rect 15191 1121 18806 1239
rect 18924 1121 19000 1239
rect 15000 1079 19000 1121
rect 15000 961 15073 1079
rect 15191 961 18806 1079
rect 18924 961 19000 1079
rect 15000 919 19000 961
rect 15000 801 15073 919
rect 15191 801 18806 919
rect 18924 801 19000 919
rect 15000 759 19000 801
rect 15000 641 15073 759
rect 15191 641 18806 759
rect 18924 641 19000 759
rect 15000 599 19000 641
rect 15000 481 15073 599
rect 15191 481 18806 599
rect 18924 481 19000 599
rect 15000 439 19000 481
rect 15000 321 15073 439
rect 15191 321 18806 439
rect 18924 321 19000 439
rect 15000 279 19000 321
rect 15000 161 15073 279
rect 15191 161 18806 279
rect 18924 161 19000 279
rect 15000 119 19000 161
rect 15000 1 15073 119
rect 15191 1 18806 119
rect 18924 1 19000 119
rect 15000 -41 19000 1
rect 15000 -159 15073 -41
rect 15191 -159 18806 -41
rect 18924 -159 19000 -41
rect 15000 -201 19000 -159
rect 15000 -319 15073 -201
rect 15191 -304 18806 -201
rect 15191 -319 15261 -304
rect 15000 -422 15261 -319
rect 15379 -422 15421 -304
rect 15539 -422 15581 -304
rect 15699 -422 15741 -304
rect 15859 -422 15901 -304
rect 16019 -422 16061 -304
rect 16179 -422 16221 -304
rect 16339 -422 16381 -304
rect 16499 -422 16541 -304
rect 16659 -422 16701 -304
rect 16819 -422 16861 -304
rect 16979 -422 17021 -304
rect 17139 -422 17181 -304
rect 17299 -422 17341 -304
rect 17459 -422 17501 -304
rect 17619 -422 17661 -304
rect 17779 -422 17821 -304
rect 17939 -422 17981 -304
rect 18099 -422 18141 -304
rect 18259 -422 18301 -304
rect 18419 -422 18461 -304
rect 18579 -422 18621 -304
rect 18739 -319 18806 -304
rect 18924 -319 19000 -201
rect 18739 -422 19000 -319
rect 15000 -500 19000 -422
rect 21000 3424 25000 3500
rect 21000 3319 21261 3424
rect 21000 3201 21073 3319
rect 21191 3306 21261 3319
rect 21379 3306 21421 3424
rect 21539 3306 21581 3424
rect 21699 3306 21741 3424
rect 21859 3306 21901 3424
rect 22019 3306 22061 3424
rect 22179 3306 22221 3424
rect 22339 3306 22381 3424
rect 22499 3306 22541 3424
rect 22659 3306 22701 3424
rect 22819 3306 22861 3424
rect 22979 3306 23021 3424
rect 23139 3306 23181 3424
rect 23299 3306 23341 3424
rect 23459 3306 23501 3424
rect 23619 3306 23661 3424
rect 23779 3306 23821 3424
rect 23939 3306 23981 3424
rect 24099 3306 24141 3424
rect 24259 3306 24301 3424
rect 24419 3306 24461 3424
rect 24579 3306 24621 3424
rect 24739 3319 25000 3424
rect 24739 3306 24806 3319
rect 21191 3201 24806 3306
rect 24924 3201 25000 3319
rect 21000 3159 25000 3201
rect 21000 3041 21073 3159
rect 21191 3041 24806 3159
rect 24924 3041 25000 3159
rect 21000 2999 25000 3041
rect 21000 2881 21073 2999
rect 21191 2881 24806 2999
rect 24924 2881 25000 2999
rect 21000 2839 25000 2881
rect 21000 2721 21073 2839
rect 21191 2721 24806 2839
rect 24924 2721 25000 2839
rect 21000 2679 25000 2721
rect 21000 2561 21073 2679
rect 21191 2561 24806 2679
rect 24924 2561 25000 2679
rect 21000 2519 25000 2561
rect 21000 2401 21073 2519
rect 21191 2401 24806 2519
rect 24924 2401 25000 2519
rect 21000 2359 25000 2401
rect 21000 2241 21073 2359
rect 21191 2241 24806 2359
rect 24924 2241 25000 2359
rect 21000 2199 25000 2241
rect 21000 2081 21073 2199
rect 21191 2081 24806 2199
rect 24924 2081 25000 2199
rect 21000 2039 25000 2081
rect 21000 1921 21073 2039
rect 21191 1921 24806 2039
rect 24924 1921 25000 2039
rect 21000 1879 25000 1921
rect 21000 1761 21073 1879
rect 21191 1761 24806 1879
rect 24924 1761 25000 1879
rect 21000 1719 25000 1761
rect 21000 1601 21073 1719
rect 21191 1601 24806 1719
rect 24924 1601 25000 1719
rect 21000 1559 25000 1601
rect 21000 1441 21073 1559
rect 21191 1441 24806 1559
rect 24924 1441 25000 1559
rect 21000 1399 25000 1441
rect 21000 1281 21073 1399
rect 21191 1281 24806 1399
rect 24924 1281 25000 1399
rect 21000 1239 25000 1281
rect 21000 1121 21073 1239
rect 21191 1121 24806 1239
rect 24924 1121 25000 1239
rect 21000 1079 25000 1121
rect 21000 961 21073 1079
rect 21191 961 24806 1079
rect 24924 961 25000 1079
rect 21000 919 25000 961
rect 21000 801 21073 919
rect 21191 801 24806 919
rect 24924 801 25000 919
rect 21000 759 25000 801
rect 21000 641 21073 759
rect 21191 641 24806 759
rect 24924 641 25000 759
rect 21000 599 25000 641
rect 21000 481 21073 599
rect 21191 481 24806 599
rect 24924 481 25000 599
rect 21000 439 25000 481
rect 21000 321 21073 439
rect 21191 321 24806 439
rect 24924 321 25000 439
rect 21000 279 25000 321
rect 21000 161 21073 279
rect 21191 161 24806 279
rect 24924 161 25000 279
rect 21000 119 25000 161
rect 21000 1 21073 119
rect 21191 1 24806 119
rect 24924 1 25000 119
rect 21000 -41 25000 1
rect 21000 -159 21073 -41
rect 21191 -159 24806 -41
rect 24924 -159 25000 -41
rect 21000 -201 25000 -159
rect 21000 -319 21073 -201
rect 21191 -304 24806 -201
rect 21191 -319 21261 -304
rect 21000 -422 21261 -319
rect 21379 -422 21421 -304
rect 21539 -422 21581 -304
rect 21699 -422 21741 -304
rect 21859 -422 21901 -304
rect 22019 -422 22061 -304
rect 22179 -422 22221 -304
rect 22339 -422 22381 -304
rect 22499 -422 22541 -304
rect 22659 -422 22701 -304
rect 22819 -422 22861 -304
rect 22979 -422 23021 -304
rect 23139 -422 23181 -304
rect 23299 -422 23341 -304
rect 23459 -422 23501 -304
rect 23619 -422 23661 -304
rect 23779 -422 23821 -304
rect 23939 -422 23981 -304
rect 24099 -422 24141 -304
rect 24259 -422 24301 -304
rect 24419 -422 24461 -304
rect 24579 -422 24621 -304
rect 24739 -319 24806 -304
rect 24924 -319 25000 -201
rect 24739 -422 25000 -319
rect 21000 -500 25000 -422
rect 22900 -1100 23100 -700
rect 22100 -1500 22300 -1100
rect 22500 -1500 22700 -1100
rect 22100 -1700 22700 -1500
rect 22900 -1300 23500 -1100
rect 22900 -1700 23100 -1300
rect 23300 -1700 23500 -1300
rect 23700 -1300 24300 -1100
rect 22100 -1900 22300 -1700
rect 22500 -1900 22700 -1700
rect 22100 -2100 22700 -1900
rect 23700 -1900 23900 -1300
rect 24100 -1900 24300 -1300
rect 23700 -2100 24300 -1900
rect 24500 -1500 24700 -1100
rect 25300 -1500 25500 -1100
rect 24500 -1700 25100 -1500
rect 24500 -2100 24700 -1700
rect 24900 -2100 25100 -1700
rect 25300 -1700 25900 -1500
rect 25300 -2100 25500 -1700
rect 25700 -2100 25900 -1700
rect 2300 -4100 2900 -3900
rect 3100 -4100 3700 -3900
rect 2700 -4300 2900 -4100
rect 3500 -4300 3700 -4100
rect 2300 -4500 2900 -4300
rect 3100 -4500 3700 -4300
rect 3900 -4100 4500 -3900
rect 2300 -4700 2500 -4500
rect 3100 -4700 3300 -4500
rect 3900 -4700 4100 -4100
rect 4300 -4700 4500 -4100
rect 5500 -4100 6100 -3900
rect 5500 -4300 5700 -4100
rect 5900 -4300 6100 -4100
rect 2300 -4900 2900 -4700
rect 3100 -4900 3700 -4700
rect 3900 -4900 4500 -4700
rect 4700 -4700 4900 -4300
rect 5100 -4700 5300 -4300
rect 4700 -4900 5300 -4700
rect 5500 -4500 6100 -4300
rect 5500 -4900 5700 -4500
rect 5900 -4900 6100 -4500
rect 5100 -5300 5300 -4900
rect 3000 -5578 7000 -5500
rect 3000 -5681 3261 -5578
rect 3000 -5799 3076 -5681
rect 3194 -5696 3261 -5681
rect 3379 -5696 3421 -5578
rect 3539 -5696 3581 -5578
rect 3699 -5696 3741 -5578
rect 3859 -5696 3901 -5578
rect 4019 -5696 4061 -5578
rect 4179 -5696 4221 -5578
rect 4339 -5696 4381 -5578
rect 4499 -5696 4541 -5578
rect 4659 -5696 4701 -5578
rect 4819 -5696 4861 -5578
rect 4979 -5696 5021 -5578
rect 5139 -5696 5181 -5578
rect 5299 -5696 5341 -5578
rect 5459 -5696 5501 -5578
rect 5619 -5696 5661 -5578
rect 5779 -5696 5821 -5578
rect 5939 -5696 5981 -5578
rect 6099 -5696 6141 -5578
rect 6259 -5696 6301 -5578
rect 6419 -5696 6461 -5578
rect 6579 -5696 6621 -5578
rect 6739 -5681 7000 -5578
rect 6739 -5696 6809 -5681
rect 3194 -5799 6809 -5696
rect 6927 -5799 7000 -5681
rect 3000 -5841 7000 -5799
rect 3000 -5959 3076 -5841
rect 3194 -5959 6809 -5841
rect 6927 -5959 7000 -5841
rect 3000 -6001 7000 -5959
rect 3000 -6119 3076 -6001
rect 3194 -6119 6809 -6001
rect 6927 -6119 7000 -6001
rect 3000 -6161 7000 -6119
rect 3000 -6279 3076 -6161
rect 3194 -6279 6809 -6161
rect 6927 -6279 7000 -6161
rect 3000 -6321 7000 -6279
rect 3000 -6439 3076 -6321
rect 3194 -6439 6809 -6321
rect 6927 -6439 7000 -6321
rect 3000 -6481 7000 -6439
rect 3000 -6599 3076 -6481
rect 3194 -6599 6809 -6481
rect 6927 -6599 7000 -6481
rect 3000 -6641 7000 -6599
rect 3000 -6759 3076 -6641
rect 3194 -6759 6809 -6641
rect 6927 -6759 7000 -6641
rect 3000 -6801 7000 -6759
rect 3000 -6919 3076 -6801
rect 3194 -6919 6809 -6801
rect 6927 -6919 7000 -6801
rect 3000 -6961 7000 -6919
rect 3000 -7079 3076 -6961
rect 3194 -7079 6809 -6961
rect 6927 -7079 7000 -6961
rect 3000 -7121 7000 -7079
rect 3000 -7239 3076 -7121
rect 3194 -7239 6809 -7121
rect 6927 -7239 7000 -7121
rect 3000 -7281 7000 -7239
rect 3000 -7399 3076 -7281
rect 3194 -7399 6809 -7281
rect 6927 -7399 7000 -7281
rect 3000 -7441 7000 -7399
rect 3000 -7559 3076 -7441
rect 3194 -7559 6809 -7441
rect 6927 -7559 7000 -7441
rect 3000 -7601 7000 -7559
rect 3000 -7719 3076 -7601
rect 3194 -7719 6809 -7601
rect 6927 -7719 7000 -7601
rect 3000 -7761 7000 -7719
rect 3000 -7879 3076 -7761
rect 3194 -7879 6809 -7761
rect 6927 -7879 7000 -7761
rect 3000 -7921 7000 -7879
rect 3000 -8039 3076 -7921
rect 3194 -8039 6809 -7921
rect 6927 -8039 7000 -7921
rect 3000 -8081 7000 -8039
rect 3000 -8199 3076 -8081
rect 3194 -8199 6809 -8081
rect 6927 -8199 7000 -8081
rect 3000 -8241 7000 -8199
rect 3000 -8359 3076 -8241
rect 3194 -8359 6809 -8241
rect 6927 -8359 7000 -8241
rect 3000 -8401 7000 -8359
rect 3000 -8519 3076 -8401
rect 3194 -8519 6809 -8401
rect 6927 -8519 7000 -8401
rect 3000 -8561 7000 -8519
rect 3000 -8679 3076 -8561
rect 3194 -8679 6809 -8561
rect 6927 -8679 7000 -8561
rect 3000 -8721 7000 -8679
rect 3000 -8839 3076 -8721
rect 3194 -8839 6809 -8721
rect 6927 -8839 7000 -8721
rect 3000 -8881 7000 -8839
rect 3000 -8999 3076 -8881
rect 3194 -8999 6809 -8881
rect 6927 -8999 7000 -8881
rect 3000 -9041 7000 -8999
rect 3000 -9159 3076 -9041
rect 3194 -9159 6809 -9041
rect 6927 -9159 7000 -9041
rect 3000 -9201 7000 -9159
rect 3000 -9319 3076 -9201
rect 3194 -9306 6809 -9201
rect 3194 -9319 3261 -9306
rect 3000 -9424 3261 -9319
rect 3379 -9424 3421 -9306
rect 3539 -9424 3581 -9306
rect 3699 -9424 3741 -9306
rect 3859 -9424 3901 -9306
rect 4019 -9424 4061 -9306
rect 4179 -9424 4221 -9306
rect 4339 -9424 4381 -9306
rect 4499 -9424 4541 -9306
rect 4659 -9424 4701 -9306
rect 4819 -9424 4861 -9306
rect 4979 -9424 5021 -9306
rect 5139 -9424 5181 -9306
rect 5299 -9424 5341 -9306
rect 5459 -9424 5501 -9306
rect 5619 -9424 5661 -9306
rect 5779 -9424 5821 -9306
rect 5939 -9424 5981 -9306
rect 6099 -9424 6141 -9306
rect 6259 -9424 6301 -9306
rect 6419 -9424 6461 -9306
rect 6579 -9424 6621 -9306
rect 6739 -9319 6809 -9306
rect 6927 -9319 7000 -9201
rect 6739 -9424 7000 -9319
rect 3000 -9500 7000 -9424
rect 9000 -5578 13000 -5500
rect 9000 -5681 9261 -5578
rect 9000 -5799 9076 -5681
rect 9194 -5696 9261 -5681
rect 9379 -5696 9421 -5578
rect 9539 -5696 9581 -5578
rect 9699 -5696 9741 -5578
rect 9859 -5696 9901 -5578
rect 10019 -5696 10061 -5578
rect 10179 -5696 10221 -5578
rect 10339 -5696 10381 -5578
rect 10499 -5696 10541 -5578
rect 10659 -5696 10701 -5578
rect 10819 -5696 10861 -5578
rect 10979 -5696 11021 -5578
rect 11139 -5696 11181 -5578
rect 11299 -5696 11341 -5578
rect 11459 -5696 11501 -5578
rect 11619 -5696 11661 -5578
rect 11779 -5696 11821 -5578
rect 11939 -5696 11981 -5578
rect 12099 -5696 12141 -5578
rect 12259 -5696 12301 -5578
rect 12419 -5696 12461 -5578
rect 12579 -5696 12621 -5578
rect 12739 -5681 13000 -5578
rect 12739 -5696 12809 -5681
rect 9194 -5799 12809 -5696
rect 12927 -5799 13000 -5681
rect 9000 -5841 13000 -5799
rect 9000 -5959 9076 -5841
rect 9194 -5959 12809 -5841
rect 12927 -5959 13000 -5841
rect 9000 -6001 13000 -5959
rect 9000 -6119 9076 -6001
rect 9194 -6119 12809 -6001
rect 12927 -6119 13000 -6001
rect 9000 -6161 13000 -6119
rect 9000 -6279 9076 -6161
rect 9194 -6279 12809 -6161
rect 12927 -6279 13000 -6161
rect 9000 -6321 13000 -6279
rect 9000 -6439 9076 -6321
rect 9194 -6439 12809 -6321
rect 12927 -6439 13000 -6321
rect 9000 -6481 13000 -6439
rect 9000 -6599 9076 -6481
rect 9194 -6599 12809 -6481
rect 12927 -6599 13000 -6481
rect 9000 -6641 13000 -6599
rect 9000 -6759 9076 -6641
rect 9194 -6759 12809 -6641
rect 12927 -6759 13000 -6641
rect 9000 -6801 13000 -6759
rect 9000 -6919 9076 -6801
rect 9194 -6919 12809 -6801
rect 12927 -6919 13000 -6801
rect 9000 -6961 13000 -6919
rect 9000 -7079 9076 -6961
rect 9194 -7079 12809 -6961
rect 12927 -7079 13000 -6961
rect 9000 -7121 13000 -7079
rect 9000 -7239 9076 -7121
rect 9194 -7239 12809 -7121
rect 12927 -7239 13000 -7121
rect 9000 -7281 13000 -7239
rect 9000 -7399 9076 -7281
rect 9194 -7399 12809 -7281
rect 12927 -7399 13000 -7281
rect 9000 -7441 13000 -7399
rect 9000 -7559 9076 -7441
rect 9194 -7559 12809 -7441
rect 12927 -7559 13000 -7441
rect 9000 -7601 13000 -7559
rect 9000 -7719 9076 -7601
rect 9194 -7719 12809 -7601
rect 12927 -7719 13000 -7601
rect 9000 -7761 13000 -7719
rect 9000 -7879 9076 -7761
rect 9194 -7879 12809 -7761
rect 12927 -7879 13000 -7761
rect 9000 -7921 13000 -7879
rect 9000 -8039 9076 -7921
rect 9194 -8039 12809 -7921
rect 12927 -8039 13000 -7921
rect 9000 -8081 13000 -8039
rect 9000 -8199 9076 -8081
rect 9194 -8199 12809 -8081
rect 12927 -8199 13000 -8081
rect 9000 -8241 13000 -8199
rect 9000 -8359 9076 -8241
rect 9194 -8359 12809 -8241
rect 12927 -8359 13000 -8241
rect 9000 -8401 13000 -8359
rect 9000 -8519 9076 -8401
rect 9194 -8519 12809 -8401
rect 12927 -8519 13000 -8401
rect 9000 -8561 13000 -8519
rect 9000 -8679 9076 -8561
rect 9194 -8679 12809 -8561
rect 12927 -8679 13000 -8561
rect 9000 -8721 13000 -8679
rect 9000 -8839 9076 -8721
rect 9194 -8839 12809 -8721
rect 12927 -8839 13000 -8721
rect 9000 -8881 13000 -8839
rect 9000 -8999 9076 -8881
rect 9194 -8999 12809 -8881
rect 12927 -8999 13000 -8881
rect 9000 -9041 13000 -8999
rect 9000 -9159 9076 -9041
rect 9194 -9159 12809 -9041
rect 12927 -9159 13000 -9041
rect 9000 -9201 13000 -9159
rect 9000 -9319 9076 -9201
rect 9194 -9306 12809 -9201
rect 9194 -9319 9261 -9306
rect 9000 -9424 9261 -9319
rect 9379 -9424 9421 -9306
rect 9539 -9424 9581 -9306
rect 9699 -9424 9741 -9306
rect 9859 -9424 9901 -9306
rect 10019 -9424 10061 -9306
rect 10179 -9424 10221 -9306
rect 10339 -9424 10381 -9306
rect 10499 -9424 10541 -9306
rect 10659 -9424 10701 -9306
rect 10819 -9424 10861 -9306
rect 10979 -9424 11021 -9306
rect 11139 -9424 11181 -9306
rect 11299 -9424 11341 -9306
rect 11459 -9424 11501 -9306
rect 11619 -9424 11661 -9306
rect 11779 -9424 11821 -9306
rect 11939 -9424 11981 -9306
rect 12099 -9424 12141 -9306
rect 12259 -9424 12301 -9306
rect 12419 -9424 12461 -9306
rect 12579 -9424 12621 -9306
rect 12739 -9319 12809 -9306
rect 12927 -9319 13000 -9201
rect 12739 -9424 13000 -9319
rect 9000 -9500 13000 -9424
rect 15000 -5578 19000 -5500
rect 15000 -5681 15261 -5578
rect 15000 -5799 15076 -5681
rect 15194 -5696 15261 -5681
rect 15379 -5696 15421 -5578
rect 15539 -5696 15581 -5578
rect 15699 -5696 15741 -5578
rect 15859 -5696 15901 -5578
rect 16019 -5696 16061 -5578
rect 16179 -5696 16221 -5578
rect 16339 -5696 16381 -5578
rect 16499 -5696 16541 -5578
rect 16659 -5696 16701 -5578
rect 16819 -5696 16861 -5578
rect 16979 -5696 17021 -5578
rect 17139 -5696 17181 -5578
rect 17299 -5696 17341 -5578
rect 17459 -5696 17501 -5578
rect 17619 -5696 17661 -5578
rect 17779 -5696 17821 -5578
rect 17939 -5696 17981 -5578
rect 18099 -5696 18141 -5578
rect 18259 -5696 18301 -5578
rect 18419 -5696 18461 -5578
rect 18579 -5696 18621 -5578
rect 18739 -5681 19000 -5578
rect 18739 -5696 18809 -5681
rect 15194 -5799 18809 -5696
rect 18927 -5799 19000 -5681
rect 15000 -5841 19000 -5799
rect 15000 -5959 15076 -5841
rect 15194 -5959 18809 -5841
rect 18927 -5959 19000 -5841
rect 15000 -6001 19000 -5959
rect 15000 -6119 15076 -6001
rect 15194 -6119 18809 -6001
rect 18927 -6119 19000 -6001
rect 15000 -6161 19000 -6119
rect 15000 -6279 15076 -6161
rect 15194 -6279 18809 -6161
rect 18927 -6279 19000 -6161
rect 15000 -6321 19000 -6279
rect 15000 -6439 15076 -6321
rect 15194 -6439 18809 -6321
rect 18927 -6439 19000 -6321
rect 15000 -6481 19000 -6439
rect 15000 -6599 15076 -6481
rect 15194 -6599 18809 -6481
rect 18927 -6599 19000 -6481
rect 15000 -6641 19000 -6599
rect 15000 -6759 15076 -6641
rect 15194 -6759 18809 -6641
rect 18927 -6759 19000 -6641
rect 15000 -6801 19000 -6759
rect 15000 -6919 15076 -6801
rect 15194 -6919 18809 -6801
rect 18927 -6919 19000 -6801
rect 15000 -6961 19000 -6919
rect 15000 -7079 15076 -6961
rect 15194 -7079 18809 -6961
rect 18927 -7079 19000 -6961
rect 15000 -7121 19000 -7079
rect 15000 -7239 15076 -7121
rect 15194 -7239 18809 -7121
rect 18927 -7239 19000 -7121
rect 15000 -7281 19000 -7239
rect 15000 -7399 15076 -7281
rect 15194 -7399 18809 -7281
rect 18927 -7399 19000 -7281
rect 15000 -7441 19000 -7399
rect 15000 -7559 15076 -7441
rect 15194 -7559 18809 -7441
rect 18927 -7559 19000 -7441
rect 15000 -7601 19000 -7559
rect 15000 -7719 15076 -7601
rect 15194 -7719 18809 -7601
rect 18927 -7719 19000 -7601
rect 15000 -7761 19000 -7719
rect 15000 -7879 15076 -7761
rect 15194 -7879 18809 -7761
rect 18927 -7879 19000 -7761
rect 15000 -7921 19000 -7879
rect 15000 -8039 15076 -7921
rect 15194 -8039 18809 -7921
rect 18927 -8039 19000 -7921
rect 15000 -8081 19000 -8039
rect 15000 -8199 15076 -8081
rect 15194 -8199 18809 -8081
rect 18927 -8199 19000 -8081
rect 15000 -8241 19000 -8199
rect 15000 -8359 15076 -8241
rect 15194 -8359 18809 -8241
rect 18927 -8359 19000 -8241
rect 15000 -8401 19000 -8359
rect 15000 -8519 15076 -8401
rect 15194 -8519 18809 -8401
rect 18927 -8519 19000 -8401
rect 15000 -8561 19000 -8519
rect 15000 -8679 15076 -8561
rect 15194 -8679 18809 -8561
rect 18927 -8679 19000 -8561
rect 15000 -8721 19000 -8679
rect 15000 -8839 15076 -8721
rect 15194 -8839 18809 -8721
rect 18927 -8839 19000 -8721
rect 15000 -8881 19000 -8839
rect 15000 -8999 15076 -8881
rect 15194 -8999 18809 -8881
rect 18927 -8999 19000 -8881
rect 15000 -9041 19000 -8999
rect 15000 -9159 15076 -9041
rect 15194 -9159 18809 -9041
rect 18927 -9159 19000 -9041
rect 15000 -9201 19000 -9159
rect 15000 -9319 15076 -9201
rect 15194 -9306 18809 -9201
rect 15194 -9319 15261 -9306
rect 15000 -9424 15261 -9319
rect 15379 -9424 15421 -9306
rect 15539 -9424 15581 -9306
rect 15699 -9424 15741 -9306
rect 15859 -9424 15901 -9306
rect 16019 -9424 16061 -9306
rect 16179 -9424 16221 -9306
rect 16339 -9424 16381 -9306
rect 16499 -9424 16541 -9306
rect 16659 -9424 16701 -9306
rect 16819 -9424 16861 -9306
rect 16979 -9424 17021 -9306
rect 17139 -9424 17181 -9306
rect 17299 -9424 17341 -9306
rect 17459 -9424 17501 -9306
rect 17619 -9424 17661 -9306
rect 17779 -9424 17821 -9306
rect 17939 -9424 17981 -9306
rect 18099 -9424 18141 -9306
rect 18259 -9424 18301 -9306
rect 18419 -9424 18461 -9306
rect 18579 -9424 18621 -9306
rect 18739 -9319 18809 -9306
rect 18927 -9319 19000 -9201
rect 18739 -9424 19000 -9319
rect 15000 -9500 19000 -9424
rect 21000 -5578 25000 -5500
rect 21000 -5681 21261 -5578
rect 21000 -5799 21076 -5681
rect 21194 -5696 21261 -5681
rect 21379 -5696 21421 -5578
rect 21539 -5696 21581 -5578
rect 21699 -5696 21741 -5578
rect 21859 -5696 21901 -5578
rect 22019 -5696 22061 -5578
rect 22179 -5696 22221 -5578
rect 22339 -5696 22381 -5578
rect 22499 -5696 22541 -5578
rect 22659 -5696 22701 -5578
rect 22819 -5696 22861 -5578
rect 22979 -5696 23021 -5578
rect 23139 -5696 23181 -5578
rect 23299 -5696 23341 -5578
rect 23459 -5696 23501 -5578
rect 23619 -5696 23661 -5578
rect 23779 -5696 23821 -5578
rect 23939 -5696 23981 -5578
rect 24099 -5696 24141 -5578
rect 24259 -5696 24301 -5578
rect 24419 -5696 24461 -5578
rect 24579 -5696 24621 -5578
rect 24739 -5681 25000 -5578
rect 24739 -5696 24809 -5681
rect 21194 -5799 24809 -5696
rect 24927 -5799 25000 -5681
rect 21000 -5841 25000 -5799
rect 21000 -5959 21076 -5841
rect 21194 -5959 24809 -5841
rect 24927 -5959 25000 -5841
rect 21000 -6001 25000 -5959
rect 21000 -6119 21076 -6001
rect 21194 -6119 24809 -6001
rect 24927 -6119 25000 -6001
rect 21000 -6161 25000 -6119
rect 21000 -6279 21076 -6161
rect 21194 -6279 24809 -6161
rect 24927 -6279 25000 -6161
rect 21000 -6321 25000 -6279
rect 21000 -6439 21076 -6321
rect 21194 -6439 24809 -6321
rect 24927 -6439 25000 -6321
rect 21000 -6481 25000 -6439
rect 21000 -6599 21076 -6481
rect 21194 -6599 24809 -6481
rect 24927 -6599 25000 -6481
rect 21000 -6641 25000 -6599
rect 21000 -6759 21076 -6641
rect 21194 -6759 24809 -6641
rect 24927 -6759 25000 -6641
rect 21000 -6801 25000 -6759
rect 21000 -6919 21076 -6801
rect 21194 -6919 24809 -6801
rect 24927 -6919 25000 -6801
rect 21000 -6961 25000 -6919
rect 21000 -7079 21076 -6961
rect 21194 -7079 24809 -6961
rect 24927 -7079 25000 -6961
rect 21000 -7121 25000 -7079
rect 21000 -7239 21076 -7121
rect 21194 -7239 24809 -7121
rect 24927 -7239 25000 -7121
rect 21000 -7281 25000 -7239
rect 21000 -7399 21076 -7281
rect 21194 -7399 24809 -7281
rect 24927 -7399 25000 -7281
rect 21000 -7441 25000 -7399
rect 21000 -7559 21076 -7441
rect 21194 -7559 24809 -7441
rect 24927 -7559 25000 -7441
rect 21000 -7601 25000 -7559
rect 21000 -7719 21076 -7601
rect 21194 -7719 24809 -7601
rect 24927 -7719 25000 -7601
rect 21000 -7761 25000 -7719
rect 21000 -7879 21076 -7761
rect 21194 -7879 24809 -7761
rect 24927 -7879 25000 -7761
rect 21000 -7921 25000 -7879
rect 21000 -8039 21076 -7921
rect 21194 -8039 24809 -7921
rect 24927 -8039 25000 -7921
rect 21000 -8081 25000 -8039
rect 21000 -8199 21076 -8081
rect 21194 -8199 24809 -8081
rect 24927 -8199 25000 -8081
rect 21000 -8241 25000 -8199
rect 21000 -8359 21076 -8241
rect 21194 -8359 24809 -8241
rect 24927 -8359 25000 -8241
rect 21000 -8401 25000 -8359
rect 21000 -8519 21076 -8401
rect 21194 -8519 24809 -8401
rect 24927 -8519 25000 -8401
rect 21000 -8561 25000 -8519
rect 21000 -8679 21076 -8561
rect 21194 -8679 24809 -8561
rect 24927 -8679 25000 -8561
rect 21000 -8721 25000 -8679
rect 21000 -8839 21076 -8721
rect 21194 -8839 24809 -8721
rect 24927 -8839 25000 -8721
rect 21000 -8881 25000 -8839
rect 21000 -8999 21076 -8881
rect 21194 -8999 24809 -8881
rect 24927 -8999 25000 -8881
rect 21000 -9041 25000 -8999
rect 21000 -9159 21076 -9041
rect 21194 -9159 24809 -9041
rect 24927 -9159 25000 -9041
rect 21000 -9201 25000 -9159
rect 21000 -9319 21076 -9201
rect 21194 -9306 24809 -9201
rect 21194 -9319 21261 -9306
rect 21000 -9424 21261 -9319
rect 21379 -9424 21421 -9306
rect 21539 -9424 21581 -9306
rect 21699 -9424 21741 -9306
rect 21859 -9424 21901 -9306
rect 22019 -9424 22061 -9306
rect 22179 -9424 22221 -9306
rect 22339 -9424 22381 -9306
rect 22499 -9424 22541 -9306
rect 22659 -9424 22701 -9306
rect 22819 -9424 22861 -9306
rect 22979 -9424 23021 -9306
rect 23139 -9424 23181 -9306
rect 23299 -9424 23341 -9306
rect 23459 -9424 23501 -9306
rect 23619 -9424 23661 -9306
rect 23779 -9424 23821 -9306
rect 23939 -9424 23981 -9306
rect 24099 -9424 24141 -9306
rect 24259 -9424 24301 -9306
rect 24419 -9424 24461 -9306
rect 24579 -9424 24621 -9306
rect 24739 -9319 24809 -9306
rect 24927 -9319 25000 -9201
rect 24739 -9424 25000 -9319
rect 21000 -9500 25000 -9424
rect 3000 -11578 7000 -11500
rect 3000 -11681 3261 -11578
rect 3000 -11799 3076 -11681
rect 3194 -11696 3261 -11681
rect 3379 -11696 3421 -11578
rect 3539 -11696 3581 -11578
rect 3699 -11696 3741 -11578
rect 3859 -11696 3901 -11578
rect 4019 -11696 4061 -11578
rect 4179 -11696 4221 -11578
rect 4339 -11696 4381 -11578
rect 4499 -11696 4541 -11578
rect 4659 -11696 4701 -11578
rect 4819 -11696 4861 -11578
rect 4979 -11696 5021 -11578
rect 5139 -11696 5181 -11578
rect 5299 -11696 5341 -11578
rect 5459 -11696 5501 -11578
rect 5619 -11696 5661 -11578
rect 5779 -11696 5821 -11578
rect 5939 -11696 5981 -11578
rect 6099 -11696 6141 -11578
rect 6259 -11696 6301 -11578
rect 6419 -11696 6461 -11578
rect 6579 -11696 6621 -11578
rect 6739 -11681 7000 -11578
rect 6739 -11696 6809 -11681
rect 3194 -11799 6809 -11696
rect 6927 -11799 7000 -11681
rect 3000 -11841 7000 -11799
rect 3000 -11959 3076 -11841
rect 3194 -11959 6809 -11841
rect 6927 -11959 7000 -11841
rect 3000 -12001 7000 -11959
rect 3000 -12119 3076 -12001
rect 3194 -12119 6809 -12001
rect 6927 -12119 7000 -12001
rect 3000 -12161 7000 -12119
rect 3000 -12279 3076 -12161
rect 3194 -12279 6809 -12161
rect 6927 -12279 7000 -12161
rect 3000 -12321 7000 -12279
rect 3000 -12439 3076 -12321
rect 3194 -12439 6809 -12321
rect 6927 -12439 7000 -12321
rect 3000 -12481 7000 -12439
rect 3000 -12599 3076 -12481
rect 3194 -12599 6809 -12481
rect 6927 -12599 7000 -12481
rect 3000 -12641 7000 -12599
rect 3000 -12759 3076 -12641
rect 3194 -12759 6809 -12641
rect 6927 -12759 7000 -12641
rect 3000 -12801 7000 -12759
rect 3000 -12919 3076 -12801
rect 3194 -12919 6809 -12801
rect 6927 -12919 7000 -12801
rect 3000 -12961 7000 -12919
rect 3000 -13079 3076 -12961
rect 3194 -13079 6809 -12961
rect 6927 -13079 7000 -12961
rect 3000 -13121 7000 -13079
rect 3000 -13239 3076 -13121
rect 3194 -13239 6809 -13121
rect 6927 -13239 7000 -13121
rect 3000 -13281 7000 -13239
rect 3000 -13399 3076 -13281
rect 3194 -13399 6809 -13281
rect 6927 -13399 7000 -13281
rect 3000 -13441 7000 -13399
rect 3000 -13559 3076 -13441
rect 3194 -13559 6809 -13441
rect 6927 -13559 7000 -13441
rect 3000 -13601 7000 -13559
rect 3000 -13719 3076 -13601
rect 3194 -13719 6809 -13601
rect 6927 -13719 7000 -13601
rect 3000 -13761 7000 -13719
rect 3000 -13879 3076 -13761
rect 3194 -13879 6809 -13761
rect 6927 -13879 7000 -13761
rect 3000 -13921 7000 -13879
rect 3000 -14039 3076 -13921
rect 3194 -14039 6809 -13921
rect 6927 -14039 7000 -13921
rect 3000 -14081 7000 -14039
rect 3000 -14199 3076 -14081
rect 3194 -14199 6809 -14081
rect 6927 -14199 7000 -14081
rect 3000 -14241 7000 -14199
rect 3000 -14359 3076 -14241
rect 3194 -14359 6809 -14241
rect 6927 -14359 7000 -14241
rect 3000 -14401 7000 -14359
rect 3000 -14519 3076 -14401
rect 3194 -14519 6809 -14401
rect 6927 -14519 7000 -14401
rect 3000 -14561 7000 -14519
rect 3000 -14679 3076 -14561
rect 3194 -14679 6809 -14561
rect 6927 -14679 7000 -14561
rect 3000 -14721 7000 -14679
rect 3000 -14839 3076 -14721
rect 3194 -14839 6809 -14721
rect 6927 -14839 7000 -14721
rect 3000 -14881 7000 -14839
rect 3000 -14999 3076 -14881
rect 3194 -14999 6809 -14881
rect 6927 -14999 7000 -14881
rect 3000 -15041 7000 -14999
rect 3000 -15159 3076 -15041
rect 3194 -15159 6809 -15041
rect 6927 -15159 7000 -15041
rect 3000 -15201 7000 -15159
rect 3000 -15319 3076 -15201
rect 3194 -15306 6809 -15201
rect 3194 -15319 3261 -15306
rect 3000 -15424 3261 -15319
rect 3379 -15424 3421 -15306
rect 3539 -15424 3581 -15306
rect 3699 -15424 3741 -15306
rect 3859 -15424 3901 -15306
rect 4019 -15424 4061 -15306
rect 4179 -15424 4221 -15306
rect 4339 -15424 4381 -15306
rect 4499 -15424 4541 -15306
rect 4659 -15424 4701 -15306
rect 4819 -15424 4861 -15306
rect 4979 -15424 5021 -15306
rect 5139 -15424 5181 -15306
rect 5299 -15424 5341 -15306
rect 5459 -15424 5501 -15306
rect 5619 -15424 5661 -15306
rect 5779 -15424 5821 -15306
rect 5939 -15424 5981 -15306
rect 6099 -15424 6141 -15306
rect 6259 -15424 6301 -15306
rect 6419 -15424 6461 -15306
rect 6579 -15424 6621 -15306
rect 6739 -15319 6809 -15306
rect 6927 -15319 7000 -15201
rect 6739 -15424 7000 -15319
rect 3000 -15500 7000 -15424
rect 9000 -11578 13000 -11500
rect 9000 -11681 9261 -11578
rect 9000 -11799 9076 -11681
rect 9194 -11696 9261 -11681
rect 9379 -11696 9421 -11578
rect 9539 -11696 9581 -11578
rect 9699 -11696 9741 -11578
rect 9859 -11696 9901 -11578
rect 10019 -11696 10061 -11578
rect 10179 -11696 10221 -11578
rect 10339 -11696 10381 -11578
rect 10499 -11696 10541 -11578
rect 10659 -11696 10701 -11578
rect 10819 -11696 10861 -11578
rect 10979 -11696 11021 -11578
rect 11139 -11696 11181 -11578
rect 11299 -11696 11341 -11578
rect 11459 -11696 11501 -11578
rect 11619 -11696 11661 -11578
rect 11779 -11696 11821 -11578
rect 11939 -11696 11981 -11578
rect 12099 -11696 12141 -11578
rect 12259 -11696 12301 -11578
rect 12419 -11696 12461 -11578
rect 12579 -11696 12621 -11578
rect 12739 -11681 13000 -11578
rect 12739 -11696 12809 -11681
rect 9194 -11799 12809 -11696
rect 12927 -11799 13000 -11681
rect 9000 -11841 13000 -11799
rect 9000 -11959 9076 -11841
rect 9194 -11959 12809 -11841
rect 12927 -11959 13000 -11841
rect 9000 -12001 13000 -11959
rect 9000 -12119 9076 -12001
rect 9194 -12119 12809 -12001
rect 12927 -12119 13000 -12001
rect 9000 -12161 13000 -12119
rect 9000 -12279 9076 -12161
rect 9194 -12279 12809 -12161
rect 12927 -12279 13000 -12161
rect 9000 -12321 13000 -12279
rect 9000 -12439 9076 -12321
rect 9194 -12439 12809 -12321
rect 12927 -12439 13000 -12321
rect 9000 -12481 13000 -12439
rect 9000 -12599 9076 -12481
rect 9194 -12599 12809 -12481
rect 12927 -12599 13000 -12481
rect 9000 -12641 13000 -12599
rect 9000 -12759 9076 -12641
rect 9194 -12759 12809 -12641
rect 12927 -12759 13000 -12641
rect 9000 -12801 13000 -12759
rect 9000 -12919 9076 -12801
rect 9194 -12919 12809 -12801
rect 12927 -12919 13000 -12801
rect 9000 -12961 13000 -12919
rect 9000 -13079 9076 -12961
rect 9194 -13079 12809 -12961
rect 12927 -13079 13000 -12961
rect 9000 -13121 13000 -13079
rect 9000 -13239 9076 -13121
rect 9194 -13239 12809 -13121
rect 12927 -13239 13000 -13121
rect 9000 -13281 13000 -13239
rect 9000 -13399 9076 -13281
rect 9194 -13399 12809 -13281
rect 12927 -13399 13000 -13281
rect 9000 -13441 13000 -13399
rect 9000 -13559 9076 -13441
rect 9194 -13559 12809 -13441
rect 12927 -13559 13000 -13441
rect 9000 -13601 13000 -13559
rect 9000 -13719 9076 -13601
rect 9194 -13719 12809 -13601
rect 12927 -13719 13000 -13601
rect 9000 -13761 13000 -13719
rect 9000 -13879 9076 -13761
rect 9194 -13879 12809 -13761
rect 12927 -13879 13000 -13761
rect 9000 -13921 13000 -13879
rect 9000 -14039 9076 -13921
rect 9194 -14039 12809 -13921
rect 12927 -14039 13000 -13921
rect 9000 -14081 13000 -14039
rect 9000 -14199 9076 -14081
rect 9194 -14199 12809 -14081
rect 12927 -14199 13000 -14081
rect 9000 -14241 13000 -14199
rect 9000 -14359 9076 -14241
rect 9194 -14359 12809 -14241
rect 12927 -14359 13000 -14241
rect 9000 -14401 13000 -14359
rect 9000 -14519 9076 -14401
rect 9194 -14519 12809 -14401
rect 12927 -14519 13000 -14401
rect 9000 -14561 13000 -14519
rect 9000 -14679 9076 -14561
rect 9194 -14679 12809 -14561
rect 12927 -14679 13000 -14561
rect 9000 -14721 13000 -14679
rect 9000 -14839 9076 -14721
rect 9194 -14839 12809 -14721
rect 12927 -14839 13000 -14721
rect 9000 -14881 13000 -14839
rect 9000 -14999 9076 -14881
rect 9194 -14999 12809 -14881
rect 12927 -14999 13000 -14881
rect 9000 -15041 13000 -14999
rect 9000 -15159 9076 -15041
rect 9194 -15159 12809 -15041
rect 12927 -15159 13000 -15041
rect 9000 -15201 13000 -15159
rect 9000 -15319 9076 -15201
rect 9194 -15306 12809 -15201
rect 9194 -15319 9261 -15306
rect 9000 -15424 9261 -15319
rect 9379 -15424 9421 -15306
rect 9539 -15424 9581 -15306
rect 9699 -15424 9741 -15306
rect 9859 -15424 9901 -15306
rect 10019 -15424 10061 -15306
rect 10179 -15424 10221 -15306
rect 10339 -15424 10381 -15306
rect 10499 -15424 10541 -15306
rect 10659 -15424 10701 -15306
rect 10819 -15424 10861 -15306
rect 10979 -15424 11021 -15306
rect 11139 -15424 11181 -15306
rect 11299 -15424 11341 -15306
rect 11459 -15424 11501 -15306
rect 11619 -15424 11661 -15306
rect 11779 -15424 11821 -15306
rect 11939 -15424 11981 -15306
rect 12099 -15424 12141 -15306
rect 12259 -15424 12301 -15306
rect 12419 -15424 12461 -15306
rect 12579 -15424 12621 -15306
rect 12739 -15319 12809 -15306
rect 12927 -15319 13000 -15201
rect 12739 -15424 13000 -15319
rect 9000 -15500 13000 -15424
rect 15000 -11578 19000 -11500
rect 15000 -11681 15261 -11578
rect 15000 -11799 15076 -11681
rect 15194 -11696 15261 -11681
rect 15379 -11696 15421 -11578
rect 15539 -11696 15581 -11578
rect 15699 -11696 15741 -11578
rect 15859 -11696 15901 -11578
rect 16019 -11696 16061 -11578
rect 16179 -11696 16221 -11578
rect 16339 -11696 16381 -11578
rect 16499 -11696 16541 -11578
rect 16659 -11696 16701 -11578
rect 16819 -11696 16861 -11578
rect 16979 -11696 17021 -11578
rect 17139 -11696 17181 -11578
rect 17299 -11696 17341 -11578
rect 17459 -11696 17501 -11578
rect 17619 -11696 17661 -11578
rect 17779 -11696 17821 -11578
rect 17939 -11696 17981 -11578
rect 18099 -11696 18141 -11578
rect 18259 -11696 18301 -11578
rect 18419 -11696 18461 -11578
rect 18579 -11696 18621 -11578
rect 18739 -11681 19000 -11578
rect 18739 -11696 18809 -11681
rect 15194 -11799 18809 -11696
rect 18927 -11799 19000 -11681
rect 15000 -11841 19000 -11799
rect 15000 -11959 15076 -11841
rect 15194 -11959 18809 -11841
rect 18927 -11959 19000 -11841
rect 15000 -12001 19000 -11959
rect 15000 -12119 15076 -12001
rect 15194 -12119 18809 -12001
rect 18927 -12119 19000 -12001
rect 15000 -12161 19000 -12119
rect 15000 -12279 15076 -12161
rect 15194 -12279 18809 -12161
rect 18927 -12279 19000 -12161
rect 15000 -12321 19000 -12279
rect 15000 -12439 15076 -12321
rect 15194 -12439 18809 -12321
rect 18927 -12439 19000 -12321
rect 15000 -12481 19000 -12439
rect 15000 -12599 15076 -12481
rect 15194 -12599 18809 -12481
rect 18927 -12599 19000 -12481
rect 15000 -12641 19000 -12599
rect 15000 -12759 15076 -12641
rect 15194 -12759 18809 -12641
rect 18927 -12759 19000 -12641
rect 15000 -12801 19000 -12759
rect 15000 -12919 15076 -12801
rect 15194 -12919 18809 -12801
rect 18927 -12919 19000 -12801
rect 15000 -12961 19000 -12919
rect 15000 -13079 15076 -12961
rect 15194 -13079 18809 -12961
rect 18927 -13079 19000 -12961
rect 15000 -13121 19000 -13079
rect 15000 -13239 15076 -13121
rect 15194 -13239 18809 -13121
rect 18927 -13239 19000 -13121
rect 15000 -13281 19000 -13239
rect 15000 -13399 15076 -13281
rect 15194 -13399 18809 -13281
rect 18927 -13399 19000 -13281
rect 15000 -13441 19000 -13399
rect 15000 -13559 15076 -13441
rect 15194 -13559 18809 -13441
rect 18927 -13559 19000 -13441
rect 15000 -13601 19000 -13559
rect 15000 -13719 15076 -13601
rect 15194 -13719 18809 -13601
rect 18927 -13719 19000 -13601
rect 15000 -13761 19000 -13719
rect 15000 -13879 15076 -13761
rect 15194 -13879 18809 -13761
rect 18927 -13879 19000 -13761
rect 15000 -13921 19000 -13879
rect 15000 -14039 15076 -13921
rect 15194 -14039 18809 -13921
rect 18927 -14039 19000 -13921
rect 15000 -14081 19000 -14039
rect 15000 -14199 15076 -14081
rect 15194 -14199 18809 -14081
rect 18927 -14199 19000 -14081
rect 15000 -14241 19000 -14199
rect 15000 -14359 15076 -14241
rect 15194 -14359 18809 -14241
rect 18927 -14359 19000 -14241
rect 15000 -14401 19000 -14359
rect 15000 -14519 15076 -14401
rect 15194 -14519 18809 -14401
rect 18927 -14519 19000 -14401
rect 15000 -14561 19000 -14519
rect 15000 -14679 15076 -14561
rect 15194 -14679 18809 -14561
rect 18927 -14679 19000 -14561
rect 15000 -14721 19000 -14679
rect 15000 -14839 15076 -14721
rect 15194 -14839 18809 -14721
rect 18927 -14839 19000 -14721
rect 15000 -14881 19000 -14839
rect 15000 -14999 15076 -14881
rect 15194 -14999 18809 -14881
rect 18927 -14999 19000 -14881
rect 15000 -15041 19000 -14999
rect 15000 -15159 15076 -15041
rect 15194 -15159 18809 -15041
rect 18927 -15159 19000 -15041
rect 15000 -15201 19000 -15159
rect 15000 -15319 15076 -15201
rect 15194 -15306 18809 -15201
rect 15194 -15319 15261 -15306
rect 15000 -15424 15261 -15319
rect 15379 -15424 15421 -15306
rect 15539 -15424 15581 -15306
rect 15699 -15424 15741 -15306
rect 15859 -15424 15901 -15306
rect 16019 -15424 16061 -15306
rect 16179 -15424 16221 -15306
rect 16339 -15424 16381 -15306
rect 16499 -15424 16541 -15306
rect 16659 -15424 16701 -15306
rect 16819 -15424 16861 -15306
rect 16979 -15424 17021 -15306
rect 17139 -15424 17181 -15306
rect 17299 -15424 17341 -15306
rect 17459 -15424 17501 -15306
rect 17619 -15424 17661 -15306
rect 17779 -15424 17821 -15306
rect 17939 -15424 17981 -15306
rect 18099 -15424 18141 -15306
rect 18259 -15424 18301 -15306
rect 18419 -15424 18461 -15306
rect 18579 -15424 18621 -15306
rect 18739 -15319 18809 -15306
rect 18927 -15319 19000 -15201
rect 18739 -15424 19000 -15319
rect 15000 -15500 19000 -15424
rect 21000 -11578 25000 -11500
rect 21000 -11681 21261 -11578
rect 21000 -11799 21076 -11681
rect 21194 -11696 21261 -11681
rect 21379 -11696 21421 -11578
rect 21539 -11696 21581 -11578
rect 21699 -11696 21741 -11578
rect 21859 -11696 21901 -11578
rect 22019 -11696 22061 -11578
rect 22179 -11696 22221 -11578
rect 22339 -11696 22381 -11578
rect 22499 -11696 22541 -11578
rect 22659 -11696 22701 -11578
rect 22819 -11696 22861 -11578
rect 22979 -11696 23021 -11578
rect 23139 -11696 23181 -11578
rect 23299 -11696 23341 -11578
rect 23459 -11696 23501 -11578
rect 23619 -11696 23661 -11578
rect 23779 -11696 23821 -11578
rect 23939 -11696 23981 -11578
rect 24099 -11696 24141 -11578
rect 24259 -11696 24301 -11578
rect 24419 -11696 24461 -11578
rect 24579 -11696 24621 -11578
rect 24739 -11681 25000 -11578
rect 24739 -11696 24809 -11681
rect 21194 -11799 24809 -11696
rect 24927 -11799 25000 -11681
rect 21000 -11841 25000 -11799
rect 21000 -11959 21076 -11841
rect 21194 -11959 24809 -11841
rect 24927 -11959 25000 -11841
rect 21000 -12001 25000 -11959
rect 21000 -12119 21076 -12001
rect 21194 -12119 24809 -12001
rect 24927 -12119 25000 -12001
rect 21000 -12161 25000 -12119
rect 21000 -12279 21076 -12161
rect 21194 -12279 24809 -12161
rect 24927 -12279 25000 -12161
rect 21000 -12321 25000 -12279
rect 21000 -12439 21076 -12321
rect 21194 -12439 24809 -12321
rect 24927 -12439 25000 -12321
rect 21000 -12481 25000 -12439
rect 21000 -12599 21076 -12481
rect 21194 -12599 24809 -12481
rect 24927 -12599 25000 -12481
rect 21000 -12641 25000 -12599
rect 21000 -12759 21076 -12641
rect 21194 -12759 24809 -12641
rect 24927 -12759 25000 -12641
rect 21000 -12801 25000 -12759
rect 21000 -12919 21076 -12801
rect 21194 -12919 24809 -12801
rect 24927 -12919 25000 -12801
rect 21000 -12961 25000 -12919
rect 21000 -13079 21076 -12961
rect 21194 -13079 24809 -12961
rect 24927 -13079 25000 -12961
rect 21000 -13121 25000 -13079
rect 21000 -13239 21076 -13121
rect 21194 -13239 24809 -13121
rect 24927 -13239 25000 -13121
rect 21000 -13281 25000 -13239
rect 21000 -13399 21076 -13281
rect 21194 -13399 24809 -13281
rect 24927 -13399 25000 -13281
rect 21000 -13441 25000 -13399
rect 21000 -13559 21076 -13441
rect 21194 -13559 24809 -13441
rect 24927 -13559 25000 -13441
rect 21000 -13601 25000 -13559
rect 21000 -13719 21076 -13601
rect 21194 -13719 24809 -13601
rect 24927 -13719 25000 -13601
rect 21000 -13761 25000 -13719
rect 21000 -13879 21076 -13761
rect 21194 -13879 24809 -13761
rect 24927 -13879 25000 -13761
rect 21000 -13921 25000 -13879
rect 21000 -14039 21076 -13921
rect 21194 -14039 24809 -13921
rect 24927 -14039 25000 -13921
rect 21000 -14081 25000 -14039
rect 21000 -14199 21076 -14081
rect 21194 -14199 24809 -14081
rect 24927 -14199 25000 -14081
rect 21000 -14241 25000 -14199
rect 21000 -14359 21076 -14241
rect 21194 -14359 24809 -14241
rect 24927 -14359 25000 -14241
rect 21000 -14401 25000 -14359
rect 21000 -14519 21076 -14401
rect 21194 -14519 24809 -14401
rect 24927 -14519 25000 -14401
rect 21000 -14561 25000 -14519
rect 21000 -14679 21076 -14561
rect 21194 -14679 24809 -14561
rect 24927 -14679 25000 -14561
rect 21000 -14721 25000 -14679
rect 21000 -14839 21076 -14721
rect 21194 -14839 24809 -14721
rect 24927 -14839 25000 -14721
rect 21000 -14881 25000 -14839
rect 21000 -14999 21076 -14881
rect 21194 -14999 24809 -14881
rect 24927 -14999 25000 -14881
rect 21000 -15041 25000 -14999
rect 21000 -15159 21076 -15041
rect 21194 -15159 24809 -15041
rect 24927 -15159 25000 -15041
rect 21000 -15201 25000 -15159
rect 21000 -15319 21076 -15201
rect 21194 -15306 24809 -15201
rect 21194 -15319 21261 -15306
rect 21000 -15424 21261 -15319
rect 21379 -15424 21421 -15306
rect 21539 -15424 21581 -15306
rect 21699 -15424 21741 -15306
rect 21859 -15424 21901 -15306
rect 22019 -15424 22061 -15306
rect 22179 -15424 22221 -15306
rect 22339 -15424 22381 -15306
rect 22499 -15424 22541 -15306
rect 22659 -15424 22701 -15306
rect 22819 -15424 22861 -15306
rect 22979 -15424 23021 -15306
rect 23139 -15424 23181 -15306
rect 23299 -15424 23341 -15306
rect 23459 -15424 23501 -15306
rect 23619 -15424 23661 -15306
rect 23779 -15424 23821 -15306
rect 23939 -15424 23981 -15306
rect 24099 -15424 24141 -15306
rect 24259 -15424 24301 -15306
rect 24419 -15424 24461 -15306
rect 24579 -15424 24621 -15306
rect 24739 -15319 24809 -15306
rect 24927 -15319 25000 -15201
rect 24739 -15424 25000 -15319
rect 21000 -15500 25000 -15424
<< glass >>
rect 3300 5800 6700 9200
rect 9300 5800 12700 9200
rect 15300 5800 18700 9200
rect 21300 5800 24700 9200
rect 3300 -200 6700 3200
rect 9300 -200 12700 3200
rect 15300 -200 18700 3200
rect 21300 -200 24700 3200
rect 3300 -9200 6700 -5800
rect 9300 -9200 12700 -5800
rect 15300 -9200 18700 -5800
rect 21300 -9200 24700 -5800
rect 3300 -15200 6700 -11800
rect 9300 -15200 12700 -11800
rect 15300 -15200 18700 -11800
rect 21300 -15200 24700 -11800
<< fillblock >>
rect 3000 -10000 4200 -9500
rect 9000 -10000 10200 -9500
rect 15000 -10000 16200 -9500
rect 21000 -10000 22200 -9500
rect 3000 -11500 3400 -10900
rect 9000 -11500 9400 -10910
rect 15000 -11500 16600 -11000
rect 21000 -11500 22200 -11000
<< comment >>
rect 27000 -700 27100 3500
rect 900 -9500 1000 -5300
use cmota_gb_rp_gp  cmota_gb_rp_gp_0
timestamp 1672206111
transform 1 0 10100 0 1 -1250
box -3500 -3900 1401 300
use cmota_gp  cmota_gp_0
timestamp 1672297736
transform -1 0 17900 0 -1 -4750
box -3800 -3900 2150 350
use sky130hd_esd  sky130hd_esd_0
timestamp 1671850507
transform 0 1 19320 1 0 -883
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_1
timestamp 1671850507
transform -1 0 16552 0 -1 -2049
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_2
timestamp 1671850507
transform -1 0 16414 0 -1 -2049
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_3
timestamp 1671850507
transform 1 0 11586 0 1 -3951
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_4
timestamp 1671850507
transform 1 0 11448 0 1 -3951
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_5
timestamp 1671850507
transform 0 -1 8680 -1 0 -5117
box 111 -30 333 290
<< labels >>
rlabel metal5 3600 -8800 6250 -6500 1 VHI
rlabel metal5 9750 -8700 12400 -6400 1 VLO
rlabel metal5 15650 -8700 18300 -6400 1 VIP
rlabel metal5 21650 -8700 24300 -6400 1 VOP
rlabel metal5 21650 -14600 24300 -12300 1 VIN
rlabel metal5 15650 -14650 18300 -12350 1 VREF
rlabel metal5 9700 -14650 12350 -12350 1 SBAR
rlabel metal5 3750 -14700 6400 -12400 1 S
rlabel metal5 21750 500 24400 2800 5 VHI
rlabel metal5 15600 400 18250 2700 5 VLO
rlabel metal5 9700 400 12350 2700 5 VIP
rlabel metal5 3700 400 6350 2700 5 VOP
rlabel metal5 3700 6300 6350 8600 5 VIN
rlabel metal5 9700 6350 12350 8650 5 VREF
rlabel metal5 15650 6350 18300 8650 5 SBAR
rlabel metal5 21600 6400 24250 8700 5 S
<< end >>
