magic
tech sky130A
magscale 1 2
timestamp 1672031511
<< error_p >>
rect -19 46 55 51
rect -19 -10 -10 46
rect -19 -15 55 -10
<< metal2 >>
rect -19 -10 -10 46
rect 46 -10 55 46
<< via2 >>
rect -10 -10 46 46
<< metal3 >>
rect -19 46 55 51
rect -19 -10 -10 46
rect 46 -10 55 46
rect -19 -15 55 -10
<< end >>
