magic
tech sky130B
timestamp 1668124831
<< metal4 >>
rect 280 5240 1080 5260
rect 280 -140 300 5240
rect 420 5030 940 5240
rect 420 -140 510 5030
rect 280 -160 510 -140
rect 540 4920 820 5000
rect 540 -140 620 4920
rect 740 -140 820 4920
rect 540 -160 820 -140
rect 850 -140 940 5030
rect 1060 -140 1080 5240
rect 850 -160 1080 -140
rect 1860 4420 2140 4520
rect 1860 -160 1920 4420
rect 1950 -160 2050 4390
rect 2080 -160 2140 4420
<< via4 >>
rect 300 -140 420 5240
rect 620 -140 740 4920
rect 940 -140 1060 5240
<< metal5 >>
rect 280 5240 1080 5260
rect 280 -140 300 5240
rect 420 5100 940 5240
rect 420 -140 440 5100
rect 280 -160 440 -140
rect 600 4920 760 4940
rect 600 -140 620 4920
rect 740 -140 760 4920
rect 600 -160 760 -140
rect 920 -140 940 5100
rect 1060 -140 1080 5240
rect 920 -160 1080 -140
<< labels >>
rlabel space 460 -160 760 0 1 B
rlabel space 480 5240 780 5400 1 A
rlabel metal5 600 -160 760 0 1 TOP
rlabel metal5 610 5100 770 5260 1 BOT
rlabel metal4 1950 -160 2050 -100 1 TOP2
rlabel metal4 1920 4420 2080 4520 1 BOT2
<< end >>
