magic
tech sky130A
magscale 1 2
timestamp 1671406405
use cmota_gp  cmota_gp_0
timestamp 1671336542
transform 1 0 11534 0 -1 -8102
box -7600 -7800 2527 600
use cmota_gp  cmota_gp_2
timestamp 1671336542
transform 1 0 11610 0 1 13366
box -7600 -7800 2527 600
use isrc  isrc_0
timestamp 1671401643
transform 1 0 10508 0 1 -1702
box -200 1760 4090 5700
use swcap_array_1  swcap_array_1_0
timestamp 1671395052
transform 0 -1 37998 1 0 -171
box -6569 -1080 7773 23570
use twcon_flat  twcon_flat_0
timestamp 1671388962
transform 1 0 5307 0 1 1620
box -5309 -1622 4974 3682
<< end >>
