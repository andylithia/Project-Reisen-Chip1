magic
tech sky130A
magscale 1 2
timestamp 1671169778
<< nwell >>
rect -163 66 5363 2504
<< pwell >>
rect -164 -2434 1350 -14
rect 1473 -1110 3727 -190
rect 1517 -3550 3683 -1130
rect 3849 -2434 5363 -14
<< nmos >>
rect 32 -2224 92 -224
rect 150 -2224 210 -224
rect 268 -2224 328 -224
rect 386 -2224 446 -224
rect 504 -2224 564 -224
rect 622 -2224 682 -224
rect 740 -2224 800 -224
rect 858 -2224 918 -224
rect 976 -2224 1036 -224
rect 1094 -2224 1154 -224
rect 1713 -3340 2113 -1340
rect 2171 -3340 2571 -1340
rect 2629 -3340 3029 -1340
rect 3087 -3340 3487 -1340
rect 4045 -2224 4105 -224
rect 4163 -2224 4223 -224
rect 4281 -2224 4341 -224
rect 4399 -2224 4459 -224
rect 4517 -2224 4577 -224
rect 4635 -2224 4695 -224
rect 4753 -2224 4813 -224
rect 4871 -2224 4931 -224
rect 4989 -2224 5049 -224
rect 5107 -2224 5167 -224
<< pmos >>
rect 33 285 93 2285
rect 151 285 211 2285
rect 269 285 329 2285
rect 387 285 447 2285
rect 505 285 565 2285
rect 623 285 683 2285
rect 741 285 801 2285
rect 859 285 919 2285
rect 977 285 1037 2285
rect 1095 285 1155 2285
rect 1213 285 1273 2285
rect 1331 285 1391 2285
rect 1449 285 1509 2285
rect 1567 285 1627 2285
rect 1685 285 1745 2285
rect 1803 285 1863 2285
rect 1921 285 1981 2285
rect 2039 285 2099 2285
rect 2157 285 2217 2285
rect 2275 285 2335 2285
rect 2393 285 2453 2285
rect 2511 285 2571 2285
rect 2629 285 2689 2285
rect 2747 285 2807 2285
rect 2865 285 2925 2285
rect 2983 285 3043 2285
rect 3101 285 3161 2285
rect 3219 285 3279 2285
rect 3337 285 3397 2285
rect 3455 285 3515 2285
rect 3573 285 3633 2285
rect 3691 285 3751 2285
rect 3809 285 3869 2285
rect 3927 285 3987 2285
rect 4045 285 4105 2285
rect 4163 285 4223 2285
rect 4281 285 4341 2285
rect 4399 285 4459 2285
rect 4517 285 4577 2285
rect 4635 285 4695 2285
rect 4753 285 4813 2285
rect 4871 285 4931 2285
rect 4989 285 5049 2285
rect 5107 285 5167 2285
<< nmoslvt >>
rect 1673 -900 1703 -400
rect 1769 -900 1799 -400
rect 1865 -900 1895 -400
rect 1961 -900 1991 -400
rect 2057 -900 2087 -400
rect 2153 -900 2183 -400
rect 2249 -900 2279 -400
rect 2345 -900 2375 -400
rect 2441 -900 2471 -400
rect 2537 -900 2567 -400
rect 2633 -900 2663 -400
rect 2729 -900 2759 -400
rect 2825 -900 2855 -400
rect 2921 -900 2951 -400
rect 3017 -900 3047 -400
rect 3113 -900 3143 -400
rect 3209 -900 3239 -400
rect 3305 -900 3335 -400
rect 3401 -900 3431 -400
rect 3497 -900 3527 -400
<< ndiff >>
rect -26 -236 32 -224
rect -26 -2212 -14 -236
rect 20 -2212 32 -236
rect -26 -2224 32 -2212
rect 92 -236 150 -224
rect 92 -2212 104 -236
rect 138 -2212 150 -236
rect 92 -2224 150 -2212
rect 210 -236 268 -224
rect 210 -2212 222 -236
rect 256 -2212 268 -236
rect 210 -2224 268 -2212
rect 328 -236 386 -224
rect 328 -2212 340 -236
rect 374 -2212 386 -236
rect 328 -2224 386 -2212
rect 446 -236 504 -224
rect 446 -2212 458 -236
rect 492 -2212 504 -236
rect 446 -2224 504 -2212
rect 564 -236 622 -224
rect 564 -2212 576 -236
rect 610 -2212 622 -236
rect 564 -2224 622 -2212
rect 682 -236 740 -224
rect 682 -2212 694 -236
rect 728 -2212 740 -236
rect 682 -2224 740 -2212
rect 800 -236 858 -224
rect 800 -2212 812 -236
rect 846 -2212 858 -236
rect 800 -2224 858 -2212
rect 918 -236 976 -224
rect 918 -2212 930 -236
rect 964 -2212 976 -236
rect 918 -2224 976 -2212
rect 1036 -236 1094 -224
rect 1036 -2212 1048 -236
rect 1082 -2212 1094 -236
rect 1036 -2224 1094 -2212
rect 1154 -236 1212 -224
rect 1154 -2212 1166 -236
rect 1200 -2212 1212 -236
rect 1154 -2224 1212 -2212
rect 1611 -412 1673 -400
rect 1611 -888 1623 -412
rect 1657 -888 1673 -412
rect 1611 -900 1673 -888
rect 1703 -412 1769 -400
rect 1703 -888 1719 -412
rect 1753 -888 1769 -412
rect 1703 -900 1769 -888
rect 1799 -412 1865 -400
rect 1799 -888 1815 -412
rect 1849 -888 1865 -412
rect 1799 -900 1865 -888
rect 1895 -412 1961 -400
rect 1895 -888 1911 -412
rect 1945 -888 1961 -412
rect 1895 -900 1961 -888
rect 1991 -412 2057 -400
rect 1991 -888 2007 -412
rect 2041 -888 2057 -412
rect 1991 -900 2057 -888
rect 2087 -412 2153 -400
rect 2087 -888 2103 -412
rect 2137 -888 2153 -412
rect 2087 -900 2153 -888
rect 2183 -412 2249 -400
rect 2183 -888 2199 -412
rect 2233 -888 2249 -412
rect 2183 -900 2249 -888
rect 2279 -412 2345 -400
rect 2279 -888 2295 -412
rect 2329 -888 2345 -412
rect 2279 -900 2345 -888
rect 2375 -412 2441 -400
rect 2375 -888 2391 -412
rect 2425 -888 2441 -412
rect 2375 -900 2441 -888
rect 2471 -412 2537 -400
rect 2471 -888 2487 -412
rect 2521 -888 2537 -412
rect 2471 -900 2537 -888
rect 2567 -412 2633 -400
rect 2567 -888 2583 -412
rect 2617 -888 2633 -412
rect 2567 -900 2633 -888
rect 2663 -412 2729 -400
rect 2663 -888 2679 -412
rect 2713 -888 2729 -412
rect 2663 -900 2729 -888
rect 2759 -412 2825 -400
rect 2759 -888 2775 -412
rect 2809 -888 2825 -412
rect 2759 -900 2825 -888
rect 2855 -412 2921 -400
rect 2855 -888 2871 -412
rect 2905 -888 2921 -412
rect 2855 -900 2921 -888
rect 2951 -412 3017 -400
rect 2951 -888 2967 -412
rect 3001 -888 3017 -412
rect 2951 -900 3017 -888
rect 3047 -412 3113 -400
rect 3047 -888 3063 -412
rect 3097 -888 3113 -412
rect 3047 -900 3113 -888
rect 3143 -412 3209 -400
rect 3143 -888 3159 -412
rect 3193 -888 3209 -412
rect 3143 -900 3209 -888
rect 3239 -412 3305 -400
rect 3239 -888 3255 -412
rect 3289 -888 3305 -412
rect 3239 -900 3305 -888
rect 3335 -412 3401 -400
rect 3335 -888 3351 -412
rect 3385 -888 3401 -412
rect 3335 -900 3401 -888
rect 3431 -412 3497 -400
rect 3431 -888 3447 -412
rect 3481 -888 3497 -412
rect 3431 -900 3497 -888
rect 3527 -412 3589 -400
rect 3527 -888 3543 -412
rect 3577 -888 3589 -412
rect 3527 -900 3589 -888
rect 1655 -1352 1713 -1340
rect 1655 -3328 1667 -1352
rect 1701 -3328 1713 -1352
rect 1655 -3340 1713 -3328
rect 2113 -1352 2171 -1340
rect 2113 -3328 2125 -1352
rect 2159 -3328 2171 -1352
rect 2113 -3340 2171 -3328
rect 2571 -1352 2629 -1340
rect 2571 -3328 2583 -1352
rect 2617 -3328 2629 -1352
rect 2571 -3340 2629 -3328
rect 3029 -1352 3087 -1340
rect 3029 -3328 3041 -1352
rect 3075 -3328 3087 -1352
rect 3029 -3340 3087 -3328
rect 3487 -1352 3545 -1340
rect 3487 -3328 3499 -1352
rect 3533 -3328 3545 -1352
rect 3487 -3340 3545 -3328
rect 3987 -236 4045 -224
rect 3987 -2212 3999 -236
rect 4033 -2212 4045 -236
rect 3987 -2224 4045 -2212
rect 4105 -236 4163 -224
rect 4105 -2212 4117 -236
rect 4151 -2212 4163 -236
rect 4105 -2224 4163 -2212
rect 4223 -236 4281 -224
rect 4223 -2212 4235 -236
rect 4269 -2212 4281 -236
rect 4223 -2224 4281 -2212
rect 4341 -236 4399 -224
rect 4341 -2212 4353 -236
rect 4387 -2212 4399 -236
rect 4341 -2224 4399 -2212
rect 4459 -236 4517 -224
rect 4459 -2212 4471 -236
rect 4505 -2212 4517 -236
rect 4459 -2224 4517 -2212
rect 4577 -236 4635 -224
rect 4577 -2212 4589 -236
rect 4623 -2212 4635 -236
rect 4577 -2224 4635 -2212
rect 4695 -236 4753 -224
rect 4695 -2212 4707 -236
rect 4741 -2212 4753 -236
rect 4695 -2224 4753 -2212
rect 4813 -236 4871 -224
rect 4813 -2212 4825 -236
rect 4859 -2212 4871 -236
rect 4813 -2224 4871 -2212
rect 4931 -236 4989 -224
rect 4931 -2212 4943 -236
rect 4977 -2212 4989 -236
rect 4931 -2224 4989 -2212
rect 5049 -236 5107 -224
rect 5049 -2212 5061 -236
rect 5095 -2212 5107 -236
rect 5049 -2224 5107 -2212
rect 5167 -236 5225 -224
rect 5167 -2212 5179 -236
rect 5213 -2212 5225 -236
rect 5167 -2224 5225 -2212
<< pdiff >>
rect -25 2273 33 2285
rect -25 297 -13 2273
rect 21 297 33 2273
rect -25 285 33 297
rect 93 2273 151 2285
rect 93 297 105 2273
rect 139 297 151 2273
rect 93 285 151 297
rect 211 2273 269 2285
rect 211 297 223 2273
rect 257 297 269 2273
rect 211 285 269 297
rect 329 2273 387 2285
rect 329 297 341 2273
rect 375 297 387 2273
rect 329 285 387 297
rect 447 2273 505 2285
rect 447 297 459 2273
rect 493 297 505 2273
rect 447 285 505 297
rect 565 2273 623 2285
rect 565 297 577 2273
rect 611 297 623 2273
rect 565 285 623 297
rect 683 2273 741 2285
rect 683 297 695 2273
rect 729 297 741 2273
rect 683 285 741 297
rect 801 2273 859 2285
rect 801 297 813 2273
rect 847 297 859 2273
rect 801 285 859 297
rect 919 2273 977 2285
rect 919 297 931 2273
rect 965 297 977 2273
rect 919 285 977 297
rect 1037 2273 1095 2285
rect 1037 297 1049 2273
rect 1083 297 1095 2273
rect 1037 285 1095 297
rect 1155 2273 1213 2285
rect 1155 297 1167 2273
rect 1201 297 1213 2273
rect 1155 285 1213 297
rect 1273 2273 1331 2285
rect 1273 297 1285 2273
rect 1319 297 1331 2273
rect 1273 285 1331 297
rect 1391 2273 1449 2285
rect 1391 297 1403 2273
rect 1437 297 1449 2273
rect 1391 285 1449 297
rect 1509 2273 1567 2285
rect 1509 297 1521 2273
rect 1555 297 1567 2273
rect 1509 285 1567 297
rect 1627 2273 1685 2285
rect 1627 297 1639 2273
rect 1673 297 1685 2273
rect 1627 285 1685 297
rect 1745 2273 1803 2285
rect 1745 297 1757 2273
rect 1791 297 1803 2273
rect 1745 285 1803 297
rect 1863 2273 1921 2285
rect 1863 297 1875 2273
rect 1909 297 1921 2273
rect 1863 285 1921 297
rect 1981 2273 2039 2285
rect 1981 297 1993 2273
rect 2027 297 2039 2273
rect 1981 285 2039 297
rect 2099 2273 2157 2285
rect 2099 297 2111 2273
rect 2145 297 2157 2273
rect 2099 285 2157 297
rect 2217 2273 2275 2285
rect 2217 297 2229 2273
rect 2263 297 2275 2273
rect 2217 285 2275 297
rect 2335 2273 2393 2285
rect 2335 297 2347 2273
rect 2381 297 2393 2273
rect 2335 285 2393 297
rect 2453 2273 2511 2285
rect 2453 297 2465 2273
rect 2499 297 2511 2273
rect 2453 285 2511 297
rect 2571 2273 2629 2285
rect 2571 297 2583 2273
rect 2617 297 2629 2273
rect 2571 285 2629 297
rect 2689 2273 2747 2285
rect 2689 297 2701 2273
rect 2735 297 2747 2273
rect 2689 285 2747 297
rect 2807 2273 2865 2285
rect 2807 297 2819 2273
rect 2853 297 2865 2273
rect 2807 285 2865 297
rect 2925 2273 2983 2285
rect 2925 297 2937 2273
rect 2971 297 2983 2273
rect 2925 285 2983 297
rect 3043 2273 3101 2285
rect 3043 297 3055 2273
rect 3089 297 3101 2273
rect 3043 285 3101 297
rect 3161 2273 3219 2285
rect 3161 297 3173 2273
rect 3207 297 3219 2273
rect 3161 285 3219 297
rect 3279 2273 3337 2285
rect 3279 297 3291 2273
rect 3325 297 3337 2273
rect 3279 285 3337 297
rect 3397 2273 3455 2285
rect 3397 297 3409 2273
rect 3443 297 3455 2273
rect 3397 285 3455 297
rect 3515 2273 3573 2285
rect 3515 297 3527 2273
rect 3561 297 3573 2273
rect 3515 285 3573 297
rect 3633 2273 3691 2285
rect 3633 297 3645 2273
rect 3679 297 3691 2273
rect 3633 285 3691 297
rect 3751 2273 3809 2285
rect 3751 297 3763 2273
rect 3797 297 3809 2273
rect 3751 285 3809 297
rect 3869 2273 3927 2285
rect 3869 297 3881 2273
rect 3915 297 3927 2273
rect 3869 285 3927 297
rect 3987 2273 4045 2285
rect 3987 297 3999 2273
rect 4033 297 4045 2273
rect 3987 285 4045 297
rect 4105 2273 4163 2285
rect 4105 297 4117 2273
rect 4151 297 4163 2273
rect 4105 285 4163 297
rect 4223 2273 4281 2285
rect 4223 297 4235 2273
rect 4269 297 4281 2273
rect 4223 285 4281 297
rect 4341 2273 4399 2285
rect 4341 297 4353 2273
rect 4387 297 4399 2273
rect 4341 285 4399 297
rect 4459 2273 4517 2285
rect 4459 297 4471 2273
rect 4505 297 4517 2273
rect 4459 285 4517 297
rect 4577 2273 4635 2285
rect 4577 297 4589 2273
rect 4623 297 4635 2273
rect 4577 285 4635 297
rect 4695 2273 4753 2285
rect 4695 297 4707 2273
rect 4741 297 4753 2273
rect 4695 285 4753 297
rect 4813 2273 4871 2285
rect 4813 297 4825 2273
rect 4859 297 4871 2273
rect 4813 285 4871 297
rect 4931 2273 4989 2285
rect 4931 297 4943 2273
rect 4977 297 4989 2273
rect 4931 285 4989 297
rect 5049 2273 5107 2285
rect 5049 297 5061 2273
rect 5095 297 5107 2273
rect 5049 285 5107 297
rect 5167 2273 5225 2285
rect 5167 297 5179 2273
rect 5213 297 5225 2273
rect 5167 285 5225 297
<< ndiffc >>
rect -14 -2212 20 -236
rect 104 -2212 138 -236
rect 222 -2212 256 -236
rect 340 -2212 374 -236
rect 458 -2212 492 -236
rect 576 -2212 610 -236
rect 694 -2212 728 -236
rect 812 -2212 846 -236
rect 930 -2212 964 -236
rect 1048 -2212 1082 -236
rect 1166 -2212 1200 -236
rect 1623 -888 1657 -412
rect 1719 -888 1753 -412
rect 1815 -888 1849 -412
rect 1911 -888 1945 -412
rect 2007 -888 2041 -412
rect 2103 -888 2137 -412
rect 2199 -888 2233 -412
rect 2295 -888 2329 -412
rect 2391 -888 2425 -412
rect 2487 -888 2521 -412
rect 2583 -888 2617 -412
rect 2679 -888 2713 -412
rect 2775 -888 2809 -412
rect 2871 -888 2905 -412
rect 2967 -888 3001 -412
rect 3063 -888 3097 -412
rect 3159 -888 3193 -412
rect 3255 -888 3289 -412
rect 3351 -888 3385 -412
rect 3447 -888 3481 -412
rect 3543 -888 3577 -412
rect 1667 -3328 1701 -1352
rect 2125 -3328 2159 -1352
rect 2583 -3328 2617 -1352
rect 3041 -3328 3075 -1352
rect 3499 -3328 3533 -1352
rect 3999 -2212 4033 -236
rect 4117 -2212 4151 -236
rect 4235 -2212 4269 -236
rect 4353 -2212 4387 -236
rect 4471 -2212 4505 -236
rect 4589 -2212 4623 -236
rect 4707 -2212 4741 -236
rect 4825 -2212 4859 -236
rect 4943 -2212 4977 -236
rect 5061 -2212 5095 -236
rect 5179 -2212 5213 -236
<< pdiffc >>
rect -13 297 21 2273
rect 105 297 139 2273
rect 223 297 257 2273
rect 341 297 375 2273
rect 459 297 493 2273
rect 577 297 611 2273
rect 695 297 729 2273
rect 813 297 847 2273
rect 931 297 965 2273
rect 1049 297 1083 2273
rect 1167 297 1201 2273
rect 1285 297 1319 2273
rect 1403 297 1437 2273
rect 1521 297 1555 2273
rect 1639 297 1673 2273
rect 1757 297 1791 2273
rect 1875 297 1909 2273
rect 1993 297 2027 2273
rect 2111 297 2145 2273
rect 2229 297 2263 2273
rect 2347 297 2381 2273
rect 2465 297 2499 2273
rect 2583 297 2617 2273
rect 2701 297 2735 2273
rect 2819 297 2853 2273
rect 2937 297 2971 2273
rect 3055 297 3089 2273
rect 3173 297 3207 2273
rect 3291 297 3325 2273
rect 3409 297 3443 2273
rect 3527 297 3561 2273
rect 3645 297 3679 2273
rect 3763 297 3797 2273
rect 3881 297 3915 2273
rect 3999 297 4033 2273
rect 4117 297 4151 2273
rect 4235 297 4269 2273
rect 4353 297 4387 2273
rect 4471 297 4505 2273
rect 4589 297 4623 2273
rect 4707 297 4741 2273
rect 4825 297 4859 2273
rect 4943 297 4977 2273
rect 5061 297 5095 2273
rect 5179 297 5213 2273
<< psubdiff >>
rect -128 -84 -32 -50
rect 1218 -84 1314 -50
rect -128 -146 -94 -84
rect 1280 -146 1314 -84
rect -128 -2364 -94 -2302
rect 3885 -84 3981 -50
rect 5231 -84 5327 -50
rect 3885 -146 3919 -84
rect 1509 -260 1605 -226
rect 3595 -260 3691 -226
rect 1509 -322 1543 -260
rect 3657 -322 3691 -260
rect 1509 -1040 1543 -978
rect 3657 -1040 3691 -978
rect 1509 -1074 1605 -1040
rect 3595 -1074 3691 -1040
rect 1280 -2364 1314 -2302
rect -128 -2398 -32 -2364
rect 1218 -2398 1314 -2364
rect 1553 -1200 1649 -1166
rect 3551 -1200 3647 -1166
rect 1553 -1262 1587 -1200
rect 3613 -1262 3647 -1200
rect 1553 -3480 1587 -3418
rect 5293 -146 5327 -84
rect 3885 -2364 3919 -2302
rect 5293 -2364 5327 -2302
rect 3885 -2398 3981 -2364
rect 5231 -2398 5327 -2364
rect 3613 -3480 3647 -3418
rect 1553 -3514 1649 -3480
rect 3551 -3514 3647 -3480
<< nsubdiff >>
rect -127 2434 -31 2468
rect 5231 2434 5327 2468
rect -127 2372 -93 2434
rect 5293 2372 5327 2434
rect -127 136 -93 198
rect 5293 136 5327 198
rect -127 102 -31 136
rect 5231 102 5327 136
<< psubdiffcont >>
rect -32 -84 1218 -50
rect -128 -2302 -94 -146
rect 1280 -2302 1314 -146
rect 3981 -84 5231 -50
rect 1605 -260 3595 -226
rect 1509 -978 1543 -322
rect 3657 -978 3691 -322
rect 1605 -1074 3595 -1040
rect -32 -2398 1218 -2364
rect 1649 -1200 3551 -1166
rect 1553 -3418 1587 -1262
rect 3613 -3418 3647 -1262
rect 3885 -2302 3919 -146
rect 5293 -2302 5327 -146
rect 3981 -2398 5231 -2364
rect 1649 -3514 3551 -3480
<< nsubdiffcont >>
rect -31 2434 5231 2468
rect -127 198 -93 2372
rect 5293 198 5327 2372
rect -31 102 5231 136
<< poly >>
rect 30 2366 96 2382
rect 30 2332 46 2366
rect 80 2332 96 2366
rect 30 2316 96 2332
rect 148 2366 214 2382
rect 148 2332 164 2366
rect 198 2332 214 2366
rect 148 2316 214 2332
rect 266 2366 332 2382
rect 266 2332 282 2366
rect 316 2332 332 2366
rect 266 2316 332 2332
rect 384 2366 450 2382
rect 384 2332 400 2366
rect 434 2332 450 2366
rect 384 2316 450 2332
rect 502 2366 568 2382
rect 502 2332 518 2366
rect 552 2332 568 2366
rect 502 2316 568 2332
rect 620 2366 686 2382
rect 620 2332 636 2366
rect 670 2332 686 2366
rect 620 2316 686 2332
rect 738 2366 804 2382
rect 738 2332 754 2366
rect 788 2332 804 2366
rect 738 2316 804 2332
rect 856 2366 922 2382
rect 856 2332 872 2366
rect 906 2332 922 2366
rect 856 2316 922 2332
rect 974 2366 1040 2382
rect 974 2332 990 2366
rect 1024 2332 1040 2366
rect 974 2316 1040 2332
rect 1092 2366 1158 2382
rect 1092 2332 1108 2366
rect 1142 2332 1158 2366
rect 1092 2316 1158 2332
rect 1210 2366 1276 2382
rect 1210 2332 1226 2366
rect 1260 2332 1276 2366
rect 1210 2316 1276 2332
rect 1328 2366 1394 2382
rect 1328 2332 1344 2366
rect 1378 2332 1394 2366
rect 1328 2316 1394 2332
rect 1446 2366 1512 2382
rect 1446 2332 1462 2366
rect 1496 2332 1512 2366
rect 1446 2316 1512 2332
rect 1564 2366 1630 2382
rect 1564 2332 1580 2366
rect 1614 2332 1630 2366
rect 1564 2316 1630 2332
rect 1682 2366 1748 2382
rect 1682 2332 1698 2366
rect 1732 2332 1748 2366
rect 1682 2316 1748 2332
rect 1800 2366 1866 2382
rect 1800 2332 1816 2366
rect 1850 2332 1866 2366
rect 1800 2316 1866 2332
rect 1918 2366 1984 2382
rect 1918 2332 1934 2366
rect 1968 2332 1984 2366
rect 1918 2316 1984 2332
rect 2036 2366 2102 2382
rect 2036 2332 2052 2366
rect 2086 2332 2102 2366
rect 2036 2316 2102 2332
rect 2154 2366 2220 2382
rect 2154 2332 2170 2366
rect 2204 2332 2220 2366
rect 2154 2316 2220 2332
rect 2272 2366 2338 2382
rect 2272 2332 2288 2366
rect 2322 2332 2338 2366
rect 2272 2316 2338 2332
rect 2390 2316 2456 2382
rect 2508 2316 2574 2382
rect 2626 2316 2692 2382
rect 2744 2316 2810 2382
rect 2862 2366 2928 2382
rect 2862 2332 2878 2366
rect 2912 2332 2928 2366
rect 2862 2316 2928 2332
rect 2980 2366 3046 2382
rect 2980 2332 2996 2366
rect 3030 2332 3046 2366
rect 2980 2316 3046 2332
rect 3098 2366 3164 2382
rect 3098 2332 3114 2366
rect 3148 2332 3164 2366
rect 3098 2316 3164 2332
rect 3216 2366 3282 2382
rect 3216 2332 3232 2366
rect 3266 2332 3282 2366
rect 3216 2316 3282 2332
rect 3334 2366 3400 2382
rect 3334 2332 3350 2366
rect 3384 2332 3400 2366
rect 3334 2316 3400 2332
rect 3452 2366 3518 2382
rect 3452 2332 3468 2366
rect 3502 2332 3518 2366
rect 3452 2316 3518 2332
rect 3570 2366 3636 2382
rect 3570 2332 3586 2366
rect 3620 2332 3636 2366
rect 3570 2316 3636 2332
rect 3688 2366 3754 2382
rect 3688 2332 3704 2366
rect 3738 2332 3754 2366
rect 3688 2316 3754 2332
rect 3806 2366 3872 2382
rect 3806 2332 3822 2366
rect 3856 2332 3872 2366
rect 3806 2316 3872 2332
rect 3924 2366 3990 2382
rect 3924 2332 3940 2366
rect 3974 2332 3990 2366
rect 3924 2316 3990 2332
rect 4042 2366 4108 2382
rect 4042 2332 4058 2366
rect 4092 2332 4108 2366
rect 4042 2316 4108 2332
rect 4160 2366 4226 2382
rect 4160 2332 4176 2366
rect 4210 2332 4226 2366
rect 4160 2316 4226 2332
rect 4278 2366 4344 2382
rect 4278 2332 4294 2366
rect 4328 2332 4344 2366
rect 4278 2316 4344 2332
rect 4396 2366 4462 2382
rect 4396 2332 4412 2366
rect 4446 2332 4462 2366
rect 4396 2316 4462 2332
rect 4514 2366 4580 2382
rect 4514 2332 4530 2366
rect 4564 2332 4580 2366
rect 4514 2316 4580 2332
rect 4632 2366 4698 2382
rect 4632 2332 4648 2366
rect 4682 2332 4698 2366
rect 4632 2316 4698 2332
rect 4750 2366 4816 2382
rect 4750 2332 4766 2366
rect 4800 2332 4816 2366
rect 4750 2316 4816 2332
rect 4868 2366 4934 2382
rect 4868 2332 4884 2366
rect 4918 2332 4934 2366
rect 4868 2316 4934 2332
rect 4986 2366 5052 2382
rect 4986 2332 5002 2366
rect 5036 2332 5052 2366
rect 4986 2316 5052 2332
rect 5104 2366 5170 2382
rect 5104 2332 5120 2366
rect 5154 2332 5170 2366
rect 5104 2316 5170 2332
rect 33 2285 93 2316
rect 151 2285 211 2316
rect 269 2285 329 2316
rect 387 2285 447 2316
rect 505 2285 565 2316
rect 623 2285 683 2316
rect 741 2285 801 2316
rect 859 2285 919 2316
rect 977 2285 1037 2316
rect 1095 2285 1155 2316
rect 1213 2285 1273 2316
rect 1331 2285 1391 2316
rect 1449 2285 1509 2316
rect 1567 2285 1627 2316
rect 1685 2285 1745 2316
rect 1803 2285 1863 2316
rect 1921 2285 1981 2316
rect 2039 2285 2099 2316
rect 2157 2285 2217 2316
rect 2275 2285 2335 2316
rect 2393 2285 2453 2316
rect 2511 2285 2571 2316
rect 2629 2285 2689 2316
rect 2747 2285 2807 2316
rect 2865 2285 2925 2316
rect 2983 2285 3043 2316
rect 3101 2285 3161 2316
rect 3219 2285 3279 2316
rect 3337 2285 3397 2316
rect 3455 2285 3515 2316
rect 3573 2285 3633 2316
rect 3691 2285 3751 2316
rect 3809 2285 3869 2316
rect 3927 2285 3987 2316
rect 4045 2285 4105 2316
rect 4163 2285 4223 2316
rect 4281 2285 4341 2316
rect 4399 2285 4459 2316
rect 4517 2285 4577 2316
rect 4635 2285 4695 2316
rect 4753 2285 4813 2316
rect 4871 2285 4931 2316
rect 4989 2285 5049 2316
rect 5107 2285 5167 2316
rect 33 254 93 285
rect 151 254 211 285
rect 269 254 329 285
rect 387 254 447 285
rect 505 254 565 285
rect 623 254 683 285
rect 741 254 801 285
rect 859 254 919 285
rect 977 254 1037 285
rect 1095 254 1155 285
rect 1213 254 1273 285
rect 1331 254 1391 285
rect 1449 254 1509 285
rect 1567 254 1627 285
rect 1685 254 1745 285
rect 1803 254 1863 285
rect 1921 254 1981 285
rect 2039 254 2099 285
rect 2157 254 2217 285
rect 2275 254 2335 285
rect 2393 254 2453 285
rect 2511 254 2571 285
rect 2629 254 2689 285
rect 2747 254 2807 285
rect 2865 254 2925 285
rect 2983 254 3043 285
rect 3101 254 3161 285
rect 3219 254 3279 285
rect 3337 254 3397 285
rect 3455 254 3515 285
rect 3573 254 3633 285
rect 3691 254 3751 285
rect 3809 254 3869 285
rect 3927 254 3987 285
rect 4045 254 4105 285
rect 4163 254 4223 285
rect 4281 254 4341 285
rect 4399 254 4459 285
rect 4517 254 4577 285
rect 4635 254 4695 285
rect 4753 254 4813 285
rect 4871 254 4931 285
rect 4989 254 5049 285
rect 5107 254 5167 285
rect 30 238 96 254
rect 30 204 46 238
rect 80 204 96 238
rect 30 188 96 204
rect 148 238 214 254
rect 148 204 164 238
rect 198 204 214 238
rect 148 188 214 204
rect 266 238 332 254
rect 266 204 282 238
rect 316 204 332 238
rect 266 188 332 204
rect 384 238 450 254
rect 384 204 400 238
rect 434 204 450 238
rect 384 188 450 204
rect 502 238 568 254
rect 502 204 518 238
rect 552 204 568 238
rect 502 188 568 204
rect 620 238 686 254
rect 620 204 636 238
rect 670 204 686 238
rect 620 188 686 204
rect 738 238 804 254
rect 738 204 754 238
rect 788 204 804 238
rect 738 188 804 204
rect 856 238 922 254
rect 856 204 872 238
rect 906 204 922 238
rect 856 188 922 204
rect 974 238 1040 254
rect 974 204 990 238
rect 1024 204 1040 238
rect 974 188 1040 204
rect 1092 238 1158 254
rect 1092 204 1108 238
rect 1142 204 1158 238
rect 1092 188 1158 204
rect 1210 238 1276 254
rect 1210 204 1226 238
rect 1260 204 1276 238
rect 1210 188 1276 204
rect 1328 238 1394 254
rect 1328 204 1344 238
rect 1378 204 1394 238
rect 1328 188 1394 204
rect 1446 238 1512 254
rect 1446 204 1462 238
rect 1496 204 1512 238
rect 1446 188 1512 204
rect 1564 238 1630 254
rect 1564 204 1580 238
rect 1614 204 1630 238
rect 1564 188 1630 204
rect 1682 238 1748 254
rect 1682 204 1698 238
rect 1732 204 1748 238
rect 1682 188 1748 204
rect 1800 238 1866 254
rect 1800 204 1816 238
rect 1850 204 1866 238
rect 1800 188 1866 204
rect 1918 238 1984 254
rect 1918 204 1934 238
rect 1968 204 1984 238
rect 1918 188 1984 204
rect 2036 238 2102 254
rect 2036 204 2052 238
rect 2086 204 2102 238
rect 2036 188 2102 204
rect 2154 238 2220 254
rect 2154 204 2170 238
rect 2204 204 2220 238
rect 2154 188 2220 204
rect 2272 238 2338 254
rect 2272 204 2288 238
rect 2322 204 2338 238
rect 2272 188 2338 204
rect 2390 238 2456 254
rect 2390 204 2406 238
rect 2440 204 2456 238
rect 2390 188 2456 204
rect 2508 238 2574 254
rect 2508 204 2524 238
rect 2558 204 2574 238
rect 2508 188 2574 204
rect 2626 238 2692 254
rect 2626 204 2642 238
rect 2676 204 2692 238
rect 2626 188 2692 204
rect 2744 238 2810 254
rect 2744 204 2760 238
rect 2794 204 2810 238
rect 2744 188 2810 204
rect 2862 238 2928 254
rect 2862 204 2878 238
rect 2912 204 2928 238
rect 2862 188 2928 204
rect 2980 238 3046 254
rect 2980 204 2996 238
rect 3030 204 3046 238
rect 2980 188 3046 204
rect 3098 238 3164 254
rect 3098 204 3114 238
rect 3148 204 3164 238
rect 3098 188 3164 204
rect 3216 238 3282 254
rect 3216 204 3232 238
rect 3266 204 3282 238
rect 3216 188 3282 204
rect 3334 238 3400 254
rect 3334 204 3350 238
rect 3384 204 3400 238
rect 3334 188 3400 204
rect 3452 238 3518 254
rect 3452 204 3468 238
rect 3502 204 3518 238
rect 3452 188 3518 204
rect 3570 238 3636 254
rect 3570 204 3586 238
rect 3620 204 3636 238
rect 3570 188 3636 204
rect 3688 238 3754 254
rect 3688 204 3704 238
rect 3738 204 3754 238
rect 3688 188 3754 204
rect 3806 238 3872 254
rect 3806 204 3822 238
rect 3856 204 3872 238
rect 3806 188 3872 204
rect 3924 238 3990 254
rect 3924 204 3940 238
rect 3974 204 3990 238
rect 3924 188 3990 204
rect 4042 238 4108 254
rect 4042 204 4058 238
rect 4092 204 4108 238
rect 4042 188 4108 204
rect 4160 238 4226 254
rect 4160 204 4176 238
rect 4210 204 4226 238
rect 4160 188 4226 204
rect 4278 238 4344 254
rect 4278 204 4294 238
rect 4328 204 4344 238
rect 4278 188 4344 204
rect 4396 238 4462 254
rect 4396 204 4412 238
rect 4446 204 4462 238
rect 4396 188 4462 204
rect 4514 238 4580 254
rect 4514 204 4530 238
rect 4564 204 4580 238
rect 4514 188 4580 204
rect 4632 238 4698 254
rect 4632 204 4648 238
rect 4682 204 4698 238
rect 4632 188 4698 204
rect 4750 238 4816 254
rect 4750 204 4766 238
rect 4800 204 4816 238
rect 4750 188 4816 204
rect 4868 238 4934 254
rect 4868 204 4884 238
rect 4918 204 4934 238
rect 4868 188 4934 204
rect 4986 238 5052 254
rect 4986 204 5002 238
rect 5036 204 5052 238
rect 4986 188 5052 204
rect 5104 238 5170 254
rect 5104 204 5120 238
rect 5154 204 5170 238
rect 5104 188 5170 204
rect 29 -152 95 -136
rect 29 -186 45 -152
rect 79 -186 95 -152
rect 29 -202 95 -186
rect 147 -152 213 -136
rect 147 -186 163 -152
rect 197 -186 213 -152
rect 147 -202 213 -186
rect 265 -152 331 -136
rect 265 -186 281 -152
rect 315 -186 331 -152
rect 265 -202 331 -186
rect 383 -152 449 -136
rect 383 -186 399 -152
rect 433 -186 449 -152
rect 383 -202 449 -186
rect 501 -152 567 -136
rect 501 -186 517 -152
rect 551 -186 567 -152
rect 501 -202 567 -186
rect 619 -152 685 -136
rect 619 -186 635 -152
rect 669 -186 685 -152
rect 619 -202 685 -186
rect 737 -152 803 -136
rect 737 -186 753 -152
rect 787 -186 803 -152
rect 737 -202 803 -186
rect 855 -152 921 -136
rect 855 -186 871 -152
rect 905 -186 921 -152
rect 855 -202 921 -186
rect 973 -152 1039 -136
rect 973 -186 989 -152
rect 1023 -186 1039 -152
rect 973 -202 1039 -186
rect 1091 -152 1157 -136
rect 1091 -186 1107 -152
rect 1141 -186 1157 -152
rect 1091 -202 1157 -186
rect 32 -224 92 -202
rect 150 -224 210 -202
rect 268 -224 328 -202
rect 386 -224 446 -202
rect 504 -224 564 -202
rect 622 -224 682 -202
rect 740 -224 800 -202
rect 858 -224 918 -202
rect 976 -224 1036 -202
rect 1094 -224 1154 -202
rect 32 -2246 92 -2224
rect 150 -2246 210 -2224
rect 268 -2246 328 -2224
rect 386 -2246 446 -2224
rect 504 -2246 564 -2224
rect 622 -2246 682 -2224
rect 740 -2246 800 -2224
rect 858 -2246 918 -2224
rect 976 -2246 1036 -2224
rect 1094 -2246 1154 -2224
rect 29 -2262 95 -2246
rect 29 -2296 45 -2262
rect 79 -2296 95 -2262
rect 29 -2312 95 -2296
rect 147 -2262 213 -2246
rect 147 -2296 163 -2262
rect 197 -2296 213 -2262
rect 147 -2312 213 -2296
rect 265 -2262 331 -2246
rect 265 -2296 281 -2262
rect 315 -2296 331 -2262
rect 265 -2312 331 -2296
rect 383 -2262 449 -2246
rect 383 -2296 399 -2262
rect 433 -2296 449 -2262
rect 383 -2312 449 -2296
rect 501 -2262 567 -2246
rect 501 -2296 517 -2262
rect 551 -2296 567 -2262
rect 501 -2312 567 -2296
rect 619 -2262 685 -2246
rect 619 -2296 635 -2262
rect 669 -2296 685 -2262
rect 619 -2312 685 -2296
rect 737 -2262 803 -2246
rect 737 -2296 753 -2262
rect 787 -2296 803 -2262
rect 737 -2312 803 -2296
rect 855 -2262 921 -2246
rect 855 -2296 871 -2262
rect 905 -2296 921 -2262
rect 855 -2312 921 -2296
rect 973 -2262 1039 -2246
rect 973 -2296 989 -2262
rect 1023 -2296 1039 -2262
rect 973 -2312 1039 -2296
rect 1091 -2262 1157 -2246
rect 1091 -2296 1107 -2262
rect 1141 -2296 1157 -2262
rect 1091 -2312 1157 -2296
rect 1673 -324 1799 -296
rect 1673 -358 1719 -324
rect 1753 -358 1799 -324
rect 1673 -374 1799 -358
rect 3401 -324 3527 -296
rect 3401 -358 3447 -324
rect 3481 -358 3527 -324
rect 3401 -374 3527 -358
rect 1673 -400 1703 -374
rect 1769 -400 1799 -374
rect 1865 -400 1895 -374
rect 1961 -400 1991 -374
rect 2057 -400 2087 -374
rect 2153 -400 2183 -374
rect 2249 -400 2279 -374
rect 2345 -400 2375 -374
rect 2441 -400 2471 -374
rect 2537 -400 2567 -374
rect 2633 -400 2663 -374
rect 2729 -400 2759 -374
rect 2825 -400 2855 -374
rect 2921 -400 2951 -374
rect 3017 -400 3047 -374
rect 3113 -400 3143 -374
rect 3209 -400 3239 -374
rect 3305 -400 3335 -374
rect 3401 -400 3431 -374
rect 3497 -400 3527 -374
rect 1673 -926 1703 -900
rect 1769 -926 1799 -900
rect 1865 -922 1895 -900
rect 1961 -922 1991 -900
rect 1865 -950 1991 -922
rect 1865 -984 1911 -950
rect 1945 -984 1991 -950
rect 1865 -1000 1991 -984
rect 2057 -922 2087 -900
rect 2153 -922 2183 -900
rect 2057 -950 2183 -922
rect 2057 -984 2103 -950
rect 2137 -984 2183 -950
rect 2057 -1000 2183 -984
rect 2249 -922 2279 -900
rect 2345 -922 2375 -900
rect 2249 -950 2375 -922
rect 2249 -984 2295 -950
rect 2329 -984 2375 -950
rect 2249 -1000 2375 -984
rect 2441 -922 2471 -900
rect 2537 -922 2567 -900
rect 2441 -950 2567 -922
rect 2441 -984 2487 -950
rect 2521 -984 2567 -950
rect 2441 -1000 2567 -984
rect 2633 -922 2663 -900
rect 2729 -922 2759 -900
rect 2633 -950 2759 -922
rect 2633 -984 2679 -950
rect 2713 -984 2759 -950
rect 2633 -1000 2759 -984
rect 2825 -922 2855 -900
rect 2921 -922 2951 -900
rect 2825 -950 2951 -922
rect 2825 -984 2871 -950
rect 2905 -984 2951 -950
rect 2825 -1000 2951 -984
rect 3017 -922 3047 -900
rect 3113 -922 3143 -900
rect 3017 -950 3143 -922
rect 3017 -984 3063 -950
rect 3097 -984 3143 -950
rect 3017 -1000 3143 -984
rect 3209 -922 3239 -900
rect 3305 -922 3335 -900
rect 3209 -950 3335 -922
rect 3401 -926 3431 -900
rect 3497 -926 3527 -900
rect 3209 -984 3255 -950
rect 3289 -984 3335 -950
rect 3209 -1000 3335 -984
rect 1713 -1268 2113 -1252
rect 1713 -1302 1729 -1268
rect 2097 -1302 2113 -1268
rect 1713 -1340 2113 -1302
rect 2171 -1268 2571 -1252
rect 2171 -1302 2187 -1268
rect 2555 -1302 2571 -1268
rect 2171 -1340 2571 -1302
rect 2629 -1268 3029 -1252
rect 2629 -1302 2645 -1268
rect 3013 -1302 3029 -1268
rect 2629 -1340 3029 -1302
rect 3087 -1268 3487 -1252
rect 3087 -1302 3103 -1268
rect 3471 -1302 3487 -1268
rect 3087 -1340 3487 -1302
rect 1713 -3378 2113 -3340
rect 1713 -3412 1729 -3378
rect 2097 -3412 2113 -3378
rect 1713 -3428 2113 -3412
rect 2171 -3378 2571 -3340
rect 2171 -3412 2187 -3378
rect 2555 -3412 2571 -3378
rect 2171 -3428 2571 -3412
rect 2629 -3378 3029 -3340
rect 2629 -3412 2645 -3378
rect 3013 -3412 3029 -3378
rect 2629 -3428 3029 -3412
rect 3087 -3378 3487 -3340
rect 3087 -3412 3103 -3378
rect 3471 -3412 3487 -3378
rect 3087 -3428 3487 -3412
rect 4042 -152 4108 -136
rect 4042 -186 4058 -152
rect 4092 -186 4108 -152
rect 4042 -202 4108 -186
rect 4160 -152 4226 -136
rect 4160 -186 4176 -152
rect 4210 -186 4226 -152
rect 4160 -202 4226 -186
rect 4278 -152 4344 -136
rect 4278 -186 4294 -152
rect 4328 -186 4344 -152
rect 4278 -202 4344 -186
rect 4396 -152 4462 -136
rect 4396 -186 4412 -152
rect 4446 -186 4462 -152
rect 4396 -202 4462 -186
rect 4514 -152 4580 -136
rect 4514 -186 4530 -152
rect 4564 -186 4580 -152
rect 4514 -202 4580 -186
rect 4632 -152 4698 -136
rect 4632 -186 4648 -152
rect 4682 -186 4698 -152
rect 4632 -202 4698 -186
rect 4750 -152 4816 -136
rect 4750 -186 4766 -152
rect 4800 -186 4816 -152
rect 4750 -202 4816 -186
rect 4868 -152 4934 -136
rect 4868 -186 4884 -152
rect 4918 -186 4934 -152
rect 4868 -202 4934 -186
rect 4986 -152 5052 -136
rect 4986 -186 5002 -152
rect 5036 -186 5052 -152
rect 4986 -202 5052 -186
rect 5104 -152 5170 -136
rect 5104 -186 5120 -152
rect 5154 -186 5170 -152
rect 5104 -202 5170 -186
rect 4045 -224 4105 -202
rect 4163 -224 4223 -202
rect 4281 -224 4341 -202
rect 4399 -224 4459 -202
rect 4517 -224 4577 -202
rect 4635 -224 4695 -202
rect 4753 -224 4813 -202
rect 4871 -224 4931 -202
rect 4989 -224 5049 -202
rect 5107 -224 5167 -202
rect 4045 -2246 4105 -2224
rect 4163 -2246 4223 -2224
rect 4281 -2246 4341 -2224
rect 4399 -2246 4459 -2224
rect 4517 -2246 4577 -2224
rect 4635 -2246 4695 -2224
rect 4753 -2246 4813 -2224
rect 4871 -2246 4931 -2224
rect 4989 -2246 5049 -2224
rect 5107 -2246 5167 -2224
rect 4042 -2262 4108 -2246
rect 4042 -2296 4058 -2262
rect 4092 -2296 4108 -2262
rect 4042 -2312 4108 -2296
rect 4160 -2262 4226 -2246
rect 4160 -2296 4176 -2262
rect 4210 -2296 4226 -2262
rect 4160 -2312 4226 -2296
rect 4278 -2262 4344 -2246
rect 4278 -2296 4294 -2262
rect 4328 -2296 4344 -2262
rect 4278 -2312 4344 -2296
rect 4396 -2262 4462 -2246
rect 4396 -2296 4412 -2262
rect 4446 -2296 4462 -2262
rect 4396 -2312 4462 -2296
rect 4514 -2262 4580 -2246
rect 4514 -2296 4530 -2262
rect 4564 -2296 4580 -2262
rect 4514 -2312 4580 -2296
rect 4632 -2262 4698 -2246
rect 4632 -2296 4648 -2262
rect 4682 -2296 4698 -2262
rect 4632 -2312 4698 -2296
rect 4750 -2262 4816 -2246
rect 4750 -2296 4766 -2262
rect 4800 -2296 4816 -2262
rect 4750 -2312 4816 -2296
rect 4868 -2262 4934 -2246
rect 4868 -2296 4884 -2262
rect 4918 -2296 4934 -2262
rect 4868 -2312 4934 -2296
rect 4986 -2262 5052 -2246
rect 4986 -2296 5002 -2262
rect 5036 -2296 5052 -2262
rect 4986 -2312 5052 -2296
rect 5104 -2262 5170 -2246
rect 5104 -2296 5120 -2262
rect 5154 -2296 5170 -2262
rect 5104 -2312 5170 -2296
<< polycont >>
rect 46 2332 80 2366
rect 164 2332 198 2366
rect 282 2332 316 2366
rect 400 2332 434 2366
rect 518 2332 552 2366
rect 636 2332 670 2366
rect 754 2332 788 2366
rect 872 2332 906 2366
rect 990 2332 1024 2366
rect 1108 2332 1142 2366
rect 1226 2332 1260 2366
rect 1344 2332 1378 2366
rect 1462 2332 1496 2366
rect 1580 2332 1614 2366
rect 1698 2332 1732 2366
rect 1816 2332 1850 2366
rect 1934 2332 1968 2366
rect 2052 2332 2086 2366
rect 2170 2332 2204 2366
rect 2288 2332 2322 2366
rect 2878 2332 2912 2366
rect 2996 2332 3030 2366
rect 3114 2332 3148 2366
rect 3232 2332 3266 2366
rect 3350 2332 3384 2366
rect 3468 2332 3502 2366
rect 3586 2332 3620 2366
rect 3704 2332 3738 2366
rect 3822 2332 3856 2366
rect 3940 2332 3974 2366
rect 4058 2332 4092 2366
rect 4176 2332 4210 2366
rect 4294 2332 4328 2366
rect 4412 2332 4446 2366
rect 4530 2332 4564 2366
rect 4648 2332 4682 2366
rect 4766 2332 4800 2366
rect 4884 2332 4918 2366
rect 5002 2332 5036 2366
rect 5120 2332 5154 2366
rect 46 204 80 238
rect 164 204 198 238
rect 282 204 316 238
rect 400 204 434 238
rect 518 204 552 238
rect 636 204 670 238
rect 754 204 788 238
rect 872 204 906 238
rect 990 204 1024 238
rect 1108 204 1142 238
rect 1226 204 1260 238
rect 1344 204 1378 238
rect 1462 204 1496 238
rect 1580 204 1614 238
rect 1698 204 1732 238
rect 1816 204 1850 238
rect 1934 204 1968 238
rect 2052 204 2086 238
rect 2170 204 2204 238
rect 2288 204 2322 238
rect 2406 204 2440 238
rect 2524 204 2558 238
rect 2642 204 2676 238
rect 2760 204 2794 238
rect 2878 204 2912 238
rect 2996 204 3030 238
rect 3114 204 3148 238
rect 3232 204 3266 238
rect 3350 204 3384 238
rect 3468 204 3502 238
rect 3586 204 3620 238
rect 3704 204 3738 238
rect 3822 204 3856 238
rect 3940 204 3974 238
rect 4058 204 4092 238
rect 4176 204 4210 238
rect 4294 204 4328 238
rect 4412 204 4446 238
rect 4530 204 4564 238
rect 4648 204 4682 238
rect 4766 204 4800 238
rect 4884 204 4918 238
rect 5002 204 5036 238
rect 5120 204 5154 238
rect 45 -186 79 -152
rect 163 -186 197 -152
rect 281 -186 315 -152
rect 399 -186 433 -152
rect 517 -186 551 -152
rect 635 -186 669 -152
rect 753 -186 787 -152
rect 871 -186 905 -152
rect 989 -186 1023 -152
rect 1107 -186 1141 -152
rect 45 -2296 79 -2262
rect 163 -2296 197 -2262
rect 281 -2296 315 -2262
rect 399 -2296 433 -2262
rect 517 -2296 551 -2262
rect 635 -2296 669 -2262
rect 753 -2296 787 -2262
rect 871 -2296 905 -2262
rect 989 -2296 1023 -2262
rect 1107 -2296 1141 -2262
rect 1719 -358 1753 -324
rect 3447 -358 3481 -324
rect 1911 -984 1945 -950
rect 2103 -984 2137 -950
rect 2295 -984 2329 -950
rect 2487 -984 2521 -950
rect 2679 -984 2713 -950
rect 2871 -984 2905 -950
rect 3063 -984 3097 -950
rect 3255 -984 3289 -950
rect 1729 -1302 2097 -1268
rect 2187 -1302 2555 -1268
rect 2645 -1302 3013 -1268
rect 3103 -1302 3471 -1268
rect 1729 -3412 2097 -3378
rect 2187 -3412 2555 -3378
rect 2645 -3412 3013 -3378
rect 3103 -3412 3471 -3378
rect 4058 -186 4092 -152
rect 4176 -186 4210 -152
rect 4294 -186 4328 -152
rect 4412 -186 4446 -152
rect 4530 -186 4564 -152
rect 4648 -186 4682 -152
rect 4766 -186 4800 -152
rect 4884 -186 4918 -152
rect 5002 -186 5036 -152
rect 5120 -186 5154 -152
rect 4058 -2296 4092 -2262
rect 4176 -2296 4210 -2262
rect 4294 -2296 4328 -2262
rect 4412 -2296 4446 -2262
rect 4530 -2296 4564 -2262
rect 4648 -2296 4682 -2262
rect 4766 -2296 4800 -2262
rect 4884 -2296 4918 -2262
rect 5002 -2296 5036 -2262
rect 5120 -2296 5154 -2262
<< locali >>
rect -127 2434 -31 2468
rect 5231 2434 5327 2468
rect -127 2372 -93 2434
rect 5293 2372 5327 2434
rect 30 2332 46 2366
rect 80 2332 96 2366
rect 148 2332 164 2366
rect 198 2332 214 2366
rect 266 2332 282 2366
rect 316 2332 332 2366
rect 384 2332 400 2366
rect 434 2332 450 2366
rect 502 2332 518 2366
rect 552 2332 568 2366
rect 620 2332 636 2366
rect 670 2332 686 2366
rect 738 2332 754 2366
rect 788 2332 804 2366
rect 856 2332 872 2366
rect 906 2332 922 2366
rect 974 2332 990 2366
rect 1024 2332 1040 2366
rect 1092 2332 1108 2366
rect 1142 2332 1158 2366
rect 1210 2332 1226 2366
rect 1260 2332 1276 2366
rect 1328 2332 1344 2366
rect 1378 2332 1394 2366
rect 1446 2332 1462 2366
rect 1496 2332 1512 2366
rect 1564 2332 1580 2366
rect 1614 2332 1630 2366
rect 1682 2332 1698 2366
rect 1732 2332 1748 2366
rect 1800 2332 1816 2366
rect 1850 2332 1866 2366
rect 1918 2332 1934 2366
rect 1968 2332 1984 2366
rect 2036 2332 2052 2366
rect 2086 2332 2102 2366
rect 2154 2332 2170 2366
rect 2204 2332 2220 2366
rect 2272 2332 2288 2366
rect 2322 2332 2338 2366
rect 2862 2332 2878 2366
rect 2912 2332 2928 2366
rect 2980 2332 2996 2366
rect 3030 2332 3046 2366
rect 3098 2332 3114 2366
rect 3148 2332 3164 2366
rect 3216 2332 3232 2366
rect 3266 2332 3282 2366
rect 3334 2332 3350 2366
rect 3384 2332 3400 2366
rect 3452 2332 3468 2366
rect 3502 2332 3518 2366
rect 3570 2332 3586 2366
rect 3620 2332 3636 2366
rect 3688 2332 3704 2366
rect 3738 2332 3754 2366
rect 3806 2332 3822 2366
rect 3856 2332 3872 2366
rect 3924 2332 3940 2366
rect 3974 2332 3990 2366
rect 4042 2332 4058 2366
rect 4092 2332 4108 2366
rect 4160 2332 4176 2366
rect 4210 2332 4226 2366
rect 4278 2332 4294 2366
rect 4328 2332 4344 2366
rect 4396 2332 4412 2366
rect 4446 2332 4462 2366
rect 4514 2332 4530 2366
rect 4564 2332 4580 2366
rect 4632 2332 4648 2366
rect 4682 2332 4698 2366
rect 4750 2332 4766 2366
rect 4800 2332 4816 2366
rect 4868 2332 4884 2366
rect 4918 2332 4934 2366
rect 4986 2332 5002 2366
rect 5036 2332 5052 2366
rect 5104 2332 5120 2366
rect 5154 2332 5170 2366
rect -13 2273 21 2289
rect -13 281 21 297
rect 105 2273 139 2289
rect 105 281 139 297
rect 223 2273 257 2289
rect 223 281 257 297
rect 341 2273 375 2289
rect 341 281 375 297
rect 459 2273 493 2289
rect 459 281 493 297
rect 577 2273 611 2289
rect 577 281 611 297
rect 695 2273 729 2289
rect 695 281 729 297
rect 813 2273 847 2289
rect 813 281 847 297
rect 931 2273 965 2289
rect 931 281 965 297
rect 1049 2273 1083 2289
rect 1049 281 1083 297
rect 1167 2273 1201 2289
rect 1167 281 1201 297
rect 1285 2273 1319 2289
rect 1285 281 1319 297
rect 1403 2273 1437 2289
rect 1403 281 1437 297
rect 1521 2273 1555 2289
rect 1521 281 1555 297
rect 1639 2273 1673 2289
rect 1639 281 1673 297
rect 1757 2273 1791 2289
rect 1757 281 1791 297
rect 1875 2273 1909 2289
rect 1875 281 1909 297
rect 1993 2273 2027 2289
rect 1993 281 2027 297
rect 2111 2273 2145 2289
rect 2111 281 2145 297
rect 2229 2273 2263 2289
rect 2229 281 2263 297
rect 2347 2273 2381 2289
rect 2347 281 2381 297
rect 2465 2273 2499 2289
rect 2465 281 2499 297
rect 2583 2273 2617 2289
rect 2583 281 2617 297
rect 2701 2273 2735 2289
rect 2701 281 2735 297
rect 2819 2273 2853 2289
rect 2819 281 2853 297
rect 2937 2273 2971 2289
rect 2937 281 2971 297
rect 3055 2273 3089 2289
rect 3055 281 3089 297
rect 3173 2273 3207 2289
rect 3173 281 3207 297
rect 3291 2273 3325 2289
rect 3291 281 3325 297
rect 3409 2273 3443 2289
rect 3409 281 3443 297
rect 3527 2273 3561 2289
rect 3527 281 3561 297
rect 3645 2273 3679 2289
rect 3645 281 3679 297
rect 3763 2273 3797 2289
rect 3763 281 3797 297
rect 3881 2273 3915 2289
rect 3881 281 3915 297
rect 3999 2273 4033 2289
rect 3999 281 4033 297
rect 4117 2273 4151 2289
rect 4117 281 4151 297
rect 4235 2273 4269 2289
rect 4235 281 4269 297
rect 4353 2273 4387 2289
rect 4353 281 4387 297
rect 4471 2273 4505 2289
rect 4471 281 4505 297
rect 4589 2273 4623 2289
rect 4589 281 4623 297
rect 4707 2273 4741 2289
rect 4707 281 4741 297
rect 4825 2273 4859 2289
rect 4825 281 4859 297
rect 4943 2273 4977 2289
rect 4943 281 4977 297
rect 5061 2273 5095 2289
rect 5061 281 5095 297
rect 5179 2273 5213 2289
rect 5179 281 5213 297
rect 30 204 46 238
rect 80 204 96 238
rect 148 204 164 238
rect 198 204 214 238
rect 266 204 282 238
rect 316 204 332 238
rect 384 204 400 238
rect 434 204 450 238
rect 502 204 518 238
rect 552 204 568 238
rect 620 204 636 238
rect 670 204 686 238
rect 738 204 754 238
rect 788 204 804 238
rect 856 204 872 238
rect 906 204 922 238
rect 974 204 990 238
rect 1024 204 1040 238
rect 1092 204 1108 238
rect 1142 204 1158 238
rect 1210 204 1226 238
rect 1260 204 1276 238
rect 1328 204 1344 238
rect 1378 204 1394 238
rect 1446 204 1462 238
rect 1496 204 1512 238
rect 1564 204 1580 238
rect 1614 204 1630 238
rect 1682 204 1698 238
rect 1732 204 1748 238
rect 1800 204 1816 238
rect 1850 204 1866 238
rect 1918 204 1934 238
rect 1968 204 1984 238
rect 2036 204 2052 238
rect 2086 204 2102 238
rect 2154 204 2170 238
rect 2204 204 2220 238
rect 2272 204 2288 238
rect 2322 204 2338 238
rect 2390 204 2406 238
rect 2440 204 2456 238
rect 2508 204 2524 238
rect 2558 204 2574 238
rect 2626 204 2642 238
rect 2676 204 2692 238
rect 2744 204 2760 238
rect 2794 204 2810 238
rect 2862 204 2878 238
rect 2912 204 2928 238
rect 2980 204 2996 238
rect 3030 204 3046 238
rect 3098 204 3114 238
rect 3148 204 3164 238
rect 3216 204 3232 238
rect 3266 204 3282 238
rect 3334 204 3350 238
rect 3384 204 3400 238
rect 3452 204 3468 238
rect 3502 204 3518 238
rect 3570 204 3586 238
rect 3620 204 3636 238
rect 3688 204 3704 238
rect 3738 204 3754 238
rect 3806 204 3822 238
rect 3856 204 3872 238
rect 3924 204 3940 238
rect 3974 204 3990 238
rect 4042 204 4058 238
rect 4092 204 4108 238
rect 4160 204 4176 238
rect 4210 204 4226 238
rect 4278 204 4294 238
rect 4328 204 4344 238
rect 4396 204 4412 238
rect 4446 204 4462 238
rect 4514 204 4530 238
rect 4564 204 4580 238
rect 4632 204 4648 238
rect 4682 204 4698 238
rect 4750 204 4766 238
rect 4800 204 4816 238
rect 4868 204 4884 238
rect 4918 204 4934 238
rect 4986 204 5002 238
rect 5036 204 5052 238
rect 5104 204 5120 238
rect 5154 204 5170 238
rect -127 136 -93 198
rect 5293 136 5327 198
rect -127 102 -31 136
rect 5231 102 5327 136
rect -128 -84 -32 -50
rect 1218 -84 1314 -50
rect -128 -146 -94 -84
rect 1280 -146 1314 -84
rect 29 -186 45 -152
rect 79 -186 95 -152
rect 147 -186 163 -152
rect 197 -186 213 -152
rect 265 -186 281 -152
rect 315 -186 331 -152
rect 383 -186 399 -152
rect 433 -186 449 -152
rect 501 -186 517 -152
rect 551 -186 567 -152
rect 619 -186 635 -152
rect 669 -186 685 -152
rect 737 -186 753 -152
rect 787 -186 803 -152
rect 855 -186 871 -152
rect 905 -186 921 -152
rect 973 -186 989 -152
rect 1023 -186 1039 -152
rect 1091 -186 1107 -152
rect 1141 -186 1157 -152
rect -14 -236 20 -220
rect -14 -2228 20 -2212
rect 104 -236 138 -220
rect 104 -2228 138 -2212
rect 222 -236 256 -220
rect 222 -2228 256 -2212
rect 340 -236 374 -220
rect 340 -2228 374 -2212
rect 458 -236 492 -220
rect 458 -2228 492 -2212
rect 576 -236 610 -220
rect 576 -2228 610 -2212
rect 694 -236 728 -220
rect 694 -2228 728 -2212
rect 812 -236 846 -220
rect 812 -2228 846 -2212
rect 930 -236 964 -220
rect 930 -2228 964 -2212
rect 1048 -236 1082 -220
rect 1048 -2228 1082 -2212
rect 1166 -236 1200 -220
rect 1166 -2228 1200 -2212
rect 3885 -84 3981 -50
rect 5231 -84 5327 -50
rect 3885 -146 3919 -84
rect 5293 -146 5327 -84
rect 4042 -186 4058 -152
rect 4092 -186 4108 -152
rect 4160 -186 4176 -152
rect 4210 -186 4226 -152
rect 4278 -186 4294 -152
rect 4328 -186 4344 -152
rect 4396 -186 4412 -152
rect 4446 -186 4462 -152
rect 4514 -186 4530 -152
rect 4564 -186 4580 -152
rect 4632 -186 4648 -152
rect 4682 -186 4698 -152
rect 4750 -186 4766 -152
rect 4800 -186 4816 -152
rect 4868 -186 4884 -152
rect 4918 -186 4934 -152
rect 4986 -186 5002 -152
rect 5036 -186 5052 -152
rect 5104 -186 5120 -152
rect 5154 -186 5170 -152
rect 1509 -260 1605 -226
rect 3595 -260 3691 -226
rect 1509 -322 1543 -260
rect 3657 -322 3691 -260
rect 1703 -358 1719 -324
rect 1753 -358 1769 -324
rect 3431 -358 3447 -324
rect 3481 -358 3497 -324
rect 1623 -412 1657 -396
rect 1623 -904 1657 -888
rect 1719 -412 1753 -396
rect 1719 -904 1753 -888
rect 1815 -412 1849 -396
rect 1815 -904 1849 -888
rect 1911 -412 1945 -396
rect 1911 -904 1945 -888
rect 2007 -412 2041 -396
rect 2007 -904 2041 -888
rect 2103 -412 2137 -396
rect 2103 -904 2137 -888
rect 2199 -412 2233 -396
rect 2199 -904 2233 -888
rect 2295 -412 2329 -396
rect 2295 -904 2329 -888
rect 2391 -412 2425 -396
rect 2391 -904 2425 -888
rect 2487 -412 2521 -396
rect 2487 -904 2521 -888
rect 2583 -412 2617 -396
rect 2583 -904 2617 -888
rect 2679 -412 2713 -396
rect 2679 -904 2713 -888
rect 2775 -412 2809 -396
rect 2775 -904 2809 -888
rect 2871 -412 2905 -396
rect 2871 -904 2905 -888
rect 2967 -412 3001 -396
rect 2967 -904 3001 -888
rect 3063 -412 3097 -396
rect 3063 -904 3097 -888
rect 3159 -412 3193 -396
rect 3159 -904 3193 -888
rect 3255 -412 3289 -396
rect 3255 -904 3289 -888
rect 3351 -412 3385 -396
rect 3351 -904 3385 -888
rect 3447 -412 3481 -396
rect 3447 -904 3481 -888
rect 3543 -412 3577 -396
rect 3543 -904 3577 -888
rect 1509 -1040 1543 -978
rect 1895 -984 1911 -950
rect 1945 -984 1961 -950
rect 2087 -984 2103 -950
rect 2137 -984 2153 -950
rect 2279 -984 2295 -950
rect 2329 -984 2345 -950
rect 2471 -984 2487 -950
rect 2521 -984 2537 -950
rect 2663 -984 2679 -950
rect 2713 -984 2729 -950
rect 2855 -984 2871 -950
rect 2905 -984 2921 -950
rect 3047 -984 3063 -950
rect 3097 -984 3113 -950
rect 3239 -984 3255 -950
rect 3289 -984 3305 -950
rect 3657 -1040 3691 -978
rect 1509 -1074 1605 -1040
rect 3595 -1074 3691 -1040
rect 29 -2296 45 -2262
rect 79 -2296 95 -2262
rect 147 -2296 163 -2262
rect 197 -2296 213 -2262
rect 265 -2296 281 -2262
rect 315 -2296 331 -2262
rect 383 -2296 399 -2262
rect 433 -2296 449 -2262
rect 501 -2296 517 -2262
rect 551 -2296 567 -2262
rect 619 -2296 635 -2262
rect 669 -2296 685 -2262
rect 737 -2296 753 -2262
rect 787 -2296 803 -2262
rect 855 -2296 871 -2262
rect 905 -2296 921 -2262
rect 973 -2296 989 -2262
rect 1023 -2296 1039 -2262
rect 1091 -2296 1107 -2262
rect 1141 -2296 1157 -2262
rect -128 -2364 -94 -2302
rect 1280 -2364 1314 -2302
rect -128 -2398 -32 -2364
rect 1218 -2398 1314 -2364
rect 1553 -1200 1649 -1166
rect 3551 -1200 3647 -1166
rect 1553 -1262 1587 -1200
rect 3613 -1262 3647 -1200
rect 1713 -1302 1729 -1268
rect 2097 -1302 2113 -1268
rect 2171 -1302 2187 -1268
rect 2555 -1302 2571 -1268
rect 2629 -1302 2645 -1268
rect 3013 -1302 3029 -1268
rect 3087 -1302 3103 -1268
rect 3471 -1302 3487 -1268
rect 1667 -1352 1701 -1336
rect 1667 -3344 1701 -3328
rect 2125 -1352 2159 -1336
rect 2125 -3344 2159 -3328
rect 2583 -1352 2617 -1336
rect 2583 -3344 2617 -3328
rect 3041 -1352 3075 -1336
rect 3041 -3344 3075 -3328
rect 3499 -1352 3533 -1336
rect 3499 -3344 3533 -3328
rect 3999 -236 4033 -220
rect 3999 -2228 4033 -2212
rect 4117 -236 4151 -220
rect 4117 -2228 4151 -2212
rect 4235 -236 4269 -220
rect 4235 -2228 4269 -2212
rect 4353 -236 4387 -220
rect 4353 -2228 4387 -2212
rect 4471 -236 4505 -220
rect 4471 -2228 4505 -2212
rect 4589 -236 4623 -220
rect 4589 -2228 4623 -2212
rect 4707 -236 4741 -220
rect 4707 -2228 4741 -2212
rect 4825 -236 4859 -220
rect 4825 -2228 4859 -2212
rect 4943 -236 4977 -220
rect 4943 -2228 4977 -2212
rect 5061 -236 5095 -220
rect 5061 -2228 5095 -2212
rect 5179 -236 5213 -220
rect 5179 -2228 5213 -2212
rect 4042 -2296 4058 -2262
rect 4092 -2296 4108 -2262
rect 4160 -2296 4176 -2262
rect 4210 -2296 4226 -2262
rect 4278 -2296 4294 -2262
rect 4328 -2296 4344 -2262
rect 4396 -2296 4412 -2262
rect 4446 -2296 4462 -2262
rect 4514 -2296 4530 -2262
rect 4564 -2296 4580 -2262
rect 4632 -2296 4648 -2262
rect 4682 -2296 4698 -2262
rect 4750 -2296 4766 -2262
rect 4800 -2296 4816 -2262
rect 4868 -2296 4884 -2262
rect 4918 -2296 4934 -2262
rect 4986 -2296 5002 -2262
rect 5036 -2296 5052 -2262
rect 5104 -2296 5120 -2262
rect 5154 -2296 5170 -2262
rect 3885 -2364 3919 -2302
rect 5293 -2364 5327 -2302
rect 3885 -2398 3981 -2364
rect 5231 -2398 5327 -2364
rect 1713 -3412 1729 -3378
rect 2097 -3412 2113 -3378
rect 2171 -3412 2187 -3378
rect 2555 -3412 2571 -3378
rect 2629 -3412 2645 -3378
rect 3013 -3412 3029 -3378
rect 3087 -3412 3103 -3378
rect 3471 -3412 3487 -3378
rect 1553 -3480 1587 -3418
rect 3613 -3480 3647 -3418
rect 1553 -3514 1649 -3480
rect 3551 -3514 3647 -3480
<< viali >>
rect 46 2332 80 2366
rect 164 2332 198 2366
rect 282 2332 316 2366
rect 400 2332 434 2366
rect 518 2332 552 2366
rect 636 2332 670 2366
rect 754 2332 788 2366
rect 872 2332 906 2366
rect 990 2332 1024 2366
rect 1108 2332 1142 2366
rect 1226 2332 1260 2366
rect 1344 2332 1378 2366
rect 1462 2332 1496 2366
rect 1580 2332 1614 2366
rect 1698 2332 1732 2366
rect 1816 2332 1850 2366
rect 1934 2332 1968 2366
rect 2052 2332 2086 2366
rect 2170 2332 2204 2366
rect 2288 2332 2322 2366
rect 2878 2332 2912 2366
rect 2996 2332 3030 2366
rect 3114 2332 3148 2366
rect 3232 2332 3266 2366
rect 3350 2332 3384 2366
rect 3468 2332 3502 2366
rect 3586 2332 3620 2366
rect 3704 2332 3738 2366
rect 3822 2332 3856 2366
rect 3940 2332 3974 2366
rect 4058 2332 4092 2366
rect 4176 2332 4210 2366
rect 4294 2332 4328 2366
rect 4412 2332 4446 2366
rect 4530 2332 4564 2366
rect 4648 2332 4682 2366
rect 4766 2332 4800 2366
rect 4884 2332 4918 2366
rect 5002 2332 5036 2366
rect 5120 2332 5154 2366
rect -127 1885 -93 2285
rect -127 285 -93 685
rect -13 297 21 2273
rect 105 297 139 2273
rect 223 297 257 2273
rect 341 297 375 2273
rect 459 297 493 2273
rect 577 297 611 2273
rect 695 297 729 2273
rect 813 297 847 2273
rect 931 297 965 2273
rect 1049 297 1083 2273
rect 1167 297 1201 2273
rect 1285 297 1319 2273
rect 1403 297 1437 2273
rect 1521 297 1555 2273
rect 1639 297 1673 2273
rect 1757 297 1791 2273
rect 1875 297 1909 2273
rect 1993 297 2027 2273
rect 2111 297 2145 2273
rect 2229 297 2263 2273
rect 2347 297 2381 2273
rect 2465 297 2499 2273
rect 2583 297 2617 2273
rect 2701 297 2735 2273
rect 2819 297 2853 2273
rect 2937 297 2971 2273
rect 3055 297 3089 2273
rect 3173 297 3207 2273
rect 3291 297 3325 2273
rect 3409 297 3443 2273
rect 3527 297 3561 2273
rect 3645 297 3679 2273
rect 3763 297 3797 2273
rect 3881 297 3915 2273
rect 3999 297 4033 2273
rect 4117 297 4151 2273
rect 4235 297 4269 2273
rect 4353 297 4387 2273
rect 4471 297 4505 2273
rect 4589 297 4623 2273
rect 4707 297 4741 2273
rect 4825 297 4859 2273
rect 4943 297 4977 2273
rect 5061 297 5095 2273
rect 5179 297 5213 2273
rect 5293 1885 5327 2285
rect 5293 285 5327 685
rect 46 204 80 238
rect 164 204 198 238
rect 282 204 316 238
rect 400 204 434 238
rect 518 204 552 238
rect 636 204 670 238
rect 754 204 788 238
rect 872 204 906 238
rect 990 204 1024 238
rect 1108 204 1142 238
rect 1226 204 1260 238
rect 1344 204 1378 238
rect 1462 204 1496 238
rect 1580 204 1614 238
rect 1698 204 1732 238
rect 1816 204 1850 238
rect 1934 204 1968 238
rect 2052 204 2086 238
rect 2170 204 2204 238
rect 2288 204 2322 238
rect 2406 204 2440 238
rect 2524 204 2558 238
rect 2642 204 2676 238
rect 2760 204 2794 238
rect 2878 204 2912 238
rect 2996 204 3030 238
rect 3114 204 3148 238
rect 3232 204 3266 238
rect 3350 204 3384 238
rect 3468 204 3502 238
rect 3586 204 3620 238
rect 3704 204 3738 238
rect 3822 204 3856 238
rect 3940 204 3974 238
rect 4058 204 4092 238
rect 4176 204 4210 238
rect 4294 204 4328 238
rect 4412 204 4446 238
rect 4530 204 4564 238
rect 4648 204 4682 238
rect 4766 204 4800 238
rect 4884 204 4918 238
rect 5002 204 5036 238
rect 5120 204 5154 238
rect 45 -186 79 -152
rect 163 -186 197 -152
rect 281 -186 315 -152
rect 399 -186 433 -152
rect 517 -186 551 -152
rect 635 -186 669 -152
rect 753 -186 787 -152
rect 871 -186 905 -152
rect 989 -186 1023 -152
rect 1107 -186 1141 -152
rect -128 -624 -94 -224
rect -128 -2224 -94 -1824
rect -14 -2212 20 -236
rect 104 -2212 138 -236
rect 222 -2212 256 -236
rect 340 -2212 374 -236
rect 458 -2212 492 -236
rect 576 -2212 610 -236
rect 694 -2212 728 -236
rect 812 -2212 846 -236
rect 930 -2212 964 -236
rect 1048 -2212 1082 -236
rect 1166 -2212 1200 -236
rect 1280 -624 1314 -224
rect 4058 -186 4092 -152
rect 4176 -186 4210 -152
rect 4294 -186 4328 -152
rect 4412 -186 4446 -152
rect 4530 -186 4564 -152
rect 4648 -186 4682 -152
rect 4766 -186 4800 -152
rect 4884 -186 4918 -152
rect 5002 -186 5036 -152
rect 5120 -186 5154 -152
rect 1719 -358 1753 -324
rect 3447 -358 3481 -324
rect 1509 -900 1543 -400
rect 1623 -888 1657 -412
rect 1719 -888 1753 -412
rect 1815 -888 1849 -412
rect 1911 -888 1945 -412
rect 2007 -888 2041 -412
rect 2103 -888 2137 -412
rect 2199 -888 2233 -412
rect 2295 -888 2329 -412
rect 2391 -888 2425 -412
rect 2487 -888 2521 -412
rect 2583 -888 2617 -412
rect 2679 -888 2713 -412
rect 2775 -888 2809 -412
rect 2871 -888 2905 -412
rect 2967 -888 3001 -412
rect 3063 -888 3097 -412
rect 3159 -888 3193 -412
rect 3255 -888 3289 -412
rect 3351 -888 3385 -412
rect 3447 -888 3481 -412
rect 3543 -888 3577 -412
rect 3657 -900 3691 -400
rect 1911 -984 1945 -950
rect 2103 -984 2137 -950
rect 2295 -984 2329 -950
rect 2487 -984 2521 -950
rect 2679 -984 2713 -950
rect 2871 -984 2905 -950
rect 3063 -984 3097 -950
rect 3255 -984 3289 -950
rect 3885 -624 3919 -224
rect 1280 -2224 1314 -1824
rect 45 -2296 79 -2262
rect 163 -2296 197 -2262
rect 281 -2296 315 -2262
rect 399 -2296 433 -2262
rect 517 -2296 551 -2262
rect 635 -2296 669 -2262
rect 753 -2296 787 -2262
rect 871 -2296 905 -2262
rect 989 -2296 1023 -2262
rect 1107 -2296 1141 -2262
rect 1729 -1302 2097 -1268
rect 2187 -1302 2555 -1268
rect 2645 -1302 3013 -1268
rect 3103 -1302 3471 -1268
rect 1553 -1740 1587 -1340
rect 1553 -3340 1587 -2940
rect 1667 -3328 1701 -1352
rect 2125 -3328 2159 -1352
rect 2583 -3328 2617 -1352
rect 3041 -3328 3075 -1352
rect 3499 -3328 3533 -1352
rect 3613 -1740 3647 -1340
rect 3885 -2224 3919 -1824
rect 3999 -2212 4033 -236
rect 4117 -2212 4151 -236
rect 4235 -2212 4269 -236
rect 4353 -2212 4387 -236
rect 4471 -2212 4505 -236
rect 4589 -2212 4623 -236
rect 4707 -2212 4741 -236
rect 4825 -2212 4859 -236
rect 4943 -2212 4977 -236
rect 5061 -2212 5095 -236
rect 5179 -2212 5213 -236
rect 5293 -624 5327 -224
rect 5293 -2224 5327 -1824
rect 4058 -2296 4092 -2262
rect 4176 -2296 4210 -2262
rect 4294 -2296 4328 -2262
rect 4412 -2296 4446 -2262
rect 4530 -2296 4564 -2262
rect 4648 -2296 4682 -2262
rect 4766 -2296 4800 -2262
rect 4884 -2296 4918 -2262
rect 5002 -2296 5036 -2262
rect 5120 -2296 5154 -2262
rect 3613 -3340 3647 -2940
rect 1729 -3412 2097 -3378
rect 2187 -3412 2555 -3378
rect 2645 -3412 3013 -3378
rect 3103 -3412 3471 -3378
<< metal1 >>
rect -22 2366 210 2372
rect -22 2332 46 2366
rect 80 2332 164 2366
rect 198 2332 210 2366
rect -22 2326 210 2332
rect 270 2366 2334 2372
rect 270 2332 282 2366
rect 316 2332 400 2366
rect 434 2332 518 2366
rect 552 2332 636 2366
rect 670 2332 754 2366
rect 788 2332 872 2366
rect 906 2332 990 2366
rect 1024 2332 1108 2366
rect 1142 2332 1226 2366
rect 1260 2332 1344 2366
rect 1378 2332 1462 2366
rect 1496 2332 1580 2366
rect 1614 2332 1698 2366
rect 1732 2332 1816 2366
rect 1850 2332 1934 2366
rect 1968 2332 2052 2366
rect 2086 2332 2170 2366
rect 2204 2332 2288 2366
rect 2322 2332 2334 2366
rect 270 2326 2334 2332
rect 2866 2366 4930 2372
rect 2866 2332 2878 2366
rect 2912 2332 2996 2366
rect 3030 2332 3114 2366
rect 3148 2332 3232 2366
rect 3266 2332 3350 2366
rect 3384 2332 3468 2366
rect 3502 2332 3586 2366
rect 3620 2332 3704 2366
rect 3738 2332 3822 2366
rect 3856 2332 3940 2366
rect 3974 2332 4058 2366
rect 4092 2332 4176 2366
rect 4210 2332 4294 2366
rect 4328 2332 4412 2366
rect 4446 2332 4530 2366
rect 4564 2332 4648 2366
rect 4682 2332 4766 2366
rect 4800 2332 4884 2366
rect 4918 2332 4930 2366
rect 2866 2326 4930 2332
rect 4990 2366 5222 2372
rect 4990 2332 5002 2366
rect 5036 2332 5120 2366
rect 5154 2332 5222 2366
rect 4990 2326 5222 2332
rect -133 2285 -87 2297
rect -22 2285 30 2326
rect -133 1885 -127 2285
rect -93 2273 30 2285
rect -93 1885 -22 2273
rect -133 1873 -87 1885
rect -133 685 -87 697
rect -133 285 -127 685
rect -93 297 -22 685
rect -93 285 30 297
rect -133 273 -87 285
rect -22 244 30 285
rect 96 2273 148 2285
rect 96 244 148 297
rect 214 2273 266 2285
rect 214 285 266 297
rect 332 2273 384 2285
rect 332 285 384 297
rect 450 2273 502 2285
rect 450 285 502 297
rect 568 2273 620 2285
rect 568 285 620 297
rect 686 2273 738 2285
rect 686 285 738 297
rect 804 2273 856 2285
rect 804 285 856 297
rect 922 2273 974 2285
rect 922 285 974 297
rect 1040 2273 1092 2285
rect 1040 285 1092 297
rect 1158 2273 1210 2285
rect 1158 285 1210 297
rect 1276 2273 1328 2285
rect 1276 285 1328 297
rect 1394 2273 1446 2285
rect 1394 285 1446 297
rect 1512 2273 1564 2285
rect 1512 285 1564 297
rect 1630 2273 1682 2285
rect 1630 285 1682 297
rect 1748 2273 1800 2285
rect 1748 285 1800 297
rect 1866 2273 1918 2285
rect 1866 285 1918 297
rect 1984 2273 2036 2285
rect 1984 285 2036 297
rect 2102 2273 2154 2285
rect 2102 285 2154 297
rect 2220 2273 2272 2326
rect 2220 244 2272 297
rect 2338 2273 2390 2285
rect 2338 285 2390 297
rect 2456 2273 2508 2285
rect 2456 285 2508 297
rect 2574 2273 2626 2285
rect 2574 285 2626 297
rect 2692 2273 2744 2285
rect 2692 285 2744 297
rect 2810 2273 2862 2285
rect 2810 285 2862 297
rect 2928 2273 2980 2326
rect 2508 244 2574 250
rect 2928 244 2980 297
rect 3046 2273 3098 2285
rect 3046 285 3098 297
rect 3164 2273 3216 2285
rect 3164 285 3216 297
rect 3282 2273 3334 2285
rect 3282 285 3334 297
rect 3400 2273 3452 2285
rect 3400 285 3452 297
rect 3518 2273 3570 2285
rect 3518 285 3570 297
rect 3636 2273 3688 2285
rect 3636 285 3688 297
rect 3754 2273 3806 2285
rect 3754 285 3806 297
rect 3872 2273 3924 2285
rect 3872 285 3924 297
rect 3990 2273 4042 2285
rect 3990 285 4042 297
rect 4108 2273 4160 2285
rect 4108 285 4160 297
rect 4226 2273 4278 2285
rect 4226 285 4278 297
rect 4344 2273 4396 2285
rect 4344 285 4396 297
rect 4462 2273 4514 2285
rect 4462 285 4514 297
rect 4580 2273 4632 2285
rect 4580 285 4632 297
rect 4698 2273 4750 2285
rect 4698 285 4750 297
rect 4816 2273 4868 2285
rect 4816 285 4868 297
rect 4934 2273 4986 2285
rect 4934 285 4986 297
rect 5052 2273 5104 2326
rect 5052 244 5104 297
rect 5170 2285 5222 2326
rect 5287 2285 5333 2297
rect 5170 2273 5293 2285
rect 5222 1885 5293 2273
rect 5327 1885 5333 2285
rect 5287 1873 5333 1885
rect 5287 685 5333 697
rect 5222 297 5293 685
rect 5170 285 5293 297
rect 5327 285 5333 685
rect 5170 244 5222 285
rect 5287 273 5333 285
rect -22 238 210 244
rect -22 204 46 238
rect 80 204 164 238
rect 198 204 210 238
rect -22 198 210 204
rect 270 238 2338 244
rect 270 204 282 238
rect 316 204 400 238
rect 434 204 518 238
rect 552 204 636 238
rect 670 204 754 238
rect 788 204 872 238
rect 906 204 990 238
rect 1024 204 1108 238
rect 1142 204 1226 238
rect 1260 204 1344 238
rect 1378 204 1462 238
rect 1496 204 1580 238
rect 1614 204 1698 238
rect 1732 204 1816 238
rect 1850 204 1934 238
rect 1968 204 2052 238
rect 2086 204 2170 238
rect 2204 204 2288 238
rect 2322 204 2338 238
rect 270 198 2338 204
rect 2390 238 2512 244
rect 2390 204 2406 238
rect 2440 204 2512 238
rect 2390 198 2512 204
rect 2508 187 2512 198
rect 2571 187 2574 244
rect 2508 181 2574 187
rect 2630 238 2810 244
rect 2630 204 2642 238
rect 2676 204 2760 238
rect 2794 204 2810 238
rect 2630 198 2810 204
rect 2862 238 4930 244
rect 2862 204 2878 238
rect 2912 204 2996 238
rect 3030 204 3114 238
rect 3148 204 3232 238
rect 3266 204 3350 238
rect 3384 204 3468 238
rect 3502 204 3586 238
rect 3620 204 3704 238
rect 3738 204 3822 238
rect 3856 204 3940 238
rect 3974 204 4058 238
rect 4092 204 4176 238
rect 4210 204 4294 238
rect 4328 204 4412 238
rect 4446 204 4530 238
rect 4564 204 4648 238
rect 4682 204 4766 238
rect 4800 204 4884 238
rect 4918 204 4930 238
rect 2862 198 4930 204
rect 4990 238 5222 244
rect 4990 204 5002 238
rect 5036 204 5120 238
rect 5154 204 5222 238
rect 4990 198 5222 204
rect 2630 187 2689 198
rect 2630 124 2689 130
rect 331 -42 383 -36
rect 331 -146 383 -94
rect 567 -42 619 -36
rect 567 -146 619 -94
rect 803 -42 855 -36
rect 803 -146 855 -94
rect 4344 -42 4396 -36
rect 4344 -146 4396 -94
rect 4580 -42 4632 -36
rect 4580 -146 4632 -94
rect 4816 -42 4868 -36
rect 4816 -146 4868 -94
rect -23 -152 91 -146
rect -23 -186 45 -152
rect 79 -186 91 -152
rect -23 -192 91 -186
rect 151 -152 1035 -146
rect 151 -186 163 -152
rect 197 -186 281 -152
rect 315 -186 399 -152
rect 433 -186 517 -152
rect 551 -186 635 -152
rect 669 -186 753 -152
rect 787 -186 871 -152
rect 905 -186 989 -152
rect 1023 -186 1035 -152
rect 151 -192 1035 -186
rect 1095 -152 1209 -146
rect 1095 -186 1107 -152
rect 1141 -186 1209 -152
rect 1095 -192 1209 -186
rect -134 -224 -88 -212
rect -23 -224 29 -192
rect 1157 -224 1209 -192
rect 3990 -152 4104 -146
rect 3990 -186 4058 -152
rect 4092 -186 4104 -152
rect 3990 -192 4104 -186
rect 4164 -152 5048 -146
rect 4164 -186 4176 -152
rect 4210 -186 4294 -152
rect 4328 -186 4412 -152
rect 4446 -186 4530 -152
rect 4564 -186 4648 -152
rect 4682 -186 4766 -152
rect 4800 -186 4884 -152
rect 4918 -186 5002 -152
rect 5036 -186 5048 -152
rect 4164 -192 5048 -186
rect 5108 -152 5222 -146
rect 5108 -186 5120 -152
rect 5154 -186 5222 -152
rect 5108 -192 5222 -186
rect 1300 -212 1400 -200
rect 1274 -224 1400 -212
rect -134 -624 -128 -224
rect -94 -236 29 -224
rect -94 -624 -23 -236
rect -134 -636 -88 -624
rect -134 -1824 -88 -1812
rect -134 -2224 -128 -1824
rect -94 -2212 -23 -1824
rect -94 -2224 29 -2212
rect 95 -236 147 -224
rect 95 -2224 147 -2212
rect 213 -236 265 -224
rect 213 -2224 265 -2212
rect 331 -236 383 -224
rect 331 -2224 383 -2212
rect 449 -236 501 -224
rect 449 -2224 501 -2212
rect 567 -236 619 -224
rect 567 -2224 619 -2212
rect 685 -236 737 -224
rect 685 -2224 737 -2212
rect 803 -236 855 -224
rect 803 -2224 855 -2212
rect 921 -236 973 -224
rect 921 -2224 973 -2212
rect 1039 -236 1091 -224
rect 1039 -2224 1091 -2212
rect 1157 -236 1280 -224
rect 1209 -624 1280 -236
rect 1314 -300 1400 -224
rect 3800 -212 3900 -200
rect 3800 -224 3925 -212
rect 3990 -224 4042 -192
rect 5170 -224 5222 -192
rect 5287 -224 5333 -212
rect 3800 -300 3885 -224
rect 1314 -400 1560 -300
rect 1617 -324 1769 -318
rect 1617 -358 1719 -324
rect 1753 -358 1769 -324
rect 1617 -364 1769 -358
rect 3431 -324 3583 -318
rect 3431 -358 3447 -324
rect 3481 -358 3583 -324
rect 3431 -364 3583 -358
rect 1617 -400 1663 -364
rect 1713 -400 1759 -364
rect 3441 -400 3487 -364
rect 3537 -400 3583 -364
rect 3640 -400 3885 -300
rect 1314 -624 1509 -400
rect 1274 -636 1509 -624
rect 1300 -800 1509 -636
rect 1400 -900 1509 -800
rect 1543 -900 1613 -400
rect 1667 -900 1673 -400
rect 1703 -900 1709 -400
rect 1763 -900 1769 -400
rect 1799 -900 1805 -400
rect 1859 -900 1865 -400
rect 1895 -900 1901 -400
rect 1955 -900 1961 -400
rect 1991 -900 1997 -400
rect 2051 -900 2057 -400
rect 2087 -900 2093 -400
rect 2147 -900 2153 -400
rect 2183 -900 2189 -400
rect 2243 -900 2249 -400
rect 2279 -900 2285 -400
rect 2339 -900 2345 -400
rect 2375 -900 2381 -400
rect 2435 -900 2441 -400
rect 2471 -900 2477 -400
rect 2531 -900 2537 -400
rect 2567 -900 2573 -400
rect 2627 -900 2633 -400
rect 2663 -900 2669 -400
rect 2723 -900 2729 -400
rect 2759 -900 2765 -400
rect 2819 -900 2825 -400
rect 2855 -900 2861 -400
rect 2915 -900 2921 -400
rect 2951 -900 2957 -400
rect 3011 -900 3017 -400
rect 3047 -900 3053 -400
rect 3107 -900 3113 -400
rect 3143 -900 3149 -400
rect 3203 -900 3209 -400
rect 3239 -900 3245 -400
rect 3299 -900 3305 -400
rect 3335 -900 3341 -400
rect 3395 -900 3401 -400
rect 3431 -900 3437 -400
rect 3491 -900 3497 -400
rect 3527 -900 3533 -400
rect 3587 -900 3657 -400
rect 3691 -624 3885 -400
rect 3919 -236 4042 -224
rect 3919 -624 3990 -236
rect 3691 -636 3925 -624
rect 3691 -800 3900 -636
rect 3691 -900 3800 -800
rect 1400 -1200 1560 -900
rect 1889 -1000 1895 -944
rect 1961 -1000 1967 -944
rect 2081 -1000 2087 -944
rect 2153 -1000 2159 -944
rect 2273 -1000 2279 -944
rect 2345 -1000 2351 -944
rect 2465 -1000 2471 -944
rect 2537 -1000 2543 -944
rect 2657 -1000 2663 -944
rect 2729 -1000 2735 -944
rect 2849 -1000 2855 -944
rect 2921 -1000 2927 -944
rect 3041 -1000 3047 -944
rect 3113 -1000 3119 -944
rect 3233 -1000 3239 -944
rect 3305 -1000 3311 -944
rect 1400 -1340 1600 -1200
rect 1717 -1308 1729 -1216
rect 3471 -1308 3483 -1216
rect 3640 -1328 3800 -900
rect 3607 -1340 3800 -1328
rect 1400 -1700 1553 -1340
rect 1300 -1740 1553 -1700
rect 1587 -1352 1710 -1340
rect 1587 -1740 1658 -1352
rect 1300 -1800 1600 -1740
rect 1300 -1812 1560 -1800
rect 1274 -1824 1560 -1812
rect 1209 -2212 1280 -1824
rect 1157 -2224 1280 -2212
rect 1314 -2224 1560 -1824
rect -134 -2236 -88 -2224
rect -23 -2256 29 -2224
rect 1157 -2256 1209 -2224
rect 1274 -2236 1560 -2224
rect -23 -2262 91 -2256
rect -23 -2296 45 -2262
rect 79 -2296 91 -2262
rect -23 -2302 91 -2296
rect 151 -2262 1035 -2256
rect 151 -2296 163 -2262
rect 197 -2296 281 -2262
rect 315 -2296 399 -2262
rect 433 -2296 517 -2262
rect 551 -2296 635 -2262
rect 669 -2296 753 -2262
rect 787 -2296 871 -2262
rect 905 -2296 989 -2262
rect 1023 -2296 1035 -2262
rect 151 -2302 1035 -2296
rect 1095 -2262 1209 -2256
rect 1095 -2296 1107 -2262
rect 1141 -2296 1209 -2262
rect 1095 -2302 1209 -2296
rect 1300 -2300 1560 -2236
rect 1400 -2360 1560 -2300
rect 1400 -3580 1420 -2360
rect 1480 -2928 1560 -2360
rect 1480 -2940 1593 -2928
rect 1480 -3340 1553 -2940
rect 1587 -3328 1658 -2940
rect 1587 -3340 1710 -3328
rect 2116 -1352 2168 -1340
rect 2116 -3340 2168 -3328
rect 2574 -1352 2626 -1340
rect 2574 -3340 2626 -3328
rect 3032 -1352 3084 -1340
rect 3032 -3340 3084 -3328
rect 3490 -1352 3613 -1340
rect 3542 -1740 3613 -1352
rect 3647 -1700 3800 -1340
rect 3647 -1740 3900 -1700
rect 3607 -1752 3900 -1740
rect 3640 -1812 3900 -1752
rect 3640 -1824 3925 -1812
rect 3640 -2224 3885 -1824
rect 3919 -2212 3990 -1824
rect 3919 -2224 4042 -2212
rect 4108 -236 4160 -224
rect 4108 -2224 4160 -2212
rect 4226 -236 4278 -224
rect 4226 -2224 4278 -2212
rect 4344 -236 4396 -224
rect 4344 -2224 4396 -2212
rect 4462 -236 4514 -224
rect 4462 -2224 4514 -2212
rect 4580 -236 4632 -224
rect 4580 -2224 4632 -2212
rect 4698 -236 4750 -224
rect 4698 -2224 4750 -2212
rect 4816 -236 4868 -224
rect 4816 -2224 4868 -2212
rect 4934 -236 4986 -224
rect 4934 -2224 4986 -2212
rect 5052 -236 5104 -224
rect 5052 -2224 5104 -2212
rect 5170 -236 5293 -224
rect 5222 -624 5293 -236
rect 5327 -624 5333 -224
rect 5287 -636 5333 -624
rect 5287 -1824 5333 -1812
rect 5222 -2212 5293 -1824
rect 5170 -2224 5293 -2212
rect 5327 -2224 5333 -1824
rect 3640 -2236 3925 -2224
rect 3640 -2300 3900 -2236
rect 3990 -2256 4042 -2224
rect 5170 -2256 5222 -2224
rect 5287 -2236 5333 -2224
rect 3990 -2262 4104 -2256
rect 3990 -2296 4058 -2262
rect 4092 -2296 4104 -2262
rect 3640 -2360 3800 -2300
rect 3990 -2302 4104 -2296
rect 4164 -2262 5048 -2256
rect 4164 -2296 4176 -2262
rect 4210 -2296 4294 -2262
rect 4328 -2296 4412 -2262
rect 4446 -2296 4530 -2262
rect 4564 -2296 4648 -2262
rect 4682 -2296 4766 -2262
rect 4800 -2296 4884 -2262
rect 4918 -2296 5002 -2262
rect 5036 -2296 5048 -2262
rect 4164 -2302 5048 -2296
rect 5108 -2262 5222 -2256
rect 5108 -2296 5120 -2262
rect 5154 -2296 5222 -2262
rect 5108 -2302 5222 -2296
rect 3640 -2928 3720 -2360
rect 3607 -2940 3720 -2928
rect 3542 -3328 3613 -2940
rect 3490 -3340 3613 -3328
rect 3647 -3340 3720 -2940
rect 1480 -3352 1593 -3340
rect 3607 -3352 3720 -3340
rect 1480 -3580 1560 -3352
rect 1717 -3378 3483 -3372
rect 1717 -3412 1729 -3378
rect 2097 -3412 2187 -3378
rect 2555 -3412 2645 -3378
rect 3013 -3412 3103 -3378
rect 3471 -3412 3483 -3378
rect 1717 -3418 3483 -3412
rect 1400 -3600 1560 -3580
rect 3640 -3580 3720 -3352
rect 3780 -3580 3800 -2360
rect 3640 -3600 3800 -3580
<< via1 >>
rect -22 297 -13 2273
rect -13 297 21 2273
rect 21 297 30 2273
rect 96 297 105 2273
rect 105 297 139 2273
rect 139 297 148 2273
rect 214 297 223 2273
rect 223 297 257 2273
rect 257 297 266 2273
rect 332 297 341 2273
rect 341 297 375 2273
rect 375 297 384 2273
rect 450 297 459 2273
rect 459 297 493 2273
rect 493 297 502 2273
rect 568 297 577 2273
rect 577 297 611 2273
rect 611 297 620 2273
rect 686 297 695 2273
rect 695 297 729 2273
rect 729 297 738 2273
rect 804 297 813 2273
rect 813 297 847 2273
rect 847 297 856 2273
rect 922 297 931 2273
rect 931 297 965 2273
rect 965 297 974 2273
rect 1040 297 1049 2273
rect 1049 297 1083 2273
rect 1083 297 1092 2273
rect 1158 297 1167 2273
rect 1167 297 1201 2273
rect 1201 297 1210 2273
rect 1276 297 1285 2273
rect 1285 297 1319 2273
rect 1319 297 1328 2273
rect 1394 297 1403 2273
rect 1403 297 1437 2273
rect 1437 297 1446 2273
rect 1512 297 1521 2273
rect 1521 297 1555 2273
rect 1555 297 1564 2273
rect 1630 297 1639 2273
rect 1639 297 1673 2273
rect 1673 297 1682 2273
rect 1748 297 1757 2273
rect 1757 297 1791 2273
rect 1791 297 1800 2273
rect 1866 297 1875 2273
rect 1875 297 1909 2273
rect 1909 297 1918 2273
rect 1984 297 1993 2273
rect 1993 297 2027 2273
rect 2027 297 2036 2273
rect 2102 297 2111 2273
rect 2111 297 2145 2273
rect 2145 297 2154 2273
rect 2220 297 2229 2273
rect 2229 297 2263 2273
rect 2263 297 2272 2273
rect 2338 297 2347 2273
rect 2347 297 2381 2273
rect 2381 297 2390 2273
rect 2456 297 2465 2273
rect 2465 297 2499 2273
rect 2499 297 2508 2273
rect 2574 297 2583 2273
rect 2583 297 2617 2273
rect 2617 297 2626 2273
rect 2692 297 2701 2273
rect 2701 297 2735 2273
rect 2735 297 2744 2273
rect 2810 297 2819 2273
rect 2819 297 2853 2273
rect 2853 297 2862 2273
rect 2928 297 2937 2273
rect 2937 297 2971 2273
rect 2971 297 2980 2273
rect 3046 297 3055 2273
rect 3055 297 3089 2273
rect 3089 297 3098 2273
rect 3164 297 3173 2273
rect 3173 297 3207 2273
rect 3207 297 3216 2273
rect 3282 297 3291 2273
rect 3291 297 3325 2273
rect 3325 297 3334 2273
rect 3400 297 3409 2273
rect 3409 297 3443 2273
rect 3443 297 3452 2273
rect 3518 297 3527 2273
rect 3527 297 3561 2273
rect 3561 297 3570 2273
rect 3636 297 3645 2273
rect 3645 297 3679 2273
rect 3679 297 3688 2273
rect 3754 297 3763 2273
rect 3763 297 3797 2273
rect 3797 297 3806 2273
rect 3872 297 3881 2273
rect 3881 297 3915 2273
rect 3915 297 3924 2273
rect 3990 297 3999 2273
rect 3999 297 4033 2273
rect 4033 297 4042 2273
rect 4108 297 4117 2273
rect 4117 297 4151 2273
rect 4151 297 4160 2273
rect 4226 297 4235 2273
rect 4235 297 4269 2273
rect 4269 297 4278 2273
rect 4344 297 4353 2273
rect 4353 297 4387 2273
rect 4387 297 4396 2273
rect 4462 297 4471 2273
rect 4471 297 4505 2273
rect 4505 297 4514 2273
rect 4580 297 4589 2273
rect 4589 297 4623 2273
rect 4623 297 4632 2273
rect 4698 297 4707 2273
rect 4707 297 4741 2273
rect 4741 297 4750 2273
rect 4816 297 4825 2273
rect 4825 297 4859 2273
rect 4859 297 4868 2273
rect 4934 297 4943 2273
rect 4943 297 4977 2273
rect 4977 297 4986 2273
rect 5052 297 5061 2273
rect 5061 297 5095 2273
rect 5095 297 5104 2273
rect 5170 297 5179 2273
rect 5179 297 5213 2273
rect 5213 297 5222 2273
rect 2512 238 2571 244
rect 2512 204 2524 238
rect 2524 204 2558 238
rect 2558 204 2571 238
rect 2512 187 2571 204
rect 2630 130 2689 187
rect 331 -94 383 -42
rect 567 -94 619 -42
rect 803 -94 855 -42
rect 4344 -94 4396 -42
rect 4580 -94 4632 -42
rect 4816 -94 4868 -42
rect -23 -2212 -14 -236
rect -14 -2212 20 -236
rect 20 -2212 29 -236
rect 95 -2212 104 -236
rect 104 -2212 138 -236
rect 138 -2212 147 -236
rect 213 -2212 222 -236
rect 222 -2212 256 -236
rect 256 -2212 265 -236
rect 331 -2212 340 -236
rect 340 -2212 374 -236
rect 374 -2212 383 -236
rect 449 -2212 458 -236
rect 458 -2212 492 -236
rect 492 -2212 501 -236
rect 567 -2212 576 -236
rect 576 -2212 610 -236
rect 610 -2212 619 -236
rect 685 -2212 694 -236
rect 694 -2212 728 -236
rect 728 -2212 737 -236
rect 803 -2212 812 -236
rect 812 -2212 846 -236
rect 846 -2212 855 -236
rect 921 -2212 930 -236
rect 930 -2212 964 -236
rect 964 -2212 973 -236
rect 1039 -2212 1048 -236
rect 1048 -2212 1082 -236
rect 1082 -2212 1091 -236
rect 1157 -2212 1166 -236
rect 1166 -2212 1200 -236
rect 1200 -2212 1209 -236
rect 1613 -412 1667 -400
rect 1613 -888 1623 -412
rect 1623 -888 1657 -412
rect 1657 -888 1667 -412
rect 1613 -900 1667 -888
rect 1709 -412 1763 -400
rect 1709 -888 1719 -412
rect 1719 -888 1753 -412
rect 1753 -888 1763 -412
rect 1709 -900 1763 -888
rect 1805 -412 1859 -400
rect 1805 -888 1815 -412
rect 1815 -888 1849 -412
rect 1849 -888 1859 -412
rect 1805 -900 1859 -888
rect 1901 -412 1955 -400
rect 1901 -888 1911 -412
rect 1911 -888 1945 -412
rect 1945 -888 1955 -412
rect 1901 -900 1955 -888
rect 1997 -412 2051 -400
rect 1997 -888 2007 -412
rect 2007 -888 2041 -412
rect 2041 -888 2051 -412
rect 1997 -900 2051 -888
rect 2093 -412 2147 -400
rect 2093 -888 2103 -412
rect 2103 -888 2137 -412
rect 2137 -888 2147 -412
rect 2093 -900 2147 -888
rect 2189 -412 2243 -400
rect 2189 -888 2199 -412
rect 2199 -888 2233 -412
rect 2233 -888 2243 -412
rect 2189 -900 2243 -888
rect 2285 -412 2339 -400
rect 2285 -888 2295 -412
rect 2295 -888 2329 -412
rect 2329 -888 2339 -412
rect 2285 -900 2339 -888
rect 2381 -412 2435 -400
rect 2381 -888 2391 -412
rect 2391 -888 2425 -412
rect 2425 -888 2435 -412
rect 2381 -900 2435 -888
rect 2477 -412 2531 -400
rect 2477 -888 2487 -412
rect 2487 -888 2521 -412
rect 2521 -888 2531 -412
rect 2477 -900 2531 -888
rect 2573 -412 2627 -400
rect 2573 -888 2583 -412
rect 2583 -888 2617 -412
rect 2617 -888 2627 -412
rect 2573 -900 2627 -888
rect 2669 -412 2723 -400
rect 2669 -888 2679 -412
rect 2679 -888 2713 -412
rect 2713 -888 2723 -412
rect 2669 -900 2723 -888
rect 2765 -412 2819 -400
rect 2765 -888 2775 -412
rect 2775 -888 2809 -412
rect 2809 -888 2819 -412
rect 2765 -900 2819 -888
rect 2861 -412 2915 -400
rect 2861 -888 2871 -412
rect 2871 -888 2905 -412
rect 2905 -888 2915 -412
rect 2861 -900 2915 -888
rect 2957 -412 3011 -400
rect 2957 -888 2967 -412
rect 2967 -888 3001 -412
rect 3001 -888 3011 -412
rect 2957 -900 3011 -888
rect 3053 -412 3107 -400
rect 3053 -888 3063 -412
rect 3063 -888 3097 -412
rect 3097 -888 3107 -412
rect 3053 -900 3107 -888
rect 3149 -412 3203 -400
rect 3149 -888 3159 -412
rect 3159 -888 3193 -412
rect 3193 -888 3203 -412
rect 3149 -900 3203 -888
rect 3245 -412 3299 -400
rect 3245 -888 3255 -412
rect 3255 -888 3289 -412
rect 3289 -888 3299 -412
rect 3245 -900 3299 -888
rect 3341 -412 3395 -400
rect 3341 -888 3351 -412
rect 3351 -888 3385 -412
rect 3385 -888 3395 -412
rect 3341 -900 3395 -888
rect 3437 -412 3491 -400
rect 3437 -888 3447 -412
rect 3447 -888 3481 -412
rect 3481 -888 3491 -412
rect 3437 -900 3491 -888
rect 3533 -412 3587 -400
rect 3533 -888 3543 -412
rect 3543 -888 3577 -412
rect 3577 -888 3587 -412
rect 3533 -900 3587 -888
rect 1895 -950 1961 -944
rect 1895 -984 1911 -950
rect 1911 -984 1945 -950
rect 1945 -984 1961 -950
rect 1895 -1000 1961 -984
rect 2087 -950 2153 -944
rect 2087 -984 2103 -950
rect 2103 -984 2137 -950
rect 2137 -984 2153 -950
rect 2087 -1000 2153 -984
rect 2279 -950 2345 -944
rect 2279 -984 2295 -950
rect 2295 -984 2329 -950
rect 2329 -984 2345 -950
rect 2279 -1000 2345 -984
rect 2471 -950 2537 -944
rect 2471 -984 2487 -950
rect 2487 -984 2521 -950
rect 2521 -984 2537 -950
rect 2471 -1000 2537 -984
rect 2663 -950 2729 -944
rect 2663 -984 2679 -950
rect 2679 -984 2713 -950
rect 2713 -984 2729 -950
rect 2663 -1000 2729 -984
rect 2855 -950 2921 -944
rect 2855 -984 2871 -950
rect 2871 -984 2905 -950
rect 2905 -984 2921 -950
rect 2855 -1000 2921 -984
rect 3047 -950 3113 -944
rect 3047 -984 3063 -950
rect 3063 -984 3097 -950
rect 3097 -984 3113 -950
rect 3047 -1000 3113 -984
rect 3239 -950 3305 -944
rect 3239 -984 3255 -950
rect 3255 -984 3289 -950
rect 3289 -984 3305 -950
rect 3239 -1000 3305 -984
rect 1729 -1268 3471 -1216
rect 1729 -1302 2097 -1268
rect 2097 -1302 2187 -1268
rect 2187 -1302 2555 -1268
rect 2555 -1302 2645 -1268
rect 2645 -1302 3013 -1268
rect 3013 -1302 3103 -1268
rect 3103 -1302 3471 -1268
rect 1729 -1308 3471 -1302
rect 1420 -3580 1480 -2360
rect 1658 -3328 1667 -1352
rect 1667 -3328 1701 -1352
rect 1701 -3328 1710 -1352
rect 2116 -3328 2125 -1352
rect 2125 -3328 2159 -1352
rect 2159 -3328 2168 -1352
rect 2574 -3328 2583 -1352
rect 2583 -3328 2617 -1352
rect 2617 -3328 2626 -1352
rect 3032 -3328 3041 -1352
rect 3041 -3328 3075 -1352
rect 3075 -3328 3084 -1352
rect 3490 -3328 3499 -1352
rect 3499 -3328 3533 -1352
rect 3533 -3328 3542 -1352
rect 3990 -2212 3999 -236
rect 3999 -2212 4033 -236
rect 4033 -2212 4042 -236
rect 4108 -2212 4117 -236
rect 4117 -2212 4151 -236
rect 4151 -2212 4160 -236
rect 4226 -2212 4235 -236
rect 4235 -2212 4269 -236
rect 4269 -2212 4278 -236
rect 4344 -2212 4353 -236
rect 4353 -2212 4387 -236
rect 4387 -2212 4396 -236
rect 4462 -2212 4471 -236
rect 4471 -2212 4505 -236
rect 4505 -2212 4514 -236
rect 4580 -2212 4589 -236
rect 4589 -2212 4623 -236
rect 4623 -2212 4632 -236
rect 4698 -2212 4707 -236
rect 4707 -2212 4741 -236
rect 4741 -2212 4750 -236
rect 4816 -2212 4825 -236
rect 4825 -2212 4859 -236
rect 4859 -2212 4868 -236
rect 4934 -2212 4943 -236
rect 4943 -2212 4977 -236
rect 4977 -2212 4986 -236
rect 5052 -2212 5061 -236
rect 5061 -2212 5095 -236
rect 5095 -2212 5104 -236
rect 5170 -2212 5179 -236
rect 5179 -2212 5213 -236
rect 5213 -2212 5222 -236
rect 3720 -3580 3780 -2360
<< metal2 >>
rect 0 2600 5200 2800
rect 0 2536 100 2600
rect 400 2536 500 2600
rect 800 2536 900 2600
rect 1200 2536 1300 2600
rect 1600 2536 1700 2600
rect 2000 2536 2100 2600
rect 2400 2536 2500 2600
rect 2700 2536 2800 2600
rect 3100 2536 3200 2600
rect 3500 2536 3600 2600
rect 3900 2536 4000 2600
rect 4300 2536 4400 2600
rect 4700 2536 4800 2600
rect 5100 2536 5200 2600
rect -22 2434 5222 2536
rect -22 2273 30 2434
rect -22 285 30 297
rect 96 2273 148 2434
rect 96 285 148 297
rect 214 2273 266 2434
rect 214 285 266 297
rect 332 2273 384 2285
rect 332 136 384 297
rect 450 2273 502 2434
rect 450 285 502 297
rect 568 2273 620 2285
rect 568 136 620 297
rect 686 2273 738 2434
rect 686 285 738 297
rect 804 2273 856 2285
rect 804 136 856 297
rect 922 2273 974 2434
rect 922 285 974 297
rect 1040 2273 1092 2285
rect 1040 136 1092 297
rect 1158 2273 1210 2434
rect 1158 285 1210 297
rect 1276 2273 1328 2285
rect 1276 136 1328 297
rect 1394 2273 1446 2434
rect 1394 285 1446 297
rect 1512 2273 1564 2285
rect 1512 136 1564 297
rect 1630 2273 1682 2434
rect 1630 285 1682 297
rect 1748 2273 1800 2285
rect 1748 136 1800 297
rect 1866 2273 1918 2434
rect 1866 285 1918 297
rect 1984 2273 2036 2285
rect 1984 136 2036 297
rect 2102 2273 2154 2434
rect 2102 285 2154 297
rect 2220 2273 2272 2285
rect 213 34 2036 136
rect 2220 105 2272 297
rect 2338 2273 2390 2434
rect 2338 285 2390 297
rect 2456 2273 2508 2285
rect 2456 281 2508 297
rect 2574 2273 2626 2434
rect 2574 285 2626 297
rect 2692 2273 2744 2285
rect 2692 285 2744 297
rect 2810 2273 2862 2434
rect 2810 285 2862 297
rect 2928 2273 2980 2285
rect 2456 152 2484 281
rect 2715 250 2743 285
rect 2512 244 2743 250
rect 2571 222 2743 244
rect 2571 187 2574 222
rect 2512 181 2574 187
rect 2630 187 2689 193
rect 2456 130 2630 152
rect 2456 124 2689 130
rect 2928 105 2980 297
rect 3046 2273 3098 2434
rect 3164 2273 3216 2285
rect 3046 285 3098 297
rect 3163 297 3164 365
rect 3163 285 3216 297
rect 3282 2273 3334 2434
rect 3400 2273 3452 2285
rect 3282 285 3334 297
rect 3399 297 3400 365
rect 3399 285 3452 297
rect 3518 2273 3570 2434
rect 3636 2273 3688 2285
rect 3518 285 3570 297
rect 3635 297 3636 365
rect 3635 285 3688 297
rect 3754 2273 3806 2434
rect 3872 2273 3924 2285
rect 3754 285 3806 297
rect 3871 297 3872 365
rect 3871 285 3924 297
rect 3990 2273 4042 2434
rect 4108 2273 4160 2285
rect 3990 285 4042 297
rect 4107 297 4108 365
rect 4107 285 4160 297
rect 4226 2273 4278 2434
rect 4344 2273 4396 2285
rect 4226 285 4278 297
rect 4343 297 4344 365
rect 4343 285 4396 297
rect 4462 2273 4514 2434
rect 4580 2273 4632 2285
rect 4462 285 4514 297
rect 4579 297 4580 365
rect 4579 285 4632 297
rect 4698 2273 4750 2434
rect 4816 2273 4868 2285
rect 4698 285 4750 297
rect 4815 297 4816 365
rect 4815 285 4868 297
rect 4934 2273 4986 2434
rect 5052 2273 5104 2434
rect 4934 285 4986 297
rect 5051 297 5052 365
rect 5051 285 5104 297
rect 5170 2273 5222 2434
rect 5170 285 5222 297
rect 213 -31 265 34
rect 449 -31 501 34
rect 685 -31 737 34
rect 921 -31 973 34
rect 213 -40 973 -31
rect 213 -96 329 -40
rect 385 -96 565 -40
rect 621 -96 801 -40
rect 857 -96 973 -40
rect 213 -105 973 -96
rect -23 -236 29 -224
rect -23 -2364 29 -2212
rect 95 -236 147 -224
rect 95 -2364 147 -2212
rect 213 -236 265 -105
rect 213 -2224 265 -2212
rect 331 -236 383 -224
rect 331 -2364 383 -2212
rect 449 -236 501 -105
rect 449 -2224 501 -2212
rect 567 -236 619 -224
rect 567 -2364 619 -2212
rect 685 -236 737 -105
rect 685 -2224 737 -2212
rect 803 -236 855 -224
rect 803 -2364 855 -2212
rect 921 -236 973 -105
rect 2220 -190 2324 105
rect 2876 -190 2980 105
rect 3163 136 3215 285
rect 3399 136 3451 285
rect 3635 136 3687 285
rect 3871 136 3923 285
rect 4107 136 4159 285
rect 4343 136 4395 285
rect 4579 136 4631 285
rect 4815 136 4867 285
rect 3163 34 4986 136
rect 921 -2224 973 -2212
rect 1039 -236 1091 -224
rect 1039 -2340 1091 -2212
rect 1157 -236 1209 -224
rect 1895 -330 2537 -190
rect 1895 -400 1961 -330
rect 2087 -400 2153 -330
rect 2279 -400 2345 -330
rect 2471 -400 2537 -330
rect 2663 -330 3305 -190
rect 2663 -400 2729 -330
rect 2855 -400 2921 -330
rect 3047 -400 3113 -330
rect 3239 -400 3305 -330
rect 3990 -236 4042 -224
rect 1607 -900 1613 -400
rect 1667 -900 1673 -400
rect 1703 -900 1709 -400
rect 1763 -900 1769 -400
rect 1799 -900 1805 -400
rect 1859 -900 1865 -400
rect 1895 -900 1901 -400
rect 1955 -900 1961 -400
rect 1991 -900 1997 -400
rect 2051 -900 2057 -400
rect 2087 -900 2093 -400
rect 2147 -900 2153 -400
rect 2183 -900 2189 -400
rect 2243 -900 2249 -400
rect 2279 -900 2285 -400
rect 2339 -900 2345 -400
rect 2375 -900 2381 -400
rect 2435 -900 2441 -400
rect 2471 -900 2477 -400
rect 2531 -900 2537 -400
rect 2567 -900 2573 -400
rect 2627 -900 2633 -400
rect 2663 -900 2669 -400
rect 2723 -900 2729 -400
rect 2759 -900 2765 -400
rect 2819 -900 2825 -400
rect 2855 -900 2861 -400
rect 2915 -900 2921 -400
rect 2951 -900 2957 -400
rect 3011 -900 3017 -400
rect 3047 -900 3053 -400
rect 3107 -900 3113 -400
rect 3143 -900 3149 -400
rect 3203 -900 3209 -400
rect 3239 -900 3245 -400
rect 3299 -900 3305 -400
rect 3335 -900 3341 -400
rect 3395 -900 3401 -400
rect 3431 -900 3437 -400
rect 3491 -900 3497 -400
rect 3527 -900 3533 -400
rect 3587 -900 3593 -400
rect 1805 -1060 1859 -900
rect 1895 -944 1961 -938
rect 1895 -1020 1961 -1006
rect 1997 -1060 2051 -900
rect 2087 -944 2153 -938
rect 2087 -1020 2153 -1006
rect 2189 -1060 2243 -900
rect 2279 -944 2345 -938
rect 2279 -1020 2345 -1006
rect 2381 -1060 2435 -900
rect 2471 -944 2537 -938
rect 2471 -1020 2537 -1006
rect 2573 -1060 2627 -900
rect 2663 -944 2729 -938
rect 2663 -1020 2729 -1006
rect 2765 -1060 2819 -900
rect 2855 -944 2921 -938
rect 2855 -1020 2921 -1006
rect 2957 -1060 3011 -900
rect 3047 -944 3113 -938
rect 3047 -1020 3113 -1006
rect 3149 -1060 3203 -900
rect 3239 -944 3305 -938
rect 3239 -1020 3305 -1006
rect 3341 -1060 3395 -900
rect 1805 -1130 3395 -1060
rect 1805 -1216 1859 -1130
rect 1997 -1216 2051 -1130
rect 2189 -1216 2243 -1130
rect 2381 -1216 2435 -1130
rect 2573 -1216 2627 -1130
rect 2765 -1216 2819 -1130
rect 2957 -1216 3011 -1130
rect 3149 -1216 3203 -1130
rect 3341 -1216 3395 -1130
rect 1717 -1308 1729 -1216
rect 3471 -1308 3483 -1216
rect 1157 -2340 1209 -2212
rect 1658 -1352 1710 -1340
rect 1039 -2360 1500 -2340
rect 1039 -2364 1420 -2360
rect -23 -2434 1420 -2364
rect 0 -2600 100 -2434
rect 200 -2600 300 -2434
rect 400 -2600 500 -2434
rect 600 -2600 700 -2434
rect 800 -2600 900 -2434
rect 1000 -2440 1420 -2434
rect 1000 -2600 1100 -2440
rect 1200 -2600 1300 -2440
rect 1400 -2600 1420 -2440
rect 0 -2800 1420 -2600
rect 1100 -3100 1300 -2800
rect 1400 -3100 1420 -2800
rect 1100 -3200 1420 -3100
rect 1100 -3500 1300 -3200
rect 1400 -3500 1420 -3200
rect 1100 -3580 1420 -3500
rect 1480 -3500 1500 -2360
rect 1658 -3480 1710 -3328
rect 2116 -1352 2168 -1308
rect 2116 -3340 2168 -3328
rect 2574 -1352 2626 -1340
rect 2574 -3480 2626 -3328
rect 3032 -1352 3084 -1308
rect 3032 -3340 3084 -3328
rect 3490 -1352 3542 -1340
rect 3990 -2340 4042 -2212
rect 4108 -236 4160 -224
rect 4108 -2340 4160 -2212
rect 4226 -236 4278 34
rect 4339 -40 4400 -31
rect 4339 -96 4342 -40
rect 4398 -96 4400 -40
rect 4339 -105 4400 -96
rect 4226 -2224 4278 -2212
rect 4344 -236 4396 -224
rect 3490 -3480 3542 -3328
rect 1658 -3500 3542 -3480
rect 3700 -2360 4160 -2340
rect 3700 -3500 3720 -2360
rect 1480 -3580 3720 -3500
rect 3780 -2364 4160 -2360
rect 4344 -2364 4396 -2212
rect 4462 -236 4514 34
rect 4575 -40 4636 -31
rect 4575 -96 4578 -40
rect 4634 -96 4636 -40
rect 4575 -105 4636 -96
rect 4462 -2224 4514 -2212
rect 4580 -236 4632 -224
rect 4580 -2364 4632 -2212
rect 4698 -236 4750 34
rect 4811 -40 4872 -31
rect 4811 -96 4814 -40
rect 4870 -96 4872 -40
rect 4811 -105 4872 -96
rect 4698 -2224 4750 -2212
rect 4816 -236 4868 -224
rect 4816 -2364 4868 -2212
rect 4934 -236 4986 34
rect 4934 -2224 4986 -2212
rect 5052 -236 5104 -224
rect 5052 -2364 5104 -2212
rect 5170 -236 5222 -224
rect 5170 -2364 5222 -2212
rect 3780 -2434 5222 -2364
rect 3780 -2440 4200 -2434
rect 3780 -2700 3800 -2440
rect 3900 -2600 4000 -2440
rect 4100 -2600 4200 -2440
rect 4300 -2600 4400 -2434
rect 4500 -2600 4600 -2434
rect 4700 -2600 4800 -2434
rect 4900 -2600 5000 -2434
rect 5100 -2600 5200 -2434
rect 3900 -2700 5200 -2600
rect 3780 -2800 5200 -2700
rect 3780 -3100 3800 -2800
rect 3900 -3100 4100 -2800
rect 3780 -3200 4100 -3100
rect 3780 -3500 3800 -3200
rect 3900 -3500 4100 -3200
rect 3780 -3580 4100 -3500
rect 1100 -3800 4100 -3580
<< via2 >>
rect 329 -42 385 -40
rect 329 -94 331 -42
rect 331 -94 383 -42
rect 383 -94 385 -42
rect 329 -96 385 -94
rect 565 -42 621 -40
rect 565 -94 567 -42
rect 567 -94 619 -42
rect 619 -94 621 -42
rect 565 -96 621 -94
rect 801 -42 857 -40
rect 801 -94 803 -42
rect 803 -94 855 -42
rect 855 -94 857 -42
rect 801 -96 857 -94
rect 1895 -1000 1961 -950
rect 1895 -1006 1961 -1000
rect 2087 -1000 2153 -950
rect 2087 -1006 2153 -1000
rect 2279 -1000 2345 -950
rect 2279 -1006 2345 -1000
rect 2471 -1000 2537 -950
rect 2471 -1006 2537 -1000
rect 2663 -1000 2729 -950
rect 2663 -1006 2729 -1000
rect 2855 -1000 2921 -950
rect 2855 -1006 2921 -1000
rect 3047 -1000 3113 -950
rect 3047 -1006 3113 -1000
rect 3239 -1000 3305 -950
rect 3239 -1006 3305 -1000
rect 4342 -42 4398 -40
rect 4342 -94 4344 -42
rect 4344 -94 4396 -42
rect 4396 -94 4398 -42
rect 4342 -96 4398 -94
rect 4578 -42 4634 -40
rect 4578 -94 4580 -42
rect 4580 -94 4632 -42
rect 4632 -94 4634 -42
rect 4578 -96 4634 -94
rect 4814 -42 4870 -40
rect 4814 -94 4816 -42
rect 4816 -94 4868 -42
rect 4868 -94 4870 -42
rect 4814 -96 4870 -94
<< metal3 >>
rect 324 -40 4875 -31
rect 324 -96 329 -40
rect 385 -96 565 -40
rect 621 -96 801 -40
rect 857 -96 4342 -40
rect 4398 -96 4578 -40
rect 4634 -96 4814 -40
rect 4870 -96 4875 -40
rect 324 -105 4875 -96
rect 860 -136 4339 -105
rect 1889 -950 2543 -938
rect 1889 -1006 1895 -950
rect 1961 -1006 2087 -950
rect 2153 -1006 2279 -950
rect 2345 -1006 2471 -950
rect 2537 -1006 2543 -950
rect 1889 -1020 2543 -1006
rect 2657 -950 3311 -938
rect 2657 -1006 2663 -950
rect 2729 -1006 2855 -950
rect 2921 -1006 3047 -950
rect 3113 -1006 3239 -950
rect 3305 -1006 3311 -950
rect 2657 -1020 3311 -1006
<< labels >>
rlabel via1 1740 -1250 1810 -1220 1 VREF
rlabel metal2 4940 -10 4980 30 1 VOP
rlabel metal3 3240 -1010 3300 -950 1 VIP
rlabel metal3 1900 -1010 1960 -950 1 VIN
rlabel metal2 1100 -3700 1300 -3600 1 VLO
rlabel metal2 0 2700 200 2800 1 VHI
rlabel metal3 1534 -108 1588 -64 1 NMIRROR
rlabel metal2 1556 50 1610 94 1 PMIRROR_1
rlabel metal2 2242 -262 2296 -218 1 N1
rlabel metal2 2918 -252 2972 -208 1 N2
<< end >>
