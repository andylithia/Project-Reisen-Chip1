magic
tech sky130B
magscale 1 2
timestamp 1668536381
<< nwell >>
rect 3550 -3954 5992 -2940
<< pwell >>
rect 3582 -4728 5962 -4072
rect 30 -6050 390 -5410
<< nmos >>
rect 3653 -4582 3683 -4182
rect 3749 -4582 3779 -4182
rect 3845 -4582 3875 -4182
rect 3941 -4582 3971 -4182
rect 4037 -4582 4067 -4182
rect 4133 -4582 4163 -4182
rect 4229 -4582 4259 -4182
rect 4325 -4582 4355 -4182
rect 4421 -4582 4451 -4182
rect 4517 -4582 4547 -4182
rect 4613 -4582 4643 -4182
rect 4709 -4582 4739 -4182
rect 4805 -4582 4835 -4182
rect 4901 -4582 4931 -4182
rect 4997 -4582 5027 -4182
rect 5093 -4582 5123 -4182
rect 5189 -4582 5219 -4182
rect 5285 -4582 5315 -4182
rect 5381 -4582 5411 -4182
rect 5477 -4582 5507 -4182
rect 5573 -4582 5603 -4182
rect 5669 -4582 5699 -4182
rect 5765 -4582 5795 -4182
rect 5861 -4582 5891 -4182
rect 100 -5920 130 -5520
rect 196 -5920 226 -5520
rect 292 -5920 322 -5520
<< pmos >>
rect 3653 -3827 3683 -3107
rect 3749 -3827 3779 -3107
rect 3845 -3827 3875 -3107
rect 3941 -3827 3971 -3107
rect 4037 -3827 4067 -3107
rect 4133 -3827 4163 -3107
rect 4229 -3827 4259 -3107
rect 4325 -3827 4355 -3107
rect 4421 -3827 4451 -3107
rect 4517 -3827 4547 -3107
rect 4613 -3827 4643 -3107
rect 4709 -3827 4739 -3107
rect 4805 -3827 4835 -3107
rect 4901 -3827 4931 -3107
rect 4997 -3827 5027 -3107
rect 5093 -3827 5123 -3107
rect 5189 -3827 5219 -3107
rect 5285 -3827 5315 -3107
rect 5381 -3827 5411 -3107
rect 5477 -3827 5507 -3107
rect 5573 -3827 5603 -3107
rect 5669 -3827 5699 -3107
rect 5765 -3827 5795 -3107
rect 5861 -3827 5891 -3107
<< ndiff >>
rect 3591 -4194 3653 -4182
rect 3591 -4570 3603 -4194
rect 3637 -4570 3653 -4194
rect 3591 -4582 3653 -4570
rect 3683 -4194 3749 -4182
rect 3683 -4570 3699 -4194
rect 3733 -4570 3749 -4194
rect 3683 -4582 3749 -4570
rect 3779 -4194 3845 -4182
rect 3779 -4570 3795 -4194
rect 3829 -4570 3845 -4194
rect 3779 -4582 3845 -4570
rect 3875 -4194 3941 -4182
rect 3875 -4570 3891 -4194
rect 3925 -4570 3941 -4194
rect 3875 -4582 3941 -4570
rect 3971 -4194 4037 -4182
rect 3971 -4570 3987 -4194
rect 4021 -4570 4037 -4194
rect 3971 -4582 4037 -4570
rect 4067 -4194 4133 -4182
rect 4067 -4570 4083 -4194
rect 4117 -4570 4133 -4194
rect 4067 -4582 4133 -4570
rect 4163 -4194 4229 -4182
rect 4163 -4570 4179 -4194
rect 4213 -4570 4229 -4194
rect 4163 -4582 4229 -4570
rect 4259 -4194 4325 -4182
rect 4259 -4570 4275 -4194
rect 4309 -4570 4325 -4194
rect 4259 -4582 4325 -4570
rect 4355 -4194 4421 -4182
rect 4355 -4570 4371 -4194
rect 4405 -4570 4421 -4194
rect 4355 -4582 4421 -4570
rect 4451 -4194 4517 -4182
rect 4451 -4570 4467 -4194
rect 4501 -4570 4517 -4194
rect 4451 -4582 4517 -4570
rect 4547 -4194 4613 -4182
rect 4547 -4570 4563 -4194
rect 4597 -4570 4613 -4194
rect 4547 -4582 4613 -4570
rect 4643 -4194 4709 -4182
rect 4643 -4570 4659 -4194
rect 4693 -4570 4709 -4194
rect 4643 -4582 4709 -4570
rect 4739 -4194 4805 -4182
rect 4739 -4570 4755 -4194
rect 4789 -4570 4805 -4194
rect 4739 -4582 4805 -4570
rect 4835 -4194 4901 -4182
rect 4835 -4570 4851 -4194
rect 4885 -4570 4901 -4194
rect 4835 -4582 4901 -4570
rect 4931 -4194 4997 -4182
rect 4931 -4570 4947 -4194
rect 4981 -4570 4997 -4194
rect 4931 -4582 4997 -4570
rect 5027 -4194 5093 -4182
rect 5027 -4570 5043 -4194
rect 5077 -4570 5093 -4194
rect 5027 -4582 5093 -4570
rect 5123 -4194 5189 -4182
rect 5123 -4570 5139 -4194
rect 5173 -4570 5189 -4194
rect 5123 -4582 5189 -4570
rect 5219 -4194 5285 -4182
rect 5219 -4570 5235 -4194
rect 5269 -4570 5285 -4194
rect 5219 -4582 5285 -4570
rect 5315 -4194 5381 -4182
rect 5315 -4570 5331 -4194
rect 5365 -4570 5381 -4194
rect 5315 -4582 5381 -4570
rect 5411 -4194 5477 -4182
rect 5411 -4570 5427 -4194
rect 5461 -4570 5477 -4194
rect 5411 -4582 5477 -4570
rect 5507 -4194 5573 -4182
rect 5507 -4570 5523 -4194
rect 5557 -4570 5573 -4194
rect 5507 -4582 5573 -4570
rect 5603 -4194 5669 -4182
rect 5603 -4570 5619 -4194
rect 5653 -4570 5669 -4194
rect 5603 -4582 5669 -4570
rect 5699 -4194 5765 -4182
rect 5699 -4570 5715 -4194
rect 5749 -4570 5765 -4194
rect 5699 -4582 5765 -4570
rect 5795 -4194 5861 -4182
rect 5795 -4570 5811 -4194
rect 5845 -4570 5861 -4194
rect 5795 -4582 5861 -4570
rect 5891 -4194 5953 -4182
rect 5891 -4570 5907 -4194
rect 5941 -4570 5953 -4194
rect 5891 -4582 5953 -4570
rect 38 -5532 100 -5520
rect 38 -5908 50 -5532
rect 84 -5908 100 -5532
rect 38 -5920 100 -5908
rect 130 -5532 196 -5520
rect 130 -5908 146 -5532
rect 180 -5908 196 -5532
rect 130 -5920 196 -5908
rect 226 -5532 292 -5520
rect 226 -5908 242 -5532
rect 276 -5908 292 -5532
rect 226 -5920 292 -5908
rect 322 -5532 388 -5520
rect 322 -5908 338 -5532
rect 372 -5908 388 -5532
rect 322 -5920 388 -5908
<< pdiff >>
rect 3591 -3119 3653 -3107
rect 3591 -3815 3603 -3119
rect 3637 -3815 3653 -3119
rect 3591 -3827 3653 -3815
rect 3683 -3119 3749 -3107
rect 3683 -3815 3699 -3119
rect 3733 -3815 3749 -3119
rect 3683 -3827 3749 -3815
rect 3779 -3119 3845 -3107
rect 3779 -3815 3795 -3119
rect 3829 -3815 3845 -3119
rect 3779 -3827 3845 -3815
rect 3875 -3119 3941 -3107
rect 3875 -3815 3891 -3119
rect 3925 -3815 3941 -3119
rect 3875 -3827 3941 -3815
rect 3971 -3119 4037 -3107
rect 3971 -3815 3987 -3119
rect 4021 -3815 4037 -3119
rect 3971 -3827 4037 -3815
rect 4067 -3119 4133 -3107
rect 4067 -3815 4083 -3119
rect 4117 -3815 4133 -3119
rect 4067 -3827 4133 -3815
rect 4163 -3119 4229 -3107
rect 4163 -3815 4179 -3119
rect 4213 -3815 4229 -3119
rect 4163 -3827 4229 -3815
rect 4259 -3119 4325 -3107
rect 4259 -3815 4275 -3119
rect 4309 -3815 4325 -3119
rect 4259 -3827 4325 -3815
rect 4355 -3119 4421 -3107
rect 4355 -3815 4371 -3119
rect 4405 -3815 4421 -3119
rect 4355 -3827 4421 -3815
rect 4451 -3119 4517 -3107
rect 4451 -3815 4467 -3119
rect 4501 -3815 4517 -3119
rect 4451 -3827 4517 -3815
rect 4547 -3119 4613 -3107
rect 4547 -3815 4563 -3119
rect 4597 -3815 4613 -3119
rect 4547 -3827 4613 -3815
rect 4643 -3119 4709 -3107
rect 4643 -3815 4659 -3119
rect 4693 -3815 4709 -3119
rect 4643 -3827 4709 -3815
rect 4739 -3119 4805 -3107
rect 4739 -3815 4755 -3119
rect 4789 -3815 4805 -3119
rect 4739 -3827 4805 -3815
rect 4835 -3119 4901 -3107
rect 4835 -3815 4851 -3119
rect 4885 -3815 4901 -3119
rect 4835 -3827 4901 -3815
rect 4931 -3119 4997 -3107
rect 4931 -3815 4947 -3119
rect 4981 -3815 4997 -3119
rect 4931 -3827 4997 -3815
rect 5027 -3119 5093 -3107
rect 5027 -3815 5043 -3119
rect 5077 -3815 5093 -3119
rect 5027 -3827 5093 -3815
rect 5123 -3119 5189 -3107
rect 5123 -3815 5139 -3119
rect 5173 -3815 5189 -3119
rect 5123 -3827 5189 -3815
rect 5219 -3119 5285 -3107
rect 5219 -3815 5235 -3119
rect 5269 -3815 5285 -3119
rect 5219 -3827 5285 -3815
rect 5315 -3119 5381 -3107
rect 5315 -3815 5331 -3119
rect 5365 -3815 5381 -3119
rect 5315 -3827 5381 -3815
rect 5411 -3119 5477 -3107
rect 5411 -3815 5427 -3119
rect 5461 -3815 5477 -3119
rect 5411 -3827 5477 -3815
rect 5507 -3119 5573 -3107
rect 5507 -3815 5523 -3119
rect 5557 -3815 5573 -3119
rect 5507 -3827 5573 -3815
rect 5603 -3119 5669 -3107
rect 5603 -3815 5619 -3119
rect 5653 -3815 5669 -3119
rect 5603 -3827 5669 -3815
rect 5699 -3119 5765 -3107
rect 5699 -3815 5715 -3119
rect 5749 -3815 5765 -3119
rect 5699 -3827 5765 -3815
rect 5795 -3119 5861 -3107
rect 5795 -3815 5811 -3119
rect 5845 -3815 5861 -3119
rect 5795 -3827 5861 -3815
rect 5891 -3119 5953 -3107
rect 5891 -3815 5907 -3119
rect 5941 -3815 5953 -3119
rect 5891 -3827 5953 -3815
<< ndiffc >>
rect 3603 -4570 3637 -4194
rect 3699 -4570 3733 -4194
rect 3795 -4570 3829 -4194
rect 3891 -4570 3925 -4194
rect 3987 -4570 4021 -4194
rect 4083 -4570 4117 -4194
rect 4179 -4570 4213 -4194
rect 4275 -4570 4309 -4194
rect 4371 -4570 4405 -4194
rect 4467 -4570 4501 -4194
rect 4563 -4570 4597 -4194
rect 4659 -4570 4693 -4194
rect 4755 -4570 4789 -4194
rect 4851 -4570 4885 -4194
rect 4947 -4570 4981 -4194
rect 5043 -4570 5077 -4194
rect 5139 -4570 5173 -4194
rect 5235 -4570 5269 -4194
rect 5331 -4570 5365 -4194
rect 5427 -4570 5461 -4194
rect 5523 -4570 5557 -4194
rect 5619 -4570 5653 -4194
rect 5715 -4570 5749 -4194
rect 5811 -4570 5845 -4194
rect 5907 -4570 5941 -4194
rect 50 -5908 84 -5532
rect 146 -5908 180 -5532
rect 242 -5908 276 -5532
rect 338 -5908 372 -5532
<< pdiffc >>
rect 3603 -3815 3637 -3119
rect 3699 -3815 3733 -3119
rect 3795 -3815 3829 -3119
rect 3891 -3815 3925 -3119
rect 3987 -3815 4021 -3119
rect 4083 -3815 4117 -3119
rect 4179 -3815 4213 -3119
rect 4275 -3815 4309 -3119
rect 4371 -3815 4405 -3119
rect 4467 -3815 4501 -3119
rect 4563 -3815 4597 -3119
rect 4659 -3815 4693 -3119
rect 4755 -3815 4789 -3119
rect 4851 -3815 4885 -3119
rect 4947 -3815 4981 -3119
rect 5043 -3815 5077 -3119
rect 5139 -3815 5173 -3119
rect 5235 -3815 5269 -3119
rect 5331 -3815 5365 -3119
rect 5427 -3815 5461 -3119
rect 5523 -3815 5557 -3119
rect 5619 -3815 5653 -3119
rect 5715 -3815 5749 -3119
rect 5811 -3815 5845 -3119
rect 5907 -3815 5941 -3119
<< psubdiff >>
rect 3596 -4712 3696 -4678
rect 5848 -4712 5948 -4678
<< nsubdiff >>
rect 3596 -3010 3696 -2976
rect 5848 -3010 5948 -2976
<< psubdiffcont >>
rect 3696 -4712 5848 -4678
<< nsubdiffcont >>
rect 3696 -3010 5848 -2976
<< poly >>
rect 3653 -3107 3683 -3076
rect 3749 -3107 3779 -3081
rect 3845 -3107 3875 -3076
rect 3941 -3107 3971 -3081
rect 4037 -3107 4067 -3076
rect 4133 -3107 4163 -3081
rect 4229 -3107 4259 -3076
rect 4325 -3107 4355 -3081
rect 4421 -3107 4451 -3076
rect 4517 -3107 4547 -3081
rect 4613 -3107 4643 -3076
rect 4709 -3107 4739 -3081
rect 4805 -3107 4835 -3081
rect 4901 -3107 4931 -3076
rect 4997 -3107 5027 -3081
rect 5093 -3107 5123 -3076
rect 5189 -3107 5219 -3081
rect 5285 -3107 5315 -3076
rect 5381 -3107 5411 -3081
rect 5477 -3107 5507 -3076
rect 5573 -3107 5603 -3081
rect 5669 -3107 5699 -3076
rect 5765 -3107 5795 -3081
rect 5861 -3107 5891 -3076
rect 3653 -3858 3683 -3827
rect 3749 -3858 3779 -3827
rect 3653 -3874 3779 -3858
rect 3653 -3908 3663 -3874
rect 3768 -3908 3779 -3874
rect 3653 -3924 3779 -3908
rect 3845 -3858 3875 -3827
rect 3941 -3858 3971 -3827
rect 3845 -3874 3971 -3858
rect 3845 -3908 3855 -3874
rect 3960 -3908 3971 -3874
rect 3845 -3924 3971 -3908
rect 4037 -3858 4067 -3827
rect 4133 -3858 4163 -3827
rect 4037 -3874 4163 -3858
rect 4037 -3908 4047 -3874
rect 4152 -3908 4163 -3874
rect 4037 -3924 4163 -3908
rect 4229 -3858 4259 -3827
rect 4325 -3858 4355 -3827
rect 4229 -3874 4355 -3858
rect 4229 -3908 4239 -3874
rect 4344 -3908 4355 -3874
rect 4229 -3924 4355 -3908
rect 4421 -3858 4451 -3827
rect 4517 -3858 4547 -3827
rect 4421 -3874 4547 -3858
rect 4421 -3908 4431 -3874
rect 4536 -3908 4547 -3874
rect 4421 -3924 4547 -3908
rect 4613 -3858 4643 -3827
rect 4709 -3858 4739 -3827
rect 4613 -3874 4739 -3858
rect 4613 -3908 4623 -3874
rect 4728 -3908 4739 -3874
rect 4613 -3924 4739 -3908
rect 4805 -3858 4835 -3827
rect 4901 -3858 4931 -3827
rect 4805 -3874 4931 -3858
rect 4805 -3908 4816 -3874
rect 4921 -3908 4931 -3874
rect 4805 -3924 4931 -3908
rect 4997 -3858 5027 -3827
rect 5093 -3858 5123 -3827
rect 4997 -3874 5123 -3858
rect 4997 -3908 5008 -3874
rect 5113 -3908 5123 -3874
rect 4997 -3924 5123 -3908
rect 5189 -3858 5219 -3827
rect 5285 -3858 5315 -3827
rect 5189 -3874 5315 -3858
rect 5189 -3908 5200 -3874
rect 5305 -3908 5315 -3874
rect 5189 -3924 5315 -3908
rect 5381 -3858 5411 -3827
rect 5477 -3858 5507 -3827
rect 5381 -3874 5507 -3858
rect 5381 -3908 5392 -3874
rect 5497 -3908 5507 -3874
rect 5381 -3924 5507 -3908
rect 5573 -3858 5603 -3827
rect 5669 -3858 5699 -3827
rect 5573 -3874 5699 -3858
rect 5573 -3908 5584 -3874
rect 5689 -3908 5699 -3874
rect 5573 -3924 5699 -3908
rect 5765 -3858 5795 -3827
rect 5861 -3858 5891 -3827
rect 5765 -3874 5891 -3858
rect 5765 -3908 5776 -3874
rect 5881 -3908 5891 -3874
rect 5765 -3924 5891 -3908
rect 3653 -4110 3779 -4094
rect 3653 -4144 3663 -4110
rect 3768 -4144 3779 -4110
rect 3653 -4160 3779 -4144
rect 3653 -4182 3683 -4160
rect 3749 -4182 3779 -4160
rect 3845 -4110 3971 -4094
rect 3845 -4144 3855 -4110
rect 3960 -4144 3971 -4110
rect 3845 -4160 3971 -4144
rect 3845 -4182 3875 -4160
rect 3941 -4182 3971 -4160
rect 4037 -4110 4163 -4094
rect 4037 -4144 4047 -4110
rect 4152 -4144 4163 -4110
rect 4037 -4160 4163 -4144
rect 4037 -4182 4067 -4160
rect 4133 -4182 4163 -4160
rect 4229 -4110 4355 -4094
rect 4229 -4144 4239 -4110
rect 4344 -4144 4355 -4110
rect 4229 -4160 4355 -4144
rect 4229 -4182 4259 -4160
rect 4325 -4182 4355 -4160
rect 4421 -4110 4547 -4094
rect 4421 -4144 4431 -4110
rect 4536 -4144 4547 -4110
rect 4421 -4160 4547 -4144
rect 4421 -4182 4451 -4160
rect 4517 -4182 4547 -4160
rect 4613 -4110 4739 -4094
rect 4613 -4144 4623 -4110
rect 4728 -4144 4739 -4110
rect 4613 -4160 4739 -4144
rect 4613 -4182 4643 -4160
rect 4709 -4182 4739 -4160
rect 4805 -4110 4931 -4094
rect 4805 -4144 4816 -4110
rect 4921 -4144 4931 -4110
rect 4805 -4160 4931 -4144
rect 4805 -4182 4835 -4160
rect 4901 -4182 4931 -4160
rect 4997 -4110 5123 -4094
rect 4997 -4144 5008 -4110
rect 5113 -4144 5123 -4110
rect 4997 -4160 5123 -4144
rect 4997 -4182 5027 -4160
rect 5093 -4182 5123 -4160
rect 5189 -4110 5315 -4094
rect 5189 -4144 5200 -4110
rect 5305 -4144 5315 -4110
rect 5189 -4160 5315 -4144
rect 5189 -4182 5219 -4160
rect 5285 -4182 5315 -4160
rect 5381 -4110 5507 -4094
rect 5381 -4144 5392 -4110
rect 5497 -4144 5507 -4110
rect 5381 -4160 5507 -4144
rect 5381 -4182 5411 -4160
rect 5477 -4182 5507 -4160
rect 5573 -4110 5699 -4094
rect 5573 -4144 5584 -4110
rect 5689 -4144 5699 -4110
rect 5573 -4160 5699 -4144
rect 5573 -4182 5603 -4160
rect 5669 -4182 5699 -4160
rect 5765 -4110 5891 -4094
rect 5765 -4144 5776 -4110
rect 5881 -4144 5891 -4110
rect 5765 -4160 5891 -4144
rect 5765 -4182 5795 -4160
rect 5861 -4182 5891 -4160
rect 3653 -4608 3683 -4582
rect 3749 -4608 3779 -4582
rect 3845 -4608 3875 -4582
rect 3941 -4608 3971 -4582
rect 4037 -4608 4067 -4582
rect 4133 -4608 4163 -4582
rect 4229 -4608 4259 -4582
rect 4325 -4608 4355 -4582
rect 4421 -4608 4451 -4582
rect 4517 -4608 4547 -4582
rect 4613 -4608 4643 -4582
rect 4709 -4608 4739 -4582
rect 4805 -4608 4835 -4582
rect 4901 -4608 4931 -4582
rect 4997 -4608 5027 -4582
rect 5093 -4608 5123 -4582
rect 5189 -4608 5219 -4582
rect 5285 -4608 5315 -4582
rect 5381 -4608 5411 -4582
rect 5477 -4608 5507 -4582
rect 5573 -4608 5603 -4582
rect 5669 -4608 5699 -4582
rect 5765 -4608 5795 -4582
rect 5861 -4608 5891 -4582
rect 100 -5448 226 -5432
rect 100 -5482 110 -5448
rect 215 -5482 226 -5448
rect 100 -5498 226 -5482
rect 100 -5520 130 -5498
rect 196 -5520 226 -5498
rect 292 -5520 322 -5494
rect 100 -5946 130 -5920
rect 196 -5946 226 -5920
rect 292 -5942 322 -5920
rect 274 -6008 340 -5942
<< polycont >>
rect 3663 -3908 3768 -3874
rect 3855 -3908 3960 -3874
rect 4047 -3908 4152 -3874
rect 4239 -3908 4344 -3874
rect 4431 -3908 4536 -3874
rect 4623 -3908 4728 -3874
rect 4816 -3908 4921 -3874
rect 5008 -3908 5113 -3874
rect 5200 -3908 5305 -3874
rect 5392 -3908 5497 -3874
rect 5584 -3908 5689 -3874
rect 5776 -3908 5881 -3874
rect 3663 -4144 3768 -4110
rect 3855 -4144 3960 -4110
rect 4047 -4144 4152 -4110
rect 4239 -4144 4344 -4110
rect 4431 -4144 4536 -4110
rect 4623 -4144 4728 -4110
rect 4816 -4144 4921 -4110
rect 5008 -4144 5113 -4110
rect 5200 -4144 5305 -4110
rect 5392 -4144 5497 -4110
rect 5584 -4144 5689 -4110
rect 5776 -4144 5881 -4110
rect 110 -5482 215 -5448
<< locali >>
rect 3596 -3010 3696 -2976
rect 5848 -3010 5948 -2976
rect 3603 -3119 3637 -3103
rect 3603 -3831 3637 -3815
rect 3699 -3119 3733 -3103
rect 3699 -3831 3733 -3815
rect 3795 -3119 3829 -3103
rect 3795 -3831 3829 -3815
rect 3891 -3119 3925 -3103
rect 3891 -3831 3925 -3815
rect 3987 -3119 4021 -3103
rect 3987 -3831 4021 -3815
rect 4083 -3119 4117 -3103
rect 4083 -3831 4117 -3815
rect 4179 -3119 4213 -3103
rect 4179 -3831 4213 -3815
rect 4275 -3119 4309 -3103
rect 4275 -3831 4309 -3815
rect 4371 -3119 4405 -3103
rect 4371 -3831 4405 -3815
rect 4467 -3119 4501 -3103
rect 4467 -3831 4501 -3815
rect 4563 -3119 4597 -3103
rect 4563 -3831 4597 -3815
rect 4659 -3119 4693 -3103
rect 4659 -3831 4693 -3815
rect 4755 -3119 4789 -3103
rect 4755 -3831 4789 -3815
rect 4851 -3119 4885 -3103
rect 4851 -3831 4885 -3815
rect 4947 -3119 4981 -3103
rect 4947 -3831 4981 -3815
rect 5043 -3119 5077 -3103
rect 5043 -3831 5077 -3815
rect 5139 -3119 5173 -3103
rect 5139 -3831 5173 -3815
rect 5235 -3119 5269 -3103
rect 5235 -3831 5269 -3815
rect 5331 -3119 5365 -3103
rect 5331 -3831 5365 -3815
rect 5427 -3119 5461 -3103
rect 5427 -3831 5461 -3815
rect 5523 -3119 5557 -3103
rect 5523 -3831 5557 -3815
rect 5619 -3119 5653 -3103
rect 5619 -3831 5653 -3815
rect 5715 -3119 5749 -3103
rect 5715 -3831 5749 -3815
rect 5811 -3119 5845 -3103
rect 5811 -3831 5845 -3815
rect 5907 -3119 5941 -3103
rect 5907 -3831 5941 -3815
rect 3647 -3908 3663 -3874
rect 3768 -3908 3784 -3874
rect 3839 -3908 3855 -3874
rect 3960 -3908 3976 -3874
rect 4031 -3908 4047 -3874
rect 4152 -3908 4168 -3874
rect 4223 -3908 4239 -3874
rect 4344 -3908 4360 -3874
rect 4415 -3908 4431 -3874
rect 4536 -3908 4552 -3874
rect 4607 -3908 4623 -3874
rect 4728 -3908 4744 -3874
rect 4800 -3908 4816 -3874
rect 4921 -3908 4937 -3874
rect 4992 -3908 5008 -3874
rect 5113 -3908 5129 -3874
rect 5184 -3908 5200 -3874
rect 5305 -3908 5321 -3874
rect 5376 -3908 5392 -3874
rect 5497 -3908 5513 -3874
rect 5568 -3908 5584 -3874
rect 5689 -3908 5705 -3874
rect 5760 -3908 5776 -3874
rect 5881 -3908 5897 -3874
rect 3686 -3914 3698 -3908
rect 3732 -3914 3744 -3908
rect 3686 -3952 3744 -3914
rect 3686 -3986 3698 -3952
rect 3732 -3986 3744 -3952
rect 3686 -3992 3744 -3986
rect 3878 -3914 3890 -3908
rect 3924 -3914 3936 -3908
rect 3878 -3952 3936 -3914
rect 3878 -3986 3890 -3952
rect 3924 -3986 3936 -3952
rect 3878 -3992 3936 -3986
rect 4070 -3914 4082 -3908
rect 4116 -3914 4128 -3908
rect 4070 -3952 4128 -3914
rect 4070 -3986 4082 -3952
rect 4116 -3986 4128 -3952
rect 4070 -3992 4128 -3986
rect 4262 -3914 4274 -3908
rect 4308 -3914 4320 -3908
rect 4262 -3952 4320 -3914
rect 4262 -3986 4274 -3952
rect 4308 -3986 4320 -3952
rect 4262 -3992 4320 -3986
rect 4454 -3914 4466 -3908
rect 4500 -3914 4512 -3908
rect 4454 -3952 4512 -3914
rect 4454 -3986 4466 -3952
rect 4500 -3986 4512 -3952
rect 4454 -3992 4512 -3986
rect 4646 -3914 4658 -3908
rect 4692 -3914 4704 -3908
rect 4646 -3952 4704 -3914
rect 4646 -3986 4658 -3952
rect 4692 -3986 4704 -3952
rect 4646 -3992 4704 -3986
rect 4840 -3914 4852 -3908
rect 4886 -3914 4898 -3908
rect 4840 -3952 4898 -3914
rect 4840 -3986 4852 -3952
rect 4886 -3986 4898 -3952
rect 4840 -3992 4898 -3986
rect 5032 -3914 5044 -3908
rect 5078 -3914 5090 -3908
rect 5032 -3952 5090 -3914
rect 5032 -3986 5044 -3952
rect 5078 -3986 5090 -3952
rect 5032 -3992 5090 -3986
rect 5224 -3914 5236 -3908
rect 5270 -3914 5282 -3908
rect 5224 -3952 5282 -3914
rect 5224 -3986 5236 -3952
rect 5270 -3986 5282 -3952
rect 5224 -3992 5282 -3986
rect 5416 -3914 5428 -3908
rect 5462 -3914 5474 -3908
rect 5416 -3952 5474 -3914
rect 5416 -3986 5428 -3952
rect 5462 -3986 5474 -3952
rect 5416 -3992 5474 -3986
rect 5608 -3914 5620 -3908
rect 5654 -3914 5666 -3908
rect 5608 -3952 5666 -3914
rect 5608 -3986 5620 -3952
rect 5654 -3986 5666 -3952
rect 5608 -3992 5666 -3986
rect 5800 -3914 5812 -3908
rect 5846 -3914 5858 -3908
rect 5800 -3952 5858 -3914
rect 5800 -3986 5812 -3952
rect 5846 -3986 5858 -3952
rect 5800 -3992 5858 -3986
rect 3686 -4032 3744 -4026
rect 3686 -4066 3698 -4032
rect 3732 -4066 3744 -4032
rect 3686 -4104 3744 -4066
rect 3686 -4110 3698 -4104
rect 3732 -4110 3744 -4104
rect 3878 -4032 3936 -4026
rect 3878 -4066 3890 -4032
rect 3924 -4066 3936 -4032
rect 3878 -4104 3936 -4066
rect 3878 -4110 3890 -4104
rect 3924 -4110 3936 -4104
rect 4070 -4032 4128 -4026
rect 4070 -4066 4082 -4032
rect 4116 -4066 4128 -4032
rect 4070 -4104 4128 -4066
rect 4070 -4110 4082 -4104
rect 4116 -4110 4128 -4104
rect 4262 -4032 4320 -4026
rect 4262 -4066 4274 -4032
rect 4308 -4066 4320 -4032
rect 4262 -4104 4320 -4066
rect 4262 -4110 4274 -4104
rect 4308 -4110 4320 -4104
rect 4454 -4032 4512 -4026
rect 4454 -4066 4466 -4032
rect 4500 -4066 4512 -4032
rect 4454 -4104 4512 -4066
rect 4454 -4110 4466 -4104
rect 4500 -4110 4512 -4104
rect 4646 -4032 4704 -4026
rect 4646 -4066 4658 -4032
rect 4692 -4066 4704 -4032
rect 4646 -4104 4704 -4066
rect 4646 -4110 4658 -4104
rect 4692 -4110 4704 -4104
rect 4840 -4032 4898 -4026
rect 4840 -4066 4852 -4032
rect 4886 -4066 4898 -4032
rect 4840 -4104 4898 -4066
rect 4840 -4110 4852 -4104
rect 4886 -4110 4898 -4104
rect 5032 -4032 5090 -4026
rect 5032 -4066 5044 -4032
rect 5078 -4066 5090 -4032
rect 5032 -4104 5090 -4066
rect 5032 -4110 5044 -4104
rect 5078 -4110 5090 -4104
rect 5224 -4032 5282 -4026
rect 5224 -4066 5236 -4032
rect 5270 -4066 5282 -4032
rect 5224 -4104 5282 -4066
rect 5224 -4110 5236 -4104
rect 5270 -4110 5282 -4104
rect 5416 -4032 5474 -4026
rect 5416 -4066 5428 -4032
rect 5462 -4066 5474 -4032
rect 5416 -4104 5474 -4066
rect 5416 -4110 5428 -4104
rect 5462 -4110 5474 -4104
rect 5608 -4032 5666 -4026
rect 5608 -4066 5620 -4032
rect 5654 -4066 5666 -4032
rect 5608 -4104 5666 -4066
rect 5608 -4110 5620 -4104
rect 5654 -4110 5666 -4104
rect 5800 -4032 5858 -4026
rect 5800 -4066 5812 -4032
rect 5846 -4066 5858 -4032
rect 5800 -4104 5858 -4066
rect 5800 -4110 5812 -4104
rect 5846 -4110 5858 -4104
rect 3647 -4144 3663 -4110
rect 3768 -4144 3784 -4110
rect 3839 -4144 3855 -4110
rect 3960 -4144 3976 -4110
rect 4031 -4144 4047 -4110
rect 4152 -4144 4168 -4110
rect 4223 -4144 4239 -4110
rect 4344 -4144 4360 -4110
rect 4415 -4144 4431 -4110
rect 4536 -4144 4552 -4110
rect 4607 -4144 4623 -4110
rect 4728 -4144 4744 -4110
rect 4800 -4144 4816 -4110
rect 4921 -4144 4937 -4110
rect 4992 -4144 5008 -4110
rect 5113 -4144 5129 -4110
rect 5184 -4144 5200 -4110
rect 5305 -4144 5321 -4110
rect 5376 -4144 5392 -4110
rect 5497 -4144 5513 -4110
rect 5568 -4144 5584 -4110
rect 5689 -4144 5705 -4110
rect 5760 -4144 5776 -4110
rect 5881 -4144 5897 -4110
rect 3603 -4194 3637 -4178
rect 3603 -4586 3637 -4570
rect 3699 -4194 3733 -4178
rect 3699 -4586 3733 -4570
rect 3795 -4194 3829 -4178
rect 3795 -4586 3829 -4570
rect 3891 -4194 3925 -4178
rect 3891 -4586 3925 -4570
rect 3987 -4194 4021 -4178
rect 3987 -4586 4021 -4570
rect 4083 -4194 4117 -4178
rect 4083 -4586 4117 -4570
rect 4179 -4194 4213 -4178
rect 4179 -4586 4213 -4570
rect 4275 -4194 4309 -4178
rect 4275 -4586 4309 -4570
rect 4371 -4194 4405 -4178
rect 4371 -4586 4405 -4570
rect 4467 -4194 4501 -4178
rect 4467 -4586 4501 -4570
rect 4563 -4194 4597 -4178
rect 4563 -4586 4597 -4570
rect 4659 -4194 4693 -4178
rect 4659 -4586 4693 -4570
rect 4755 -4194 4789 -4178
rect 4755 -4586 4789 -4570
rect 4851 -4194 4885 -4178
rect 4851 -4586 4885 -4570
rect 4947 -4194 4981 -4178
rect 4947 -4586 4981 -4570
rect 5043 -4194 5077 -4178
rect 5043 -4586 5077 -4570
rect 5139 -4194 5173 -4178
rect 5139 -4586 5173 -4570
rect 5235 -4194 5269 -4178
rect 5235 -4586 5269 -4570
rect 5331 -4194 5365 -4178
rect 5331 -4586 5365 -4570
rect 5427 -4194 5461 -4178
rect 5427 -4586 5461 -4570
rect 5523 -4194 5557 -4178
rect 5523 -4586 5557 -4570
rect 5619 -4194 5653 -4178
rect 5619 -4586 5653 -4570
rect 5715 -4194 5749 -4178
rect 5715 -4586 5749 -4570
rect 5811 -4194 5845 -4178
rect 5811 -4586 5845 -4570
rect 5907 -4194 5941 -4178
rect 5907 -4586 5941 -4570
rect 3596 -4712 3696 -4678
rect 5848 -4712 5948 -4678
rect 133 -5370 191 -5364
rect 133 -5404 145 -5370
rect 179 -5404 191 -5370
rect 133 -5442 191 -5404
rect 133 -5448 145 -5442
rect 179 -5448 191 -5442
rect 94 -5482 110 -5448
rect 215 -5482 231 -5448
rect 50 -5532 84 -5516
rect 50 -5924 84 -5908
rect 146 -5532 180 -5516
rect 146 -5924 180 -5908
rect 242 -5532 276 -5516
rect 242 -5924 276 -5908
rect 338 -5532 372 -5516
rect 338 -5924 372 -5908
<< viali >>
rect 3696 -3010 5848 -2976
rect 3603 -3815 3637 -3119
rect 3699 -3815 3733 -3119
rect 3795 -3815 3829 -3119
rect 3891 -3815 3925 -3119
rect 3987 -3815 4021 -3119
rect 4083 -3815 4117 -3119
rect 4179 -3815 4213 -3119
rect 4275 -3815 4309 -3119
rect 4371 -3815 4405 -3119
rect 4467 -3815 4501 -3119
rect 4563 -3815 4597 -3119
rect 4659 -3815 4693 -3119
rect 4755 -3815 4789 -3119
rect 4851 -3815 4885 -3119
rect 4947 -3815 4981 -3119
rect 5043 -3815 5077 -3119
rect 5139 -3815 5173 -3119
rect 5235 -3815 5269 -3119
rect 5331 -3815 5365 -3119
rect 5427 -3815 5461 -3119
rect 5523 -3815 5557 -3119
rect 5619 -3815 5653 -3119
rect 5715 -3815 5749 -3119
rect 5811 -3815 5845 -3119
rect 5907 -3815 5941 -3119
rect 3698 -3908 3732 -3880
rect 3890 -3908 3924 -3880
rect 4082 -3908 4116 -3880
rect 4274 -3908 4308 -3880
rect 4466 -3908 4500 -3880
rect 4658 -3908 4692 -3880
rect 4852 -3908 4886 -3880
rect 5044 -3908 5078 -3880
rect 5236 -3908 5270 -3880
rect 5428 -3908 5462 -3880
rect 5620 -3908 5654 -3880
rect 5812 -3908 5846 -3880
rect 3698 -3914 3732 -3908
rect 3698 -3986 3732 -3952
rect 3890 -3914 3924 -3908
rect 3890 -3986 3924 -3952
rect 4082 -3914 4116 -3908
rect 4082 -3986 4116 -3952
rect 4274 -3914 4308 -3908
rect 4274 -3986 4308 -3952
rect 4466 -3914 4500 -3908
rect 4466 -3986 4500 -3952
rect 4658 -3914 4692 -3908
rect 4658 -3986 4692 -3952
rect 4852 -3914 4886 -3908
rect 4852 -3986 4886 -3952
rect 5044 -3914 5078 -3908
rect 5044 -3986 5078 -3952
rect 5236 -3914 5270 -3908
rect 5236 -3986 5270 -3952
rect 5428 -3914 5462 -3908
rect 5428 -3986 5462 -3952
rect 5620 -3914 5654 -3908
rect 5620 -3986 5654 -3952
rect 5812 -3914 5846 -3908
rect 5812 -3986 5846 -3952
rect 3698 -4066 3732 -4032
rect 3698 -4110 3732 -4104
rect 3890 -4066 3924 -4032
rect 3890 -4110 3924 -4104
rect 4082 -4066 4116 -4032
rect 4082 -4110 4116 -4104
rect 4274 -4066 4308 -4032
rect 4274 -4110 4308 -4104
rect 4466 -4066 4500 -4032
rect 4466 -4110 4500 -4104
rect 4658 -4066 4692 -4032
rect 4658 -4110 4692 -4104
rect 4852 -4066 4886 -4032
rect 4852 -4110 4886 -4104
rect 5044 -4066 5078 -4032
rect 5044 -4110 5078 -4104
rect 5236 -4066 5270 -4032
rect 5236 -4110 5270 -4104
rect 5428 -4066 5462 -4032
rect 5428 -4110 5462 -4104
rect 5620 -4066 5654 -4032
rect 5620 -4110 5654 -4104
rect 5812 -4066 5846 -4032
rect 5812 -4110 5846 -4104
rect 3698 -4138 3732 -4110
rect 3890 -4138 3924 -4110
rect 4082 -4138 4116 -4110
rect 4274 -4138 4308 -4110
rect 4466 -4138 4500 -4110
rect 4658 -4138 4692 -4110
rect 4852 -4138 4886 -4110
rect 5044 -4138 5078 -4110
rect 5236 -4138 5270 -4110
rect 5428 -4138 5462 -4110
rect 5620 -4138 5654 -4110
rect 5812 -4138 5846 -4110
rect 3603 -4570 3637 -4194
rect 3699 -4570 3733 -4194
rect 3795 -4570 3829 -4194
rect 3891 -4570 3925 -4194
rect 3987 -4570 4021 -4194
rect 4083 -4570 4117 -4194
rect 4179 -4570 4213 -4194
rect 4275 -4570 4309 -4194
rect 4371 -4570 4405 -4194
rect 4467 -4570 4501 -4194
rect 4563 -4570 4597 -4194
rect 4659 -4570 4693 -4194
rect 4755 -4570 4789 -4194
rect 4851 -4570 4885 -4194
rect 4947 -4570 4981 -4194
rect 5043 -4570 5077 -4194
rect 5139 -4570 5173 -4194
rect 5235 -4570 5269 -4194
rect 5331 -4570 5365 -4194
rect 5427 -4570 5461 -4194
rect 5523 -4570 5557 -4194
rect 5619 -4570 5653 -4194
rect 5715 -4570 5749 -4194
rect 5811 -4570 5845 -4194
rect 5907 -4570 5941 -4194
rect 3696 -4712 5848 -4678
rect 145 -5404 179 -5370
rect 145 -5448 179 -5442
rect 145 -5476 179 -5448
rect 50 -5908 84 -5532
rect 146 -5908 180 -5532
rect 242 -5908 276 -5532
rect 338 -5908 372 -5532
<< metal1 >>
rect 3596 -2976 5948 -2940
rect 3596 -3010 3696 -2976
rect 5848 -3010 5948 -2976
rect 3596 -3040 5948 -3010
rect 3596 -3119 3644 -3040
rect 3596 -3815 3603 -3119
rect 3637 -3815 3644 -3119
rect 3596 -3828 3644 -3815
rect 3693 -3119 3739 -3107
rect 3693 -3815 3699 -3119
rect 3733 -3815 3739 -3119
rect 3693 -3827 3739 -3815
rect 3788 -3119 3836 -3040
rect 3788 -3815 3795 -3119
rect 3829 -3815 3836 -3119
rect 3788 -3828 3836 -3815
rect 3885 -3119 3931 -3107
rect 3885 -3815 3891 -3119
rect 3925 -3815 3931 -3119
rect 3885 -3827 3931 -3815
rect 3980 -3119 4028 -3040
rect 3980 -3815 3987 -3119
rect 4021 -3815 4028 -3119
rect 3980 -3828 4028 -3815
rect 4077 -3119 4123 -3107
rect 4077 -3815 4083 -3119
rect 4117 -3815 4123 -3119
rect 4077 -3827 4123 -3815
rect 4172 -3119 4220 -3040
rect 4172 -3815 4179 -3119
rect 4213 -3815 4220 -3119
rect 4172 -3828 4220 -3815
rect 4269 -3119 4315 -3107
rect 4269 -3815 4275 -3119
rect 4309 -3815 4315 -3119
rect 4269 -3827 4315 -3815
rect 4364 -3119 4412 -3040
rect 4364 -3815 4371 -3119
rect 4405 -3815 4412 -3119
rect 4364 -3828 4412 -3815
rect 4461 -3119 4507 -3107
rect 4461 -3815 4467 -3119
rect 4501 -3815 4507 -3119
rect 4461 -3827 4507 -3815
rect 4556 -3119 4604 -3040
rect 4556 -3815 4563 -3119
rect 4597 -3815 4604 -3119
rect 4556 -3828 4604 -3815
rect 4653 -3119 4699 -3107
rect 4653 -3815 4659 -3119
rect 4693 -3815 4699 -3119
rect 4653 -3827 4699 -3815
rect 4748 -3119 4796 -3040
rect 4748 -3815 4755 -3119
rect 4789 -3815 4796 -3119
rect 4748 -3828 4796 -3815
rect 4845 -3119 4891 -3107
rect 4845 -3815 4851 -3119
rect 4885 -3815 4891 -3119
rect 4845 -3827 4891 -3815
rect 4940 -3119 4988 -3040
rect 4940 -3815 4947 -3119
rect 4981 -3815 4988 -3119
rect 4940 -3828 4988 -3815
rect 5037 -3119 5083 -3107
rect 5037 -3815 5043 -3119
rect 5077 -3815 5083 -3119
rect 5037 -3827 5083 -3815
rect 5132 -3119 5180 -3040
rect 5132 -3815 5139 -3119
rect 5173 -3815 5180 -3119
rect 5132 -3828 5180 -3815
rect 5229 -3119 5275 -3107
rect 5229 -3815 5235 -3119
rect 5269 -3815 5275 -3119
rect 5229 -3827 5275 -3815
rect 5324 -3119 5372 -3040
rect 5324 -3815 5331 -3119
rect 5365 -3815 5372 -3119
rect 5324 -3828 5372 -3815
rect 5421 -3119 5467 -3107
rect 5421 -3815 5427 -3119
rect 5461 -3815 5467 -3119
rect 5421 -3827 5467 -3815
rect 5516 -3119 5564 -3040
rect 5516 -3815 5523 -3119
rect 5557 -3815 5564 -3119
rect 5516 -3828 5564 -3815
rect 5613 -3119 5659 -3107
rect 5613 -3815 5619 -3119
rect 5653 -3815 5659 -3119
rect 5613 -3827 5659 -3815
rect 5708 -3119 5756 -3040
rect 5708 -3815 5715 -3119
rect 5749 -3815 5756 -3119
rect 5708 -3828 5756 -3815
rect 5805 -3119 5851 -3107
rect 5805 -3815 5811 -3119
rect 5845 -3815 5851 -3119
rect 5805 -3827 5851 -3815
rect 5900 -3119 5948 -3040
rect 5900 -3815 5907 -3119
rect 5941 -3815 5948 -3119
rect 5900 -3828 5948 -3815
rect 3686 -3880 3744 -3874
rect 3686 -3914 3698 -3880
rect 3732 -3914 3744 -3880
rect 3686 -3952 3744 -3914
rect 3878 -3880 3936 -3874
rect 3878 -3914 3890 -3880
rect 3924 -3914 3936 -3880
rect 3878 -3952 3936 -3914
rect 4070 -3880 4128 -3874
rect 4070 -3914 4082 -3880
rect 4116 -3914 4128 -3880
rect 4070 -3952 4128 -3914
rect 4262 -3880 4320 -3874
rect 4262 -3914 4274 -3880
rect 4308 -3914 4320 -3880
rect 4262 -3952 4320 -3914
rect 3686 -3986 3698 -3952
rect 3732 -3986 3890 -3952
rect 3924 -3986 4082 -3952
rect 4116 -3986 4274 -3952
rect 4308 -3986 4320 -3952
rect 3686 -4032 4320 -3986
rect 3686 -4066 3698 -4032
rect 3732 -4066 3890 -4032
rect 3924 -4066 4082 -4032
rect 4116 -4066 4274 -4032
rect 4308 -4066 4320 -4032
rect 3686 -4104 3744 -4066
rect 3686 -4138 3698 -4104
rect 3732 -4138 3744 -4104
rect 3686 -4144 3744 -4138
rect 3878 -4104 3936 -4066
rect 3878 -4138 3890 -4104
rect 3924 -4138 3936 -4104
rect 3878 -4144 3936 -4138
rect 4070 -4104 4128 -4066
rect 4070 -4138 4082 -4104
rect 4116 -4138 4128 -4104
rect 4070 -4144 4128 -4138
rect 4262 -4104 4320 -4066
rect 4262 -4138 4274 -4104
rect 4308 -4138 4320 -4104
rect 4262 -4144 4320 -4138
rect 4454 -3880 4512 -3874
rect 4454 -3914 4466 -3880
rect 4500 -3914 4512 -3880
rect 4454 -3952 4512 -3914
rect 4646 -3880 4704 -3874
rect 4646 -3914 4658 -3880
rect 4692 -3914 4704 -3880
rect 4646 -3952 4704 -3914
rect 4454 -3986 4466 -3952
rect 4500 -3986 4658 -3952
rect 4692 -3986 4704 -3952
rect 4454 -4032 4704 -3986
rect 4454 -4066 4466 -4032
rect 4500 -4066 4658 -4032
rect 4692 -4066 4704 -4032
rect 4454 -4104 4512 -4066
rect 4454 -4138 4466 -4104
rect 4500 -4138 4512 -4104
rect 4454 -4144 4512 -4138
rect 4646 -4104 4704 -4066
rect 4646 -4138 4658 -4104
rect 4692 -4138 4704 -4104
rect 4646 -4144 4704 -4138
rect 4840 -3880 4898 -3874
rect 4840 -3914 4852 -3880
rect 4886 -3914 4898 -3880
rect 4840 -3952 4898 -3914
rect 5032 -3880 5090 -3874
rect 5032 -3914 5044 -3880
rect 5078 -3914 5090 -3880
rect 5032 -3952 5090 -3914
rect 4840 -3986 4852 -3952
rect 4886 -3986 5044 -3952
rect 5078 -3986 5090 -3952
rect 4840 -4032 5090 -3986
rect 4840 -4066 4852 -4032
rect 4886 -4066 5044 -4032
rect 5078 -4066 5090 -4032
rect 4840 -4104 4898 -4066
rect 4840 -4138 4852 -4104
rect 4886 -4138 4898 -4104
rect 4840 -4144 4898 -4138
rect 5032 -4104 5090 -4066
rect 5032 -4138 5044 -4104
rect 5078 -4138 5090 -4104
rect 5032 -4144 5090 -4138
rect 5224 -3880 5282 -3874
rect 5224 -3914 5236 -3880
rect 5270 -3914 5282 -3880
rect 5224 -3952 5282 -3914
rect 5416 -3880 5474 -3874
rect 5416 -3914 5428 -3880
rect 5462 -3914 5474 -3880
rect 5416 -3952 5474 -3914
rect 5608 -3880 5666 -3874
rect 5608 -3914 5620 -3880
rect 5654 -3914 5666 -3880
rect 5608 -3952 5666 -3914
rect 5800 -3880 5858 -3874
rect 5800 -3914 5812 -3880
rect 5846 -3914 5858 -3880
rect 5800 -3952 5858 -3914
rect 5224 -3986 5236 -3952
rect 5270 -3986 5428 -3952
rect 5462 -3986 5620 -3952
rect 5654 -3986 5812 -3952
rect 5846 -3986 5858 -3952
rect 5224 -4032 5858 -3986
rect 5224 -4066 5236 -4032
rect 5270 -4066 5428 -4032
rect 5462 -4066 5620 -4032
rect 5654 -4066 5812 -4032
rect 5846 -4066 5858 -4032
rect 5224 -4104 5282 -4066
rect 5224 -4138 5236 -4104
rect 5270 -4138 5282 -4104
rect 5224 -4144 5282 -4138
rect 5416 -4104 5474 -4066
rect 5416 -4138 5428 -4104
rect 5462 -4138 5474 -4104
rect 5416 -4144 5474 -4138
rect 5608 -4104 5666 -4066
rect 5608 -4138 5620 -4104
rect 5654 -4138 5666 -4104
rect 5608 -4144 5666 -4138
rect 5800 -4104 5858 -4066
rect 5800 -4138 5812 -4104
rect 5846 -4138 5858 -4104
rect 5800 -4144 5858 -4138
rect 3596 -4194 3644 -4182
rect 3596 -4570 3603 -4194
rect 3637 -4570 3644 -4194
rect 3596 -4648 3644 -4570
rect 3690 -4194 3742 -4178
rect 3690 -4586 3742 -4572
rect 3788 -4194 3836 -4182
rect 3788 -4570 3795 -4194
rect 3829 -4570 3836 -4194
rect 3788 -4648 3836 -4570
rect 3882 -4194 3934 -4178
rect 3882 -4586 3934 -4572
rect 3980 -4194 4028 -4182
rect 3980 -4570 3987 -4194
rect 4021 -4570 4028 -4194
rect 3980 -4648 4028 -4570
rect 4074 -4194 4126 -4178
rect 4074 -4586 4126 -4572
rect 4172 -4194 4220 -4182
rect 4172 -4570 4179 -4194
rect 4213 -4570 4220 -4194
rect 4172 -4648 4220 -4570
rect 4266 -4194 4318 -4178
rect 4266 -4586 4318 -4572
rect 4364 -4194 4412 -4182
rect 4364 -4570 4371 -4194
rect 4405 -4570 4412 -4194
rect 4364 -4648 4412 -4570
rect 4458 -4194 4510 -4178
rect 4458 -4586 4510 -4572
rect 4556 -4194 4604 -4182
rect 4556 -4570 4563 -4194
rect 4597 -4570 4604 -4194
rect 4556 -4648 4604 -4570
rect 4650 -4194 4702 -4178
rect 4650 -4586 4702 -4572
rect 4748 -4194 4796 -4182
rect 4748 -4570 4755 -4194
rect 4789 -4570 4796 -4194
rect 4748 -4648 4796 -4570
rect 4842 -4194 4894 -4178
rect 4842 -4586 4894 -4572
rect 4940 -4194 4988 -4182
rect 4940 -4570 4947 -4194
rect 4981 -4570 4988 -4194
rect 4940 -4648 4988 -4570
rect 5034 -4194 5086 -4178
rect 5034 -4586 5086 -4572
rect 5132 -4194 5180 -4182
rect 5132 -4570 5139 -4194
rect 5173 -4570 5180 -4194
rect 5132 -4648 5180 -4570
rect 5226 -4194 5278 -4178
rect 5226 -4586 5278 -4572
rect 5324 -4194 5372 -4182
rect 5324 -4570 5331 -4194
rect 5365 -4570 5372 -4194
rect 5324 -4648 5372 -4570
rect 5418 -4194 5470 -4178
rect 5418 -4586 5470 -4572
rect 5516 -4194 5564 -4182
rect 5516 -4570 5523 -4194
rect 5557 -4570 5564 -4194
rect 5516 -4648 5564 -4570
rect 5610 -4194 5662 -4178
rect 5610 -4586 5662 -4572
rect 5708 -4194 5756 -4182
rect 5708 -4570 5715 -4194
rect 5749 -4570 5756 -4194
rect 5708 -4648 5756 -4570
rect 5802 -4194 5854 -4178
rect 5802 -4586 5854 -4572
rect 5900 -4194 5948 -4182
rect 5900 -4570 5907 -4194
rect 5941 -4570 5948 -4194
rect 5900 -4648 5948 -4570
rect 3596 -4678 5948 -4648
rect 3596 -4712 3696 -4678
rect 5848 -4712 5948 -4678
rect 3596 -4728 5948 -4712
rect 133 -5370 191 -5364
rect 133 -5404 145 -5370
rect 179 -5404 191 -5370
rect 133 -5442 191 -5404
rect 133 -5476 145 -5442
rect 179 -5476 191 -5442
rect 133 -5482 191 -5476
rect 44 -5532 90 -5520
rect 44 -5908 50 -5532
rect 84 -5908 90 -5532
rect 44 -5920 90 -5908
rect 137 -5532 189 -5516
rect 137 -5924 189 -5910
rect 236 -5532 282 -5520
rect 236 -5908 242 -5532
rect 276 -5908 282 -5532
rect 236 -5920 282 -5908
rect 332 -5532 378 -5520
rect 332 -5908 338 -5532
rect 372 -5908 378 -5532
rect 332 -5920 378 -5908
<< via1 >>
rect 3690 -4570 3699 -4194
rect 3699 -4570 3733 -4194
rect 3733 -4570 3742 -4194
rect 3690 -4572 3742 -4570
rect 3882 -4570 3891 -4194
rect 3891 -4570 3925 -4194
rect 3925 -4570 3934 -4194
rect 3882 -4572 3934 -4570
rect 4074 -4570 4083 -4194
rect 4083 -4570 4117 -4194
rect 4117 -4570 4126 -4194
rect 4074 -4572 4126 -4570
rect 4266 -4570 4275 -4194
rect 4275 -4570 4309 -4194
rect 4309 -4570 4318 -4194
rect 4266 -4572 4318 -4570
rect 4458 -4570 4467 -4194
rect 4467 -4570 4501 -4194
rect 4501 -4570 4510 -4194
rect 4458 -4572 4510 -4570
rect 4650 -4570 4659 -4194
rect 4659 -4570 4693 -4194
rect 4693 -4570 4702 -4194
rect 4650 -4572 4702 -4570
rect 4842 -4570 4851 -4194
rect 4851 -4570 4885 -4194
rect 4885 -4570 4894 -4194
rect 4842 -4572 4894 -4570
rect 5034 -4570 5043 -4194
rect 5043 -4570 5077 -4194
rect 5077 -4570 5086 -4194
rect 5034 -4572 5086 -4570
rect 5226 -4570 5235 -4194
rect 5235 -4570 5269 -4194
rect 5269 -4570 5278 -4194
rect 5226 -4572 5278 -4570
rect 5418 -4570 5427 -4194
rect 5427 -4570 5461 -4194
rect 5461 -4570 5470 -4194
rect 5418 -4572 5470 -4570
rect 5610 -4570 5619 -4194
rect 5619 -4570 5653 -4194
rect 5653 -4570 5662 -4194
rect 5610 -4572 5662 -4570
rect 5802 -4570 5811 -4194
rect 5811 -4570 5845 -4194
rect 5845 -4570 5854 -4194
rect 5802 -4572 5854 -4570
rect 137 -5908 146 -5532
rect 146 -5908 180 -5532
rect 180 -5908 189 -5532
rect 137 -5910 189 -5908
<< metal2 >>
rect 3687 -4194 3744 -4178
rect 3687 -4586 3744 -4572
rect 3879 -4194 3936 -4178
rect 3879 -4586 3936 -4572
rect 4071 -4194 4128 -4178
rect 4071 -4586 4128 -4572
rect 4263 -4194 4320 -4178
rect 4263 -4586 4320 -4572
rect 4455 -4194 4512 -4178
rect 4455 -4586 4512 -4572
rect 4647 -4194 4704 -4178
rect 4647 -4586 4704 -4572
rect 4840 -4194 4897 -4178
rect 4840 -4586 4897 -4572
rect 5032 -4194 5089 -4178
rect 5032 -4586 5089 -4572
rect 5224 -4194 5281 -4178
rect 5224 -4586 5281 -4572
rect 5416 -4194 5473 -4178
rect 5416 -4586 5473 -4572
rect 5608 -4194 5665 -4178
rect 5608 -4586 5665 -4572
rect 5800 -4194 5857 -4178
rect 5800 -4586 5857 -4572
rect 134 -5532 191 -5516
rect 134 -5924 191 -5910
<< via2 >>
rect 3687 -4572 3690 -4194
rect 3690 -4572 3742 -4194
rect 3742 -4572 3744 -4194
rect 3879 -4572 3882 -4194
rect 3882 -4572 3934 -4194
rect 3934 -4572 3936 -4194
rect 4071 -4572 4074 -4194
rect 4074 -4572 4126 -4194
rect 4126 -4572 4128 -4194
rect 4263 -4572 4266 -4194
rect 4266 -4572 4318 -4194
rect 4318 -4572 4320 -4194
rect 4455 -4572 4458 -4194
rect 4458 -4572 4510 -4194
rect 4510 -4572 4512 -4194
rect 4647 -4572 4650 -4194
rect 4650 -4572 4702 -4194
rect 4702 -4572 4704 -4194
rect 4840 -4572 4842 -4194
rect 4842 -4572 4894 -4194
rect 4894 -4572 4897 -4194
rect 5032 -4572 5034 -4194
rect 5034 -4572 5086 -4194
rect 5086 -4572 5089 -4194
rect 5224 -4572 5226 -4194
rect 5226 -4572 5278 -4194
rect 5278 -4572 5281 -4194
rect 5416 -4572 5418 -4194
rect 5418 -4572 5470 -4194
rect 5470 -4572 5473 -4194
rect 5608 -4572 5610 -4194
rect 5610 -4572 5662 -4194
rect 5662 -4572 5665 -4194
rect 5800 -4572 5802 -4194
rect 5802 -4572 5854 -4194
rect 5854 -4572 5857 -4194
rect 134 -5910 137 -5532
rect 137 -5910 189 -5532
rect 189 -5910 191 -5532
<< metal3 >>
rect 3682 -4194 3750 -3986
rect 3682 -4572 3687 -4194
rect 3744 -4572 3750 -4194
rect 3682 -4586 3750 -4572
rect 3874 -4194 3942 -3986
rect 3874 -4572 3879 -4194
rect 3936 -4572 3942 -4194
rect 3874 -4586 3942 -4572
rect 4066 -4194 4134 -3986
rect 4066 -4572 4071 -4194
rect 4128 -4572 4134 -4194
rect 4066 -4586 4134 -4572
rect 4258 -4194 4326 -3986
rect 4258 -4572 4263 -4194
rect 4320 -4572 4326 -4194
rect 4258 -4586 4326 -4572
rect 4450 -4194 4518 -3986
rect 4450 -4572 4455 -4194
rect 4512 -4572 4518 -4194
rect 4450 -4586 4518 -4572
rect 4642 -4194 4710 -3986
rect 4642 -4572 4647 -4194
rect 4704 -4572 4710 -4194
rect 4642 -4586 4710 -4572
rect 4834 -4194 4902 -4178
rect 4834 -4572 4840 -4194
rect 4897 -4572 4902 -4194
rect 4834 -4586 4902 -4572
rect 5026 -4194 5094 -4178
rect 5026 -4572 5032 -4194
rect 5089 -4572 5094 -4194
rect 5026 -4586 5094 -4572
rect 5218 -4194 5286 -4178
rect 5218 -4572 5224 -4194
rect 5281 -4572 5286 -4194
rect 5218 -4586 5286 -4572
rect 5410 -4194 5478 -4178
rect 5410 -4572 5416 -4194
rect 5473 -4572 5478 -4194
rect 5410 -4586 5478 -4572
rect 5602 -4194 5670 -4178
rect 5602 -4572 5608 -4194
rect 5665 -4572 5670 -4194
rect 5602 -4586 5670 -4572
rect 5794 -4194 5862 -4178
rect 5794 -4572 5800 -4194
rect 5857 -4572 5862 -4194
rect 5794 -4586 5862 -4572
rect 129 -5532 197 -5516
rect 129 -5910 134 -5532
rect 191 -5910 197 -5532
rect 129 -5924 197 -5910
<< comment >>
rect 3644 -3040 3658 -3010
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_0 ~/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hs/mag
timestamp 1666464484
transform 1 0 2390 0 -1 -3327
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_2
timestamp 1666464484
transform 1 0 2390 0 1 -4659
box -38 -49 902 715
<< end >>
