* NGSPICE file created from imirror2.ext - technology: sky130A

.subckt imirror2 IN OUT VLO VHI
X0 VHI a_4493_207# a_4493_207# VHI.t5 sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X1 a_4493_207# VLO.t6 VLO.t8 VLO.t7 sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X2 VLO.t5 VLO.t3 OUT VLO.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X3 a_5868_1637# a_5468_1540# OUT VHI.t0 sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X4 OUT OUT.t0 VLO VLO.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=2e+06u
X5 VLO IN.t0 a_4493_207# VLO.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X6 a_4493_207# a_4094_1540# a_4036_1637# VHI.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X7 OUT a_4493_207# VHI VHI.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
R0 VHI.t2 VHI.t0 178.465
R1 VHI.t5 VHI.t1 178.465
R2 VHI.t0 VHI.n1 133.656
R3 VHI.t1 VHI.n3 133.656
R4 VHI.n6 VHI.t2 89.232
R5 VHI.n6 VHI.t5 89.232
R6 VHI.n9 VHI.n8 3.388
R7 VHI VHI.n9 1.702
R8 VHI.n5 VHI.n4 0.002
R9 VHI.n6 VHI.n5 0.002
R10 VHI.n8 VHI.n7 0.002
R11 VHI.n7 VHI.n6 0.002
R12 VHI.n3 VHI.n2 0.002
R13 VHI.n1 VHI.n0 0.002
R14 VLO.n4 VLO.t4 1062.83
R15 VLO.n7 VLO.t7 1062.83
R16 VLO.n15 VLO.t0 709.577
R17 VLO.n15 VLO.t9 709.577
R18 VLO.n13 VLO.n11 344.847
R19 VLO.n13 VLO.n12 344.847
R20 VLO.n6 VLO.n5 264.873
R21 VLO.n9 VLO.n8 264.496
R22 VLO.n21 VLO.n19 202.541
R23 VLO.n2 VLO.n0 202.541
R24 VLO.t6 VLO.n20 153.089
R25 VLO.n21 VLO.t6 153.089
R26 VLO.n2 VLO.t3 153.089
R27 VLO.t3 VLO.n1 153.089
R28 VLO.n22 VLO.n21 32.935
R29 VLO.n3 VLO.n2 32.935
R30 VLO.n24 VLO.n9 10.039
R31 VLO.n24 VLO.n6 10.037
R32 VLO.n24 VLO.n18 8.178
R33 VLO.n24 VLO.n23 8.178
R34 VLO.n23 VLO.n22 8.01
R35 VLO.n6 VLO.n3 6.032
R36 VLO.n24 VLO.n17 3.765
R37 VLO.n19 VLO.t8 3.48
R38 VLO.n0 VLO.t5 3.48
R39 VLO VLO.n24 1.562
R40 VLO.n17 VLO.n10 1.127
R41 VLO.n17 VLO.n16 0.014
R42 VLO.n16 VLO.n15 0.014
R43 VLO.n8 VLO.n7 0.012
R44 VLO.n5 VLO.n4 0.012
R45 VLO.n14 VLO.n13 0.007
R46 VLO.n15 VLO.n14 0.007
R47 OUT OUT.t0 68.216
R48 IN IN.t0 67.356
C0 a_4036_1637# OUT 0.03fF
C1 a_5468_1540# OUT 0.53fF
C2 a_4036_1637# VHI 0.69fF
C3 a_4036_1637# a_4493_207# 0.63fF
C4 a_5468_1540# VHI 0.99fF
C5 a_5468_1540# a_4493_207# 0.22fF
C6 a_4036_1637# a_4094_1540# 0.15fF
C7 a_5468_1540# a_4094_1540# 0.00fF
C8 VHI OUT 1.31fF
C9 OUT a_4493_207# 0.87fF
C10 OUT a_4094_1540# 0.10fF
C11 VHI a_4493_207# 3.26fF
C12 VHI a_4094_1540# 1.00fF
C13 a_4094_1540# a_4493_207# 0.44fF
C14 a_4036_1637# IN 0.01fF
C15 OUT IN 0.25fF
C16 a_5868_1637# a_5468_1540# 0.15fF
C17 VHI IN 0.19fF
C18 IN a_4493_207# 0.76fF
C19 IN a_4094_1540# 0.16fF
C20 a_5468_1540# a_4036_1637# 0.01fF
C21 a_5868_1637# OUT 0.47fF
C22 a_5868_1637# VHI 0.45fF
C23 a_5868_1637# a_4493_207# 0.22fF
C24 a_5868_1637# a_4094_1540# 0.01fF
.ends

