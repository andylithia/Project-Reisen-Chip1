* NGSPICE file created from cmota_gb_rp_gp.ext - technology: sky130A

.subckt cmota_gb_rp_gp VIN VIP VHI VLO SBAR S VREF VOP VREF_GATED
X0 gated_iref_fix_0/imirror2_0/OUT gated_iref_fix_0/a_1444_106# VLO sky130_fd_pr__res_xhigh_po w=350000u l=1.49e+06u
X1 VLO SBAR VREF_GATED VLO sky130_fd_pr__nfet_01v8 ad=4.395e+13p pd=3.12545e+08u as=1.65e+12p ps=1.132e+07u w=2.5e+06u l=150000u
X2 VLO VREF_GATED sky130_fd_pr__cap_mim_m3_1 l=6.2e+06u w=2.76e+07u
X3 VREF_GATED VLO sky130_fd_pr__cap_mim_m3_2 l=6.2e+06u w=2.76e+07u
X4 VREF_GATED S gated_iref_fix_0/a_1444_106# VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X5 VLO VLO gated_iref_fix_0/a_1444_106# VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X6 VREF_GATED SBAR VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X7 gated_iref_fix_0/a_1444_106# S VREF_GATED VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X8 cmota_gb_rp_0/VMN cmota_gb_rp_0/li_5300_n960# VLO sky130_fd_pr__res_high_po w=690000u l=5.83e+06u
X9 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/VMN VHI sky130_fd_pr__pfet_01v8 ad=5.22e+13p pd=3.7044e+08u as=0p ps=0u w=1e+07u l=300000u
X10 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X11 VHI cmota_gb_rp_0/DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+13p ps=8.232e+07u w=1e+07u l=300000u
X12 cmota_gb_rp_0/DN VIN cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X13 cmota_gb_rp_0/COM VIN cmota_gb_rp_0/DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X14 cmota_gb_rp_0/DP VIP cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X15 cmota_gb_rp_0/VMN cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X16 cmota_gb_rp_0/VMN cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X17 VHI VHI VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X18 cmota_gb_rp_0/a_2925_285# cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X19 cmota_gb_rp_0/DP VIP cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X20 cmota_gb_rp_0/li_5300_n960# VOP sky130_fd_pr__cap_mim_m3_2 l=1.32e+07u w=3.7e+06u
X21 VOP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X22 VOP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X23 VOP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X24 cmota_gb_rp_0/COM VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X25 VLO cmota_gb_rp_0/VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.116e+07u w=1e+07u l=300000u
X26 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X27 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X28 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X29 VHI cmota_gb_rp_0/DP cmota_gb_rp_0/DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X30 cmota_gb_rp_0/COM VIP cmota_gb_rp_0/DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X31 VLO VREF_GATED cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X32 cmota_gb_rp_0/VMN VHI VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X33 cmota_gb_rp_0/DN cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X34 VHI cmota_gb_rp_0/DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X35 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X36 VLO VREF_GATED cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X37 cmota_gb_rp_0/COM VIN cmota_gb_rp_0/DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X38 cmota_gb_rp_0/DN cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X39 cmota_gb_rp_0/DP cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X40 cmota_gb_rp_0/DN cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X41 cmota_gb_rp_0/DP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X42 cmota_gb_rp_0/DN VIN cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X43 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X44 cmota_gb_rp_0/COM VIP cmota_gb_rp_0/DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X45 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X46 VOP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X47 cmota_gb_rp_0/VMN cmota_gb_rp_0/VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X48 VLO cmota_gb_rp_0/VMN cmota_gb_rp_0/VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X49 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X50 VOP cmota_gb_rp_0/VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X51 VHI cmota_gb_rp_0/DP cmota_gb_rp_0/DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X52 VLO cmota_gb_rp_0/VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X53 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X54 VLO VLO cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X55 cmota_gb_rp_0/DN VIN cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X56 VHI cmota_gb_rp_0/DP cmota_gb_rp_0/a_2217_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X57 VHI cmota_gb_rp_0/DP cmota_gb_rp_0/DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X58 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X59 cmota_gb_rp_0/COM VREF_GATED VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X60 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X61 cmota_gb_rp_0/COM VIN cmota_gb_rp_0/DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X62 cmota_gb_rp_0/COM VREF_GATED VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X63 cmota_gb_rp_0/DP VIP cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X64 cmota_gb_rp_0/COM VIN cmota_gb_rp_0/DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X65 cmota_gb_rp_0/VMN cmota_gb_rp_0/DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X66 cmota_gb_rp_0/DP cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X67 cmota_gb_rp_0/DP VIP cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X68 cmota_gb_rp_0/a_2217_285# cmota_gb_rp_0/DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X69 cmota_gb_rp_0/VMN cmota_gb_rp_0/VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X70 cmota_gb_rp_0/COM VIP cmota_gb_rp_0/DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X71 VLO cmota_gb_rp_0/VMN cmota_gb_rp_0/VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X72 VOP cmota_gb_rp_0/VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X73 cmota_gb_rp_0/COM VIP cmota_gb_rp_0/DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X74 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X75 cmota_gb_rp_0/DN VIN cmota_gb_rp_0/COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X76 VOP cmota_gb_rp_0/li_5300_n960# sky130_fd_pr__cap_mim_m3_1 l=1.32e+07u w=3.7e+06u
X77 VHI cmota_gb_rp_0/DN cmota_gb_rp_0/a_2925_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X78 VHI cmota_gb_rp_0/DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X79 VLO VHI sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=1.3e+07u
X80 VHI VLO sky130_fd_pr__cap_mim_m3_1 l=3.1e+07u w=1.3e+07u
C0 cmota_gb_rp_0/DN VHI 17.11fF
C1 gated_iref_fix_0/imirror2_0/a_4493_207# VHI 3.45fF
C2 cmota_gb_rp_0/DN cmota_gb_rp_0/COM 6.05fF
C3 cmota_gb_rp_0/a_2925_285# VHI 4.36fF
C4 VHI VOP 18.33fF
C5 cmota_gb_rp_0/DP VHI 17.03fF
C6 VREF_GATED VHI 4.36fF
C7 cmota_gb_rp_0/DP cmota_gb_rp_0/COM 6.02fF
C8 VREF_GATED cmota_gb_rp_0/COM 2.52fF
C9 cmota_gb_rp_0/VMN VHI 17.90fF
C10 cmota_gb_rp_0/a_2217_285# VHI 4.36fF
C11 VHI cmota_gb_rp_0/li_5300_n960# 2.04fF
C12 cmota_gb_rp_0/li_5300_n960# VOP 9.33fF
Xgated_iref_fix_0/imirror2_0 gated_iref_fix_0/imirror2_0/OUT imirror2
C13 VREF_GATED VLO 54.32fF
C14 cmota_gb_rp_0/COM VLO 6.15fF $ **FLOATING
C15 VOP VLO 9.34fF
C16 cmota_gb_rp_0/li_5300_n960# VLO 3.02fF $ **FLOATING
C17 cmota_gb_rp_0/VMN VLO 14.09fF $ **FLOATING
C18 gated_iref_fix_0/imirror2_0/OUT VLO 6.93fF
C19 VHI VLO 135.56fF
C20 VREF VLO 7.50fF
C21 gated_iref_fix_0/imirror2_0/a_4493_207# VLO 4.63fF
.ends
